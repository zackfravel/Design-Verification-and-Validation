
module VQS64_4 ( mX1, mX2, mX3, mX4, mY1, mY2, mY3, mY4, mCLK );
  input [63:0] mX1;
  input [63:0] mX2;
  input [63:0] mX3;
  input [63:0] mX4;
  output [63:0] mY1;
  output [63:0] mY2;
  output [63:0] mY3;
  output [63:0] mY4;
  input mCLK;
  wire   N9, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22,
         N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36,
         N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50,
         N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64,
         N65, N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78,
         N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, N92,
         N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103, N104, N105,
         N106, N107, N108, N109, N110, N111, N112, N113, N114, N115, N116,
         N117, N118, N119, N120, N121, N122, N123, N124, N125, N126, N127,
         N128, N129, N130, N131, N132, N133, N134, N135, N136, N139, N140,
         N141, N142, N143, N144, N145, N146, N147, N148, N149, N150, N151,
         N152, N153, N154, N155, N156, N157, N158, N159, N160, N161, N162,
         N163, N164, N165, N166, N167, N168, N169, N170, N171, N172, N173,
         N174, N175, N176, N177, N178, N179, N180, N181, N182, N183, N184,
         N185, N186, N187, N188, N189, N190, N191, N192, N193, N194, N195,
         N196, N197, N198, N199, N200, N201, N202, N203, N204, N205, N206,
         N207, N208, N209, N210, N211, N212, N213, N214, N215, N216, N217,
         N218, N219, N220, N221, N222, N223, N224, N225, N226, N227, N228,
         N229, N230, N231, N232, N233, N234, N235, N236, N237, N238, N239,
         N240, N241, N242, N243, N244, N245, N246, N247, N248, N249, N250,
         N251, N252, N253, N254, N255, N256, N257, N258, N259, N260, N261,
         N262, N263, N264, N265, N266, N279, N280, N281, N282, N283, N284,
         N285, N286, N287, N288, N289, N290, N291, N292, N293, N294, N295,
         N296, N297, N298, N299, N300, N301, N302, N303, N304, N305, N306,
         N307, N308, N309, N310, N311, N312, N313, N314, N315, N316, N317,
         N318, N319, N320, N321, N322, N323, N324, N325, N326, N327, N328,
         N329, N330, N331, N332, N333, N334, N335, N336, N337, N338, N339,
         N340, N341, N342, N343, N344, N345, N346, N347, N348, N349, N350,
         N351, N352, N353, N354, N355, N356, N357, N358, N359, N360, N361,
         N362, N363, N364, N365, N366, N367, N368, N369, N370, N371, N372,
         N373, N374, N375, N376, N377, N378, N379, N380, N381, N382, N383,
         N384, N385, N386, N387, N388, N389, N390, N391, N392, N393, N394,
         N395, N396, N397, N398, N399, N400, N401, N402, N403, N404, N405,
         N406, N407, N408, N409, N410, N411, N412, N413, N414, N415, N416,
         N417, N418, N419, N420, N421, N422, N423, N424, N425, N426, N427,
         N428, N429, N430, N431, N432, N433, N434, N435, N436, N437, N438,
         N439, N440, N441, N442, N443, N444, N445, N446, N447, N448, N449,
         N450, N451, N452, N453, N454, N455, N456, N457, N458, N459, N460,
         N461, N462, N463, N464, N465, N466, N467, N468, N469, N470, N471,
         N472, N473, N474, N475, N476, N477, N478, N479, N480, N481, N482,
         N483, N484, N485, N486, N487, N488, N489, N490, N491, N492, N493,
         N494, N495, N496, N497, N498, N499, N500, N501, N502, N503, N504,
         N505, N506, N507, N508, N509, N510, N511, N512, N513, N514, N515,
         N516, N517, N518, N519, N520, N521, N522, N523, N524, N525, N526,
         N527, N528, N529, N530, N531, N532, N533, N534, N537, N538, N539,
         N540, N541, N542, N543, N544, N545, N546, N547, N548, N549, N550,
         N551, N552, N553, N554, N555, N556, N557, N558, N559, N560, N561,
         N562, N563, N564, N565, N566, N567, N568, N569, N570, N571, N572,
         N573, N574, N575, N576, N577, N578, N579, N580, N581, N582, N583,
         N584, N585, N586, N587, N588, N589, N590, N591, N592, N593, N594,
         N595, N596, N597, N598, N599, N600, N601, N602, N603, N604, N605,
         N606, N607, N608, N609, N610, N611, N612, N613, N614, N615, N616,
         N617, N618, N619, N620, N621, N622, N623, N624, N625, N626, N627,
         N628, N629, N630, N631, N632, N633, N634, N635, N636, N637, N638,
         N639, N640, N641, N642, N643, N644, N645, N646, N647, N648, N649,
         N650, N651, N652, N653, N654, N655, N656, N657, N658, N659, N660,
         N661, N662, N663, N664, n1863, n1864, n1865, n1866, n1867, n1868,
         n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878,
         n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888,
         n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898,
         n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908,
         n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918,
         n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928,
         n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938,
         n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948,
         n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958,
         n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968,
         n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978,
         n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988,
         n1989, n1990, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
         n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
         n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
         n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
         n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
         n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
         n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
         n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
         n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
         n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
         n2122, n2131, n2135, n2136, n2140, n2141, n2148, n2161, n2166, n2167,
         n2179, n2181, n2183, n2192, n2198, n2209, n2213, n2214, n2217, n2218,
         n2225, n2232, n2240, n2244, n2248, n2259, n2260, n2263, n2266, n2271,
         n2276, n2327, n2331, n2336, n2337, n2405, n2413, n2420, n2427, n2436,
         n2444, n2448, n2449, n2452, n2474, n2543, n2544, n2545, n2546, n2547,
         n2548, n2549, n2550, n2551, n2552, n2553, n2555, n2556, n2557, n2558,
         n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568,
         n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578,
         n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588,
         n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598,
         n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608,
         n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618,
         n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628,
         n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638,
         n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648,
         n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658,
         n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668,
         n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678,
         n2679, n2680, n2681, n2682, n2684, n2685, n2686, n2687, n2688, n2689,
         n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699,
         n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709,
         n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719,
         n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729,
         n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739,
         n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749,
         n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759,
         n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
         n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779,
         n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789,
         n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799,
         n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809,
         n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819,
         n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829,
         n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839,
         n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849,
         n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859,
         n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869,
         n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879,
         n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889,
         n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899,
         n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909,
         n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919,
         n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929,
         n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939,
         n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949,
         n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959,
         n2960, n2970, n2972, n2978, n2979, n2983, n2984, n2985, n2986, n2987,
         n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2997, n2998, n2999,
         n3000, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015,
         n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025,
         n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035,
         n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045,
         n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055,
         n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065,
         n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075,
         n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085,
         n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095,
         n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105,
         n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115,
         n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125,
         n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135,
         n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145,
         n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155,
         n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165,
         n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175,
         n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185,
         n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195,
         n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205,
         n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215,
         n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225,
         n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235,
         n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245,
         n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255,
         n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265,
         n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275,
         n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285,
         n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295,
         n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305,
         n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315,
         n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325,
         n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335,
         n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345,
         n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355,
         n3356, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378,
         n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388,
         n3389, n3390, n3391, n3392, n3395, n3396, n3397, n3398, n3399, n3400,
         n3401, n3402, n3403, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3425, n3426, n3427, n3428, n3429, n3431, n3444, n3445, n3446, n3447,
         n3448, n3449, n3450, n3452, n3454, n3455, n3456, n3459, n3460, n3461,
         n3462, n3463, n3464, n3468, n3469, n3470, n3471, n3472, n3473, n3475,
         n3476, n3478, n3480, n3481, n3482, n3483, n3486, n3487, n3488, n3489,
         n3490, n3491, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500,
         n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510,
         n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520,
         n3521, n3522, n3523, n3524, n3525, n3598, n3606, n3609, n3610, n3611,
         n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
         n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
         n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
         n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
         n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
         n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
         n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879;
  wire   [63:0] rC1;
  wire   [63:0] rC2;
  wire   [63:0] rC3;
  wire   [63:0] rC4;
  wire   [63:0] rC5;
  wire   [63:0] rC6;
  wire   [63:0] rC7;
  wire   [63:0] rC8;

  DFF_X1 \rC1_reg[63]  ( .D(N72), .CK(mCLK), .Q(rC1[63]), .QN(n3338) );
  DFF_X1 \rC1_reg[62]  ( .D(N71), .CK(mCLK), .Q(rC1[62]), .QN(n3328) );
  DFF_X1 \rC1_reg[61]  ( .D(N70), .CK(mCLK), .Q(rC1[61]), .QN(n3206) );
  DFF_X1 \rC1_reg[60]  ( .D(N69), .CK(mCLK), .Q(rC1[60]), .QN(n3262) );
  DFF_X1 \rC1_reg[59]  ( .D(N68), .CK(mCLK), .Q(rC1[59]), .QN(n3293) );
  DFF_X1 \rC1_reg[58]  ( .D(N67), .CK(mCLK), .Q(rC1[58]), .QN(n3051) );
  DFF_X1 \rC1_reg[57]  ( .D(N66), .CK(mCLK), .Q(rC1[57]), .QN(n3197) );
  DFF_X1 \rC1_reg[56]  ( .D(N65), .CK(mCLK), .Q(rC1[56]), .QN(n3302) );
  DFF_X1 \rC1_reg[55]  ( .D(N64), .CK(mCLK), .Q(rC1[55]), .QN(n3240) );
  DFF_X1 \rC1_reg[54]  ( .D(N63), .CK(mCLK), .Q(rC1[54]), .QN(n3073) );
  DFF_X1 \rC1_reg[53]  ( .D(N62), .CK(mCLK), .Q(rC1[53]), .QN(n3230) );
  DFF_X1 \rC1_reg[52]  ( .D(N61), .CK(mCLK), .Q(rC1[52]), .QN(n3287) );
  DFF_X1 \rC1_reg[51]  ( .D(N60), .CK(mCLK), .Q(rC1[51]), .QN(n3056) );
  DFF_X1 \rC1_reg[50]  ( .D(N59), .CK(mCLK), .Q(rC1[50]), .QN(n3313) );
  DFF_X1 \rC1_reg[49]  ( .D(N58), .CK(mCLK), .Q(rC1[49]), .QN(n3172) );
  DFF_X1 \rC1_reg[48]  ( .D(N57), .CK(mCLK), .Q(rC1[48]), .QN(n3187) );
  DFF_X1 \rC1_reg[47]  ( .D(N56), .CK(mCLK), .Q(rC1[47]), .QN(n3021) );
  DFF_X1 \rC1_reg[46]  ( .D(N55), .CK(mCLK), .Q(rC1[46]), .QN(n3113) );
  DFF_X1 \rC1_reg[45]  ( .D(N54), .CK(mCLK), .Q(rC1[45]), .QN(n3226) );
  DFF_X1 \rC1_reg[44]  ( .D(N53), .CK(mCLK), .Q(rC1[44]), .QN(n3162) );
  DFF_X1 \rC1_reg[43]  ( .D(N52), .CK(mCLK), .Q(rC1[43]), .QN(n3291) );
  DFF_X1 \rC1_reg[42]  ( .D(N51), .CK(mCLK), .Q(rC1[42]), .QN(n3078) );
  DFF_X1 \rC1_reg[41]  ( .D(N50), .CK(mCLK), .Q(rC1[41]), .QN(n3228) );
  DFF_X1 \rC1_reg[40]  ( .D(N49), .CK(mCLK), .Q(rC1[40]), .QN(n3330) );
  DFF_X1 \rC1_reg[39]  ( .D(N48), .CK(mCLK), .Q(rC1[39]), .QN(n3289) );
  DFF_X1 \rC1_reg[38]  ( .D(N47), .CK(mCLK), .Q(rC1[38]), .QN(n3346) );
  DFF_X1 \rC1_reg[37]  ( .D(N46), .CK(mCLK), .Q(rC1[37]), .QN(n3245) );
  DFF_X1 \rC1_reg[36]  ( .D(N45), .CK(mCLK), .Q(rC1[36]), .QN(n3178) );
  DFF_X1 \rC1_reg[35]  ( .D(N44), .CK(mCLK), .Q(rC1[35]), .QN(n3149) );
  DFF_X1 \rC1_reg[34]  ( .D(N43), .CK(mCLK), .Q(rC1[34]), .QN(n3049) );
  DFF_X1 \rC1_reg[33]  ( .D(N42), .CK(mCLK), .Q(rC1[33]), .QN(n3195) );
  DFF_X1 \rC1_reg[32]  ( .D(N41), .CK(mCLK), .Q(rC1[32]), .QN(n3299) );
  DFF_X1 \rC1_reg[31]  ( .D(N40), .CK(mCLK), .Q(rC1[31]), .QN(n3238) );
  DFF_X1 \rC1_reg[30]  ( .D(N39), .CK(mCLK), .Q(rC1[30]), .QN(n3072) );
  DFF_X1 \rC1_reg[29]  ( .D(N38), .CK(mCLK), .Q(rC1[29]), .QN(n3229) );
  DFF_X1 \rC1_reg[28]  ( .D(N37), .CK(mCLK), .Q(rC1[28]), .QN(n3331) );
  DFF_X1 \rC1_reg[27]  ( .D(N36), .CK(mCLK), .Q(rC1[27]), .QN(n3290) );
  DFF_X1 \rC1_reg[26]  ( .D(N35), .CK(mCLK), .Q(rC1[26]), .QN(n3235) );
  DFF_X1 \rC1_reg[25]  ( .D(N34), .CK(mCLK), .Q(rC1[25]), .QN(n3079) );
  DFF_X1 \rC1_reg[24]  ( .D(N33), .CK(mCLK), .Q(rC1[24]), .QN(n3189) );
  DFF_X1 \rC1_reg[23]  ( .D(N32), .CK(mCLK), .Q(rC1[23]), .QN(n3150) );
  DFF_X1 \rC1_reg[22]  ( .D(N31), .CK(mCLK), .Q(rC1[22]), .QN(n3014) );
  DFF_X1 \rC1_reg[21]  ( .D(N30), .CK(mCLK), .Q(rC1[21]), .QN(n3130) );
  DFF_X1 \rC1_reg[20]  ( .D(N29), .CK(mCLK), .Q(rC1[20]), .QN(n3340) );
  DFF_X1 \rC1_reg[19]  ( .D(N28), .CK(mCLK), .Q(rC1[19]), .QN(n3171) );
  DFF_X1 \rC1_reg[18]  ( .D(N27), .CK(mCLK), .Q(rC1[18]), .QN(n3263) );
  DFF_X1 \rC1_reg[17]  ( .D(N26), .CK(mCLK), .Q(rC1[17]), .QN(n3294) );
  DFF_X1 \rC1_reg[16]  ( .D(N25), .CK(mCLK), .Q(rC1[16]), .QN(n3052) );
  DFF_X1 \rC1_reg[15]  ( .D(N24), .CK(mCLK), .Q(rC1[15]), .QN(n3370) );
  DFF_X1 \rC1_reg[14]  ( .D(N23), .CK(mCLK), .Q(rC1[14]), .QN(n3382) );
  DFF_X1 \rC1_reg[13]  ( .D(N22), .CK(mCLK), .Q(rC1[13]), .QN(n3118) );
  DFF_X1 \rC1_reg[12]  ( .D(N21), .CK(mCLK), .Q(rC1[12]), .QN(n3417) );
  DFF_X1 \rC1_reg[11]  ( .D(N20), .CK(mCLK), .Q(rC1[11]), .QN(n3296) );
  DFF_X1 \rC1_reg[10]  ( .D(N19), .CK(mCLK), .Q(rC1[10]), .QN(n3151) );
  DFF_X1 \rC1_reg[9]  ( .D(N18), .CK(mCLK), .Q(n3376), .QN(n3419) );
  DFF_X1 \rC1_reg[8]  ( .D(N17), .CK(mCLK), .Q(n3387), .QN(n3606) );
  DFF_X1 \rC1_reg[7]  ( .D(N16), .CK(mCLK), .Q(rC1[7]), .QN(n3420) );
  DFF_X1 \rC1_reg[6]  ( .D(N15), .CK(mCLK), .Q(rC1[6]), .QN(n3167) );
  DFF_X1 \rC1_reg[5]  ( .D(N14), .CK(mCLK), .Q(rC1[5]), .QN(n3334) );
  DFF_X1 \rC1_reg[4]  ( .D(N13), .CK(mCLK), .Q(rC1[4]), .QN(n3185) );
  DFF_X1 \rC1_reg[3]  ( .D(N12), .CK(mCLK), .Q(rC1[3]), .QN(n3252) );
  DFF_X1 \rC1_reg[2]  ( .D(N11), .CK(mCLK), .Q(rC1[2]), .QN(n3304) );
  DFF_X1 \rC1_reg[1]  ( .D(N10), .CK(mCLK), .Q(rC1[1]), .QN(n3242) );
  DFF_X1 \rC1_reg[0]  ( .D(N9), .CK(mCLK), .Q(rC1[0]), .QN(n3139) );
  DFF_X1 \rC4_reg[63]  ( .D(N266), .CK(mCLK), .Q(rC4[63]), .QN(n3077) );
  DFF_X1 \rC4_reg[62]  ( .D(N265), .CK(mCLK), .Q(rC4[62]), .QN(n3081) );
  DFF_X1 \rC4_reg[61]  ( .D(N264), .CK(mCLK), .Q(rC4[61]), .QN(n3140) );
  DFF_X1 \rC4_reg[60]  ( .D(N263), .CK(mCLK), .Q(rC4[60]), .QN(n3010) );
  DFF_X1 \rC4_reg[59]  ( .D(N262), .CK(mCLK), .Q(rC4[59]), .QN(n3082) );
  DFF_X1 \rC4_reg[58]  ( .D(N261), .CK(mCLK), .Q(rC4[58]), .QN(n3300) );
  DFF_X1 \rC4_reg[57]  ( .D(N260), .CK(mCLK), .Q(rC4[57]), .QN(n3138) );
  DFF_X1 \rC4_reg[56]  ( .D(N259), .CK(mCLK), .Q(rC4[56]), .QN(n3045) );
  DFF_X1 \rC4_reg[55]  ( .D(N258), .CK(mCLK), .Q(rC4[55]), .QN(n3156) );
  DFF_X1 \rC4_reg[54]  ( .D(N257), .CK(mCLK), .Q(rC4[54]), .QN(n3326) );
  DFF_X1 \rC4_reg[53]  ( .D(N256), .CK(mCLK), .Q(rC4[53]), .QN(n3146) );
  DFF_X1 \rC4_reg[52]  ( .D(N255), .CK(mCLK), .Q(rC4[52]), .QN(n3031) );
  DFF_X1 \rC4_reg[51]  ( .D(N254), .CK(mCLK), .Q(rC4[51]), .QN(n3323) );
  DFF_X1 \rC4_reg[50]  ( .D(N253), .CK(mCLK), .Q(rC4[50]), .QN(n3067) );
  DFF_X1 \rC4_reg[49]  ( .D(N252), .CK(mCLK), .Q(rC4[49]), .QN(n3020) );
  DFF_X1 \rC4_reg[48]  ( .D(N251), .CK(mCLK), .Q(rC4[48]), .QN(n3103) );
  DFF_X1 \rC4_reg[47]  ( .D(N250), .CK(mCLK), .Q(rC4[47]), .QN(n3316) );
  DFF_X1 \rC4_reg[46]  ( .D(N249), .CK(mCLK), .Q(rC4[46]), .QN(n3233) );
  DFF_X1 \rC4_reg[45]  ( .D(N248), .CK(mCLK), .Q(rC4[45]), .QN(n3166) );
  DFF_X1 \rC4_reg[44]  ( .D(N247), .CK(mCLK), .Q(rC4[44]), .QN(n3222) );
  DFF_X1 \rC4_reg[43]  ( .D(N246), .CK(mCLK), .Q(rC4[43]), .QN(n3070) );
  DFF_X1 \rC4_reg[42]  ( .D(N245), .CK(mCLK), .Q(rC4[42]), .QN(n3105) );
  DFF_X1 \rC4_reg[41]  ( .D(N244), .CK(mCLK), .Q(rC4[41]), .QN(n3308) );
  DFF_X1 \rC4_reg[40]  ( .D(N243), .CK(mCLK), .Q(rC4[40]), .QN(n3243) );
  DFF_X1 \rC4_reg[39]  ( .D(N242), .CK(mCLK), .Q(rC4[39]), .QN(n3121) );
  DFF_X1 \rC4_reg[38]  ( .D(N241), .CK(mCLK), .Q(rC4[38]), .QN(n3333) );
  DFF_X1 \rC4_reg[37]  ( .D(N240), .CK(mCLK), .Q(rC4[37]), .QN(n3190) );
  DFF_X1 \rC4_reg[36]  ( .D(N239), .CK(mCLK), .Q(rC4[36]), .QN(n3177) );
  DFF_X1 \rC4_reg[35]  ( .D(N238), .CK(mCLK), .Q(rC4[35]), .QN(n3319) );
  DFF_X1 \rC4_reg[34]  ( .D(N237), .CK(mCLK), .Q(rC4[34]), .QN(n3048) );
  DFF_X1 \rC4_reg[33]  ( .D(N236), .CK(mCLK), .Q(rC4[33]), .QN(n3164) );
  DFF_X1 \rC4_reg[32]  ( .D(N235), .CK(mCLK), .Q(rC4[32]), .QN(n3335) );
  DFF_X1 \rC4_reg[31]  ( .D(N234), .CK(mCLK), .Q(rC4[31]), .QN(n3104) );
  DFF_X1 \rC4_reg[30]  ( .D(N233), .CK(mCLK), .Q(rC4[30]), .QN(n3220) );
  DFF_X1 \rC4_reg[29]  ( .D(N232), .CK(mCLK), .Q(rC4[29]), .QN(n3309) );
  DFF_X1 \rC4_reg[28]  ( .D(N231), .CK(mCLK), .Q(rC4[28]), .QN(n3244) );
  DFF_X1 \rC4_reg[27]  ( .D(N230), .CK(mCLK), .Q(rC4[27]), .QN(n3122) );
  DFF_X1 \rC4_reg[26]  ( .D(N229), .CK(mCLK), .Q(rC4[26]), .QN(n3066) );
  DFF_X1 \rC4_reg[25]  ( .D(N228), .CK(mCLK), .Q(rC4[25]), .QN(n3184) );
  DFF_X1 \rC4_reg[24]  ( .D(N227), .CK(mCLK), .Q(rC4[24]), .QN(n3059) );
  DFF_X1 \rC4_reg[23]  ( .D(N226), .CK(mCLK), .Q(rC4[23]), .QN(n3318) );
  DFF_X1 \rC4_reg[22]  ( .D(N225), .CK(mCLK), .Q(rC4[22]), .QN(n3234) );
  DFF_X1 \rC4_reg[21]  ( .D(N224), .CK(mCLK), .Q(rC4[21]), .QN(n3034) );
  DFF_X1 \rC4_reg[20]  ( .D(N223), .CK(mCLK), .Q(rC4[20]), .QN(n3111) );
  DFF_X1 \rC4_reg[19]  ( .D(N222), .CK(mCLK), .Q(rC4[19]), .QN(n3341) );
  DFF_X1 \rC4_reg[18]  ( .D(N221), .CK(mCLK), .Q(rC4[18]), .QN(n3012) );
  DFF_X1 \rC4_reg[17]  ( .D(N220), .CK(mCLK), .Q(rC4[17]), .QN(n3085) );
  DFF_X1 \rC4_reg[16]  ( .D(N219), .CK(mCLK), .Q(rC4[16]), .QN(n3223) );
  DFF_X1 \rC4_reg[15]  ( .D(N218), .CK(mCLK), .Q(rC4[15]), .QN(n3464) );
  DFF_X1 \rC4_reg[14]  ( .D(N217), .CK(mCLK), .Q(rC4[14]), .QN(n3482) );
  DFF_X1 \rC4_reg[13]  ( .D(N216), .CK(mCLK), .Q(rC4[13]), .QN(n3198) );
  DFF_X1 \rC4_reg[12]  ( .D(N215), .CK(mCLK), .Q(rC4[12]), .QN(n3498) );
  DFF_X1 \rC4_reg[11]  ( .D(N214), .CK(mCLK), .Q(rC4[11]), .QN(n3396) );
  DFF_X1 \rC4_reg[10]  ( .D(N213), .CK(mCLK), .Q(rC4[10]), .QN(n3241) );
  DFF_X1 \rC4_reg[9]  ( .D(N212), .CK(mCLK), .Q(rC4[9]), .QN(n3090) );
  DFF_X1 \rC4_reg[8]  ( .D(N211), .CK(mCLK), .Q(rC4[8]) );
  DFF_X1 \rC4_reg[7]  ( .D(N210), .CK(mCLK), .Q(rC4[7]), .QN(n3169) );
  DFF_X1 \rC4_reg[6]  ( .D(N209), .CK(mCLK), .Q(rC4[6]), .QN(n3201) );
  DFF_X1 \rC4_reg[5]  ( .D(N208), .CK(mCLK), .Q(rC4[5]), .QN(n3311) );
  DFF_X1 \rC4_reg[4]  ( .D(N207), .CK(mCLK), .Q(rC4[4]), .QN(n3236) );
  DFF_X1 \rC4_reg[3]  ( .D(N206), .CK(mCLK), .Q(rC4[3]), .QN(n3450) );
  DFF_X1 \rC4_reg[2]  ( .D(N205), .CK(mCLK), .Q(rC4[2]), .QN(n3486) );
  DFF_X1 \rC4_reg[1]  ( .D(N204), .CK(mCLK), .Q(rC4[1]), .QN(n3339) );
  DFF_X1 \rC4_reg[0]  ( .D(N203), .CK(mCLK), .Q(rC4[0]), .QN(n3349) );
  DFF_X1 \rC3_reg[63]  ( .D(N202), .CK(mCLK), .Q(rC3[63]) );
  DFF_X1 \rC3_reg[62]  ( .D(N201), .CK(mCLK), .Q(rC3[62]), .QN(n3080) );
  DFF_X1 \rC3_reg[61]  ( .D(N200), .CK(mCLK), .Q(rC3[61]), .QN(n3141) );
  DFF_X1 \rC3_reg[60]  ( .D(N199), .CK(mCLK), .Q(rC3[60]), .QN(n3011) );
  DFF_X1 \rC3_reg[59]  ( .D(N198), .CK(mCLK), .Q(rC3[59]), .QN(n3083) );
  DFF_X1 \rC3_reg[58]  ( .D(N197), .CK(mCLK), .Q(rC3[58]), .QN(n3305) );
  DFF_X1 \rC3_reg[57]  ( .D(N196), .CK(mCLK), .Q(rC3[57]), .QN(n3137) );
  DFF_X1 \rC3_reg[56]  ( .D(N195), .CK(mCLK), .Q(rC3[56]), .QN(n3044) );
  DFF_X1 \rC3_reg[55]  ( .D(N194), .CK(mCLK), .Q(rC3[55]), .QN(n3155) );
  DFF_X1 \rC3_reg[54]  ( .D(N193), .CK(mCLK), .Q(rC3[54]), .QN(n3325) );
  DFF_X1 \rC3_reg[53]  ( .D(N192), .CK(mCLK), .Q(rC3[53]), .QN(n3145) );
  DFF_X1 \rC3_reg[52]  ( .D(N191), .CK(mCLK), .Q(rC3[52]), .QN(n3030) );
  DFF_X1 \rC3_reg[51]  ( .D(N190), .CK(mCLK), .Q(rC3[51]), .QN(n3320) );
  DFF_X1 \rC3_reg[50]  ( .D(N189), .CK(mCLK), .Q(rC3[50]), .QN(n3065) );
  DFF_X1 \rC3_reg[49]  ( .D(N188), .CK(mCLK), .Q(rC3[49]), .QN(n3019) );
  DFF_X1 \rC3_reg[48]  ( .D(N187), .CK(mCLK), .Q(rC3[48]), .QN(n3102) );
  DFF_X1 \rC3_reg[47]  ( .D(N186), .CK(mCLK), .Q(rC3[47]), .QN(n3314) );
  DFF_X1 \rC3_reg[46]  ( .D(N185), .CK(mCLK), .Q(rC3[46]), .QN(n3232) );
  DFF_X1 \rC3_reg[45]  ( .D(N184), .CK(mCLK), .Q(rC3[45]), .QN(n3165) );
  DFF_X1 \rC3_reg[44]  ( .D(N183), .CK(mCLK), .Q(rC3[44]), .QN(n3221) );
  DFF_X1 \rC3_reg[43]  ( .D(N182), .CK(mCLK), .Q(rC3[43]), .QN(n3068) );
  DFF_X1 \rC3_reg[42]  ( .D(N181), .CK(mCLK), .Q(rC3[42]), .QN(n3312) );
  DFF_X1 \rC3_reg[41]  ( .D(N180), .CK(mCLK), .Q(rC3[41]), .QN(n3143) );
  DFF_X1 \rC3_reg[40]  ( .D(N179), .CK(mCLK), .Q(rC3[40]), .QN(n3028) );
  DFF_X1 \rC3_reg[39]  ( .D(N178), .CK(mCLK), .Q(rC3[39]), .QN(n3069) );
  DFF_X1 \rC3_reg[38]  ( .D(N177), .CK(mCLK), .Q(rC3[38]), .QN(n3040) );
  DFF_X1 \rC3_reg[37]  ( .D(N176), .CK(mCLK), .Q(rC3[37]), .QN(n3153) );
  DFF_X1 \rC3_reg[36]  ( .D(N175), .CK(mCLK), .Q(rC3[36]), .QN(n3075) );
  DFF_X1 \rC3_reg[35]  ( .D(N174), .CK(mCLK), .Q(rC3[35]), .QN(n3209) );
  DFF_X1 \rC3_reg[34]  ( .D(N173), .CK(mCLK), .Q(rC3[34]), .QN(n3298) );
  DFF_X1 \rC3_reg[33]  ( .D(N172), .CK(mCLK), .Q(rC3[33]), .QN(n3136) );
  DFF_X1 \rC3_reg[32]  ( .D(N171), .CK(mCLK), .Q(rC3[32]), .QN(n3043) );
  DFF_X1 \rC3_reg[31]  ( .D(N170), .CK(mCLK), .Q(rC3[31]), .QN(n3154) );
  DFF_X1 \rC3_reg[30]  ( .D(N169), .CK(mCLK), .Q(rC3[30]), .QN(n3324) );
  DFF_X1 \rC3_reg[29]  ( .D(N168), .CK(mCLK), .Q(rC3[29]), .QN(n3144) );
  DFF_X1 \rC3_reg[28]  ( .D(N167), .CK(mCLK), .Q(rC3[28]), .QN(n3029) );
  DFF_X1 \rC3_reg[27]  ( .D(N166), .CK(mCLK), .Q(rC3[27]), .QN(n3007) );
  DFF_X1 \rC3_reg[26]  ( .D(N165), .CK(mCLK), .Q(rC3[26]), .QN(n3168) );
  DFF_X1 \rC3_reg[25]  ( .D(N164), .CK(mCLK), .Q(rC3[25]), .QN(n3321) );
  DFF_X1 \rC3_reg[24]  ( .D(N163), .CK(mCLK), .Q(rC3[24]), .QN(n3076) );
  DFF_X1 \rC3_reg[23]  ( .D(N162), .CK(mCLK), .Q(rC3[23]), .QN(n3210) );
  DFF_X1 \rC3_reg[22]  ( .D(N161), .CK(mCLK), .Q(rC3[22]), .QN(n3329) );
  DFF_X1 \rC3_reg[21]  ( .D(N160), .CK(mCLK), .Q(rC3[21]), .QN(n3202) );
  DFF_X1 \rC3_reg[20]  ( .D(N159), .CK(mCLK), .Q(rC3[20]), .QN(n3093) );
  DFF_X1 \rC3_reg[19]  ( .D(N158), .CK(mCLK), .Q(rC3[19]), .QN(n3256) );
  DFF_X1 \rC3_reg[18]  ( .D(N157), .CK(mCLK), .Q(rC3[18]), .QN(n3013) );
  DFF_X1 \rC3_reg[17]  ( .D(N156), .CK(mCLK), .Q(rC3[17]), .QN(n3084) );
  DFF_X1 \rC3_reg[16]  ( .D(N155), .CK(mCLK), .Q(rC3[16]), .QN(n3306) );
  DFF_X1 \rC3_reg[15]  ( .D(N154), .CK(mCLK), .Q(rC3[15]), .QN(n3416) );
  DFF_X1 \rC3_reg[14]  ( .D(N153), .CK(mCLK), .Q(n3378), .QN(n3447) );
  DFF_X1 \rC3_reg[13]  ( .D(N152), .CK(mCLK), .Q(rC3[13]), .QN(n3211) );
  DFF_X1 \rC3_reg[12]  ( .D(N151), .CK(mCLK), .Q(rC3[12]) );
  DFF_X1 \rC3_reg[11]  ( .D(N150), .CK(mCLK), .Q(rC3[11]), .QN(n3091) );
  DFF_X1 \rC3_reg[10]  ( .D(N149), .CK(mCLK), .Q(rC3[10]), .QN(n3247) );
  DFF_X1 \rC3_reg[9]  ( .D(N148), .CK(mCLK), .Q(rC3[9]), .QN(n3374) );
  DFF_X1 \rC3_reg[8]  ( .D(N147), .CK(mCLK), .Q(rC3[8]), .QN(n3384) );
  DFF_X1 \rC3_reg[7]  ( .D(N146), .CK(mCLK), .Q(rC3[7]), .QN(n3183) );
  DFF_X1 \rC3_reg[6]  ( .D(N145), .CK(mCLK), .Q(rC3[6]), .QN(n3248) );
  DFF_X1 \rC3_reg[5]  ( .D(N144), .CK(mCLK), .Q(rC3[5]), .QN(n3033) );
  DFF_X1 \rC3_reg[4]  ( .D(N143), .CK(mCLK), .Q(rC3[4]), .QN(n3107) );
  DFF_X1 \rC3_reg[3]  ( .D(N142), .CK(mCLK), .Q(rC3[3]), .QN(n3400) );
  DFF_X1 \rC3_reg[2]  ( .D(N141), .CK(mCLK), .Q(rC3[2]), .QN(n3401) );
  DFF_X1 \rC3_reg[1]  ( .D(N140), .CK(mCLK), .Q(rC3[1]), .QN(n3157) );
  DFF_X1 \rC3_reg[0]  ( .D(N139), .CK(mCLK), .Q(rC3[0]), .QN(n3348) );
  DFF_X1 \rC2_reg[63]  ( .D(N136), .CK(mCLK), .Q(rC2[63]), .QN(n3337) );
  DFF_X1 \rC2_reg[62]  ( .D(N135), .CK(mCLK), .Q(rC2[62]), .QN(n3327) );
  DFF_X1 \rC2_reg[61]  ( .D(N134), .CK(mCLK), .Q(rC2[61]), .QN(n3207) );
  DFF_X1 \rC2_reg[60]  ( .D(N133), .CK(mCLK), .Q(rC2[60]), .QN(n3261) );
  DFF_X1 \rC2_reg[59]  ( .D(N132), .CK(mCLK), .Q(rC2[59]), .QN(n3292) );
  DFF_X1 \rC2_reg[58]  ( .D(N131), .CK(mCLK), .Q(rC2[58]), .QN(n3050) );
  DFF_X1 \rC2_reg[57]  ( .D(N130), .CK(mCLK), .Q(rC2[57]), .QN(n3196) );
  DFF_X1 \rC2_reg[56]  ( .D(N129), .CK(mCLK), .Q(rC2[56]), .QN(n3301) );
  DFF_X1 \rC2_reg[55]  ( .D(N128), .CK(mCLK), .Q(rC2[55]), .QN(n3239) );
  DFF_X1 \rC2_reg[54]  ( .D(N127), .CK(mCLK), .Q(rC2[54]), .QN(n3074) );
  DFF_X1 \rC2_reg[53]  ( .D(N126), .CK(mCLK), .Q(rC2[53]), .QN(n3231) );
  DFF_X1 \rC2_reg[52]  ( .D(N125), .CK(mCLK), .Q(rC2[52]), .QN(n3288) );
  DFF_X1 \rC2_reg[51]  ( .D(N124), .CK(mCLK), .Q(rC2[51]), .QN(n3057) );
  DFF_X1 \rC2_reg[50]  ( .D(N123), .CK(mCLK), .Q(rC2[50]), .QN(n3315) );
  DFF_X1 \rC2_reg[49]  ( .D(N122), .CK(mCLK), .Q(rC2[49]), .QN(n3307) );
  DFF_X1 \rC2_reg[48]  ( .D(N121), .CK(mCLK), .Q(rC2[48]), .QN(n3188) );
  DFF_X1 \rC2_reg[47]  ( .D(N120), .CK(mCLK), .Q(rC2[47]), .QN(n3022) );
  DFF_X1 \rC2_reg[46]  ( .D(N119), .CK(mCLK), .Q(rC2[46]), .QN(n3114) );
  DFF_X1 \rC2_reg[45]  ( .D(N118), .CK(mCLK), .Q(rC2[45]), .QN(n3227) );
  DFF_X1 \rC2_reg[44]  ( .D(N117), .CK(mCLK), .Q(rC2[44]), .QN(n3163) );
  DFF_X1 \rC2_reg[43]  ( .D(N116), .CK(mCLK), .Q(rC2[43]), .QN(n3297) );
  DFF_X1 \rC2_reg[42]  ( .D(N115), .CK(mCLK), .Q(rC2[42]), .QN(n3181) );
  DFF_X1 \rC2_reg[41]  ( .D(N114), .CK(mCLK), .Q(rC2[41]), .QN(n3041) );
  DFF_X1 \rC2_reg[40]  ( .D(N113), .CK(mCLK), .Q(rC2[40]), .QN(n3158) );
  DFF_X1 \rC2_reg[39]  ( .D(N112), .CK(mCLK), .Q(rC2[39]), .QN(n3224) );
  DFF_X1 \rC2_reg[38]  ( .D(N111), .CK(mCLK), .Q(rC2[38]), .QN(n3032) );
  DFF_X1 \rC2_reg[37]  ( .D(N110), .CK(mCLK), .Q(rC2[37]), .QN(n3106) );
  DFF_X1 \rC2_reg[36]  ( .D(N109), .CK(mCLK), .Q(rC2[36]), .QN(n3017) );
  DFF_X1 \rC2_reg[35]  ( .D(N108), .CK(mCLK), .Q(rC2[35]), .QN(n3088) );
  DFF_X1 \rC2_reg[34]  ( .D(N107), .CK(mCLK), .Q(rC2[34]), .QN(n3342) );
  DFF_X1 \rC2_reg[33]  ( .D(N106), .CK(mCLK), .Q(rC2[33]), .QN(n3225) );
  DFF_X1 \rC2_reg[32]  ( .D(N105), .CK(mCLK), .Q(rC2[32]), .QN(n3086) );
  DFF_X1 \rC2_reg[31]  ( .D(N104), .CK(mCLK), .Q(rC2[31]), .QN(n3180) );
  DFF_X1 \rC2_reg[30]  ( .D(N103), .CK(mCLK), .Q(rC2[30]), .QN(n3110) );
  DFF_X1 \rC2_reg[29]  ( .D(N102), .CK(mCLK), .Q(rC2[29]), .QN(n3042) );
  DFF_X1 \rC2_reg[28]  ( .D(N101), .CK(mCLK), .Q(rC2[28]), .QN(n3159) );
  DFF_X1 \rC2_reg[27]  ( .D(N100), .CK(mCLK), .Q(rC2[27]), .QN(n3176) );
  DFF_X1 \rC2_reg[26]  ( .D(N99), .CK(mCLK), .Q(rC2[26]), .QN(n3317) );
  DFF_X1 \rC2_reg[25]  ( .D(N98), .CK(mCLK), .Q(rC2[25]), .QN(n3170) );
  DFF_X1 \rC2_reg[24]  ( .D(N97), .CK(mCLK), .Q(rC2[24]), .QN(n3303) );
  DFF_X1 \rC2_reg[23]  ( .D(N96), .CK(mCLK), .Q(rC2[23]), .QN(n3023) );
  DFF_X1 \rC2_reg[22]  ( .D(N95), .CK(mCLK), .Q(rC2[22]), .QN(n3115) );
  DFF_X1 \rC2_reg[21]  ( .D(N94), .CK(mCLK), .Q(rC2[21]), .QN(n3336) );
  DFF_X1 \rC2_reg[20]  ( .D(N93), .CK(mCLK), .Q(rC2[20]), .QN(n3253) );
  DFF_X1 \rC2_reg[19]  ( .D(N92), .CK(mCLK), .Q(rC2[19]), .QN(n3094) );
  DFF_X1 \rC2_reg[18]  ( .D(N91), .CK(mCLK), .Q(rC2[18]), .QN(n3260) );
  DFF_X1 \rC2_reg[17]  ( .D(N90), .CK(mCLK), .Q(rC2[17]), .QN(n3295) );
  DFF_X1 \rC2_reg[16]  ( .D(N89), .CK(mCLK), .Q(rC2[16]), .QN(n3112) );
  DFF_X1 \rC2_reg[15]  ( .D(N88), .CK(mCLK), .Q(rC2[15]), .QN(n3497) );
  DFF_X1 \rC2_reg[14]  ( .D(N87), .CK(mCLK), .Q(n3462), .QN(n3500) );
  DFF_X1 \rC2_reg[13]  ( .D(N86), .CK(mCLK), .Q(rC2[13]), .QN(n3108) );
  DFF_X1 \rC2_reg[12]  ( .D(N85), .CK(mCLK), .Q(rC2[12]), .QN(n3478) );
  DFF_X1 \rC2_reg[11]  ( .D(N84), .CK(mCLK), .Q(n3397), .QN(n3490) );
  DFF_X1 \rC2_reg[10]  ( .D(N83), .CK(mCLK), .Q(rC2[10]), .QN(n3142) );
  DFF_X1 \rC2_reg[9]  ( .D(N82), .CK(mCLK), .Q(rC2[9]), .QN(n3322) );
  DFF_X1 \rC2_reg[8]  ( .D(N81), .CK(mCLK), .Q(rC2[8]), .QN(n3310) );
  DFF_X1 \rC2_reg[7]  ( .D(N80), .CK(mCLK), .Q(rC2[7]), .QN(n3246) );
  DFF_X1 \rC2_reg[6]  ( .D(N79), .CK(mCLK), .Q(rC2[6]), .QN(n3109) );
  DFF_X1 \rC2_reg[5]  ( .D(N78), .CK(mCLK), .Q(rC2[5]), .QN(n3047) );
  DFF_X1 \rC2_reg[4]  ( .D(N77), .CK(mCLK), .Q(rC2[4]), .QN(n3152) );
  DFF_X1 \rC2_reg[3]  ( .D(N76), .CK(mCLK), .Q(rC2[3]), .QN(n3332) );
  DFF_X1 \rC2_reg[2]  ( .D(N75), .CK(mCLK), .Q(rC2[2]), .QN(n3381) );
  DFF_X1 \rC2_reg[1]  ( .D(N74), .CK(mCLK), .Q(rC2[1]), .QN(n3480) );
  DFF_X1 \rC2_reg[0]  ( .D(N73), .CK(mCLK), .Q(rC2[0]), .QN(n3455) );
  DFF_X1 \mY1_reg[63]  ( .D(rC5[63]), .CK(mCLK), .Q(mY1[63]) );
  DFF_X1 \mY1_reg[62]  ( .D(rC5[62]), .CK(mCLK), .Q(mY1[62]) );
  DFF_X1 \mY1_reg[61]  ( .D(rC5[61]), .CK(mCLK), .Q(mY1[61]) );
  DFF_X1 \mY1_reg[60]  ( .D(rC5[60]), .CK(mCLK), .Q(mY1[60]) );
  DFF_X1 \mY1_reg[59]  ( .D(rC5[59]), .CK(mCLK), .Q(mY1[59]) );
  DFF_X1 \mY1_reg[58]  ( .D(rC5[58]), .CK(mCLK), .Q(mY1[58]) );
  DFF_X1 \mY1_reg[57]  ( .D(rC5[57]), .CK(mCLK), .Q(mY1[57]) );
  DFF_X1 \mY1_reg[56]  ( .D(rC5[56]), .CK(mCLK), .Q(mY1[56]) );
  DFF_X1 \mY1_reg[55]  ( .D(rC5[55]), .CK(mCLK), .Q(mY1[55]) );
  DFF_X1 \mY1_reg[54]  ( .D(rC5[54]), .CK(mCLK), .Q(mY1[54]) );
  DFF_X1 \mY1_reg[53]  ( .D(rC5[53]), .CK(mCLK), .Q(mY1[53]) );
  DFF_X1 \mY1_reg[52]  ( .D(rC5[52]), .CK(mCLK), .Q(mY1[52]) );
  DFF_X1 \mY1_reg[51]  ( .D(rC5[51]), .CK(mCLK), .Q(mY1[51]) );
  DFF_X1 \rC5_reg[50]  ( .D(N329), .CK(mCLK), .Q(rC5[50]) );
  DFF_X1 \mY1_reg[50]  ( .D(rC5[50]), .CK(mCLK), .Q(mY1[50]) );
  DFF_X1 \mY1_reg[49]  ( .D(rC5[49]), .CK(mCLK), .Q(mY1[49]) );
  DFF_X1 \mY1_reg[48]  ( .D(rC5[48]), .CK(mCLK), .Q(mY1[48]) );
  DFF_X1 \mY1_reg[47]  ( .D(rC5[47]), .CK(mCLK), .Q(mY1[47]) );
  DFF_X1 \mY1_reg[46]  ( .D(rC5[46]), .CK(mCLK), .Q(mY1[46]) );
  DFF_X1 \mY1_reg[45]  ( .D(rC5[45]), .CK(mCLK), .Q(mY1[45]) );
  DFF_X1 \mY1_reg[44]  ( .D(rC5[44]), .CK(mCLK), .Q(mY1[44]) );
  DFF_X1 \mY1_reg[43]  ( .D(rC5[43]), .CK(mCLK), .Q(mY1[43]) );
  DFF_X1 \mY1_reg[42]  ( .D(rC5[42]), .CK(mCLK), .Q(mY1[42]) );
  DFF_X1 \rC5_reg[41]  ( .D(N320), .CK(mCLK), .Q(rC5[41]) );
  DFF_X1 \mY1_reg[41]  ( .D(rC5[41]), .CK(mCLK), .Q(mY1[41]) );
  DFF_X1 \rC5_reg[40]  ( .D(N319), .CK(mCLK), .Q(rC5[40]) );
  DFF_X1 \mY1_reg[40]  ( .D(rC5[40]), .CK(mCLK), .Q(mY1[40]) );
  DFF_X1 \rC5_reg[39]  ( .D(N318), .CK(mCLK), .Q(rC5[39]) );
  DFF_X1 \mY1_reg[39]  ( .D(rC5[39]), .CK(mCLK), .Q(mY1[39]) );
  DFF_X1 \rC5_reg[38]  ( .D(N317), .CK(mCLK), .Q(rC5[38]) );
  DFF_X1 \mY1_reg[38]  ( .D(rC5[38]), .CK(mCLK), .Q(mY1[38]) );
  DFF_X1 \rC5_reg[37]  ( .D(N316), .CK(mCLK), .Q(rC5[37]) );
  DFF_X1 \mY1_reg[37]  ( .D(rC5[37]), .CK(mCLK), .Q(mY1[37]) );
  DFF_X1 \rC5_reg[36]  ( .D(N315), .CK(mCLK), .Q(rC5[36]) );
  DFF_X1 \mY1_reg[36]  ( .D(rC5[36]), .CK(mCLK), .Q(mY1[36]) );
  DFF_X1 \rC5_reg[35]  ( .D(N314), .CK(mCLK), .Q(rC5[35]) );
  DFF_X1 \mY1_reg[35]  ( .D(rC5[35]), .CK(mCLK), .Q(mY1[35]) );
  DFF_X1 \mY1_reg[34]  ( .D(rC5[34]), .CK(mCLK), .Q(mY1[34]) );
  DFF_X1 \rC5_reg[33]  ( .D(N312), .CK(mCLK), .Q(rC5[33]) );
  DFF_X1 \mY1_reg[33]  ( .D(rC5[33]), .CK(mCLK), .Q(mY1[33]) );
  DFF_X1 \rC5_reg[32]  ( .D(N311), .CK(mCLK), .Q(rC5[32]) );
  DFF_X1 \mY1_reg[32]  ( .D(rC5[32]), .CK(mCLK), .Q(mY1[32]) );
  DFF_X1 \mY1_reg[31]  ( .D(rC5[31]), .CK(mCLK), .Q(mY1[31]) );
  DFF_X1 \rC5_reg[30]  ( .D(N309), .CK(mCLK), .Q(rC5[30]) );
  DFF_X1 \mY1_reg[30]  ( .D(rC5[30]), .CK(mCLK), .Q(mY1[30]) );
  DFF_X1 \rC5_reg[29]  ( .D(N308), .CK(mCLK), .Q(rC5[29]) );
  DFF_X1 \mY1_reg[29]  ( .D(rC5[29]), .CK(mCLK), .Q(mY1[29]) );
  DFF_X1 \rC5_reg[28]  ( .D(N307), .CK(mCLK), .Q(rC5[28]) );
  DFF_X1 \mY1_reg[28]  ( .D(rC5[28]), .CK(mCLK), .Q(mY1[28]) );
  DFF_X1 \rC5_reg[27]  ( .D(N306), .CK(mCLK), .Q(rC5[27]) );
  DFF_X1 \mY1_reg[27]  ( .D(rC5[27]), .CK(mCLK), .Q(mY1[27]) );
  DFF_X1 \rC5_reg[26]  ( .D(N305), .CK(mCLK), .Q(rC5[26]) );
  DFF_X1 \mY1_reg[26]  ( .D(rC5[26]), .CK(mCLK), .Q(mY1[26]) );
  DFF_X1 \rC5_reg[25]  ( .D(N304), .CK(mCLK), .Q(rC5[25]) );
  DFF_X1 \mY1_reg[25]  ( .D(rC5[25]), .CK(mCLK), .Q(mY1[25]) );
  DFF_X1 \rC5_reg[24]  ( .D(N303), .CK(mCLK), .Q(rC5[24]) );
  DFF_X1 \mY1_reg[24]  ( .D(rC5[24]), .CK(mCLK), .Q(mY1[24]) );
  DFF_X1 \rC5_reg[23]  ( .D(N302), .CK(mCLK), .Q(rC5[23]) );
  DFF_X1 \mY1_reg[23]  ( .D(rC5[23]), .CK(mCLK), .Q(mY1[23]) );
  DFF_X1 \rC5_reg[22]  ( .D(N301), .CK(mCLK), .Q(rC5[22]) );
  DFF_X1 \mY1_reg[22]  ( .D(rC5[22]), .CK(mCLK), .Q(mY1[22]) );
  DFF_X1 \rC5_reg[21]  ( .D(N300), .CK(mCLK), .Q(rC5[21]) );
  DFF_X1 \mY1_reg[21]  ( .D(rC5[21]), .CK(mCLK), .Q(mY1[21]) );
  DFF_X1 \mY1_reg[20]  ( .D(rC5[20]), .CK(mCLK), .Q(mY1[20]) );
  DFF_X1 \mY1_reg[19]  ( .D(rC5[19]), .CK(mCLK), .Q(mY1[19]) );
  DFF_X1 \mY1_reg[18]  ( .D(rC5[18]), .CK(mCLK), .Q(mY1[18]) );
  DFF_X1 \rC5_reg[17]  ( .D(N296), .CK(mCLK), .Q(rC5[17]) );
  DFF_X1 \mY1_reg[17]  ( .D(rC5[17]), .CK(mCLK), .Q(mY1[17]) );
  DFF_X1 \rC5_reg[16]  ( .D(N295), .CK(mCLK), .Q(rC5[16]) );
  DFF_X1 \mY1_reg[16]  ( .D(rC5[16]), .CK(mCLK), .Q(mY1[16]) );
  DFF_X1 \mY1_reg[15]  ( .D(rC5[15]), .CK(mCLK), .Q(mY1[15]) );
  DFF_X1 \mY1_reg[14]  ( .D(rC5[14]), .CK(mCLK), .Q(mY1[14]) );
  DFF_X1 \mY1_reg[13]  ( .D(rC5[13]), .CK(mCLK), .Q(mY1[13]) );
  DFF_X1 \mY1_reg[12]  ( .D(rC5[12]), .CK(mCLK), .Q(mY1[12]) );
  DFF_X1 \rC5_reg[11]  ( .D(N290), .CK(mCLK), .Q(rC5[11]) );
  DFF_X1 \mY1_reg[11]  ( .D(rC5[11]), .CK(mCLK), .Q(mY1[11]) );
  DFF_X1 \mY1_reg[10]  ( .D(rC5[10]), .CK(mCLK), .Q(mY1[10]) );
  DFF_X1 \mY1_reg[9]  ( .D(rC5[9]), .CK(mCLK), .Q(mY1[9]) );
  DFF_X1 \mY1_reg[8]  ( .D(rC5[8]), .CK(mCLK), .Q(mY1[8]) );
  DFF_X1 \mY1_reg[7]  ( .D(rC5[7]), .CK(mCLK), .Q(mY1[7]) );
  DFF_X1 \mY1_reg[6]  ( .D(rC5[6]), .CK(mCLK), .Q(mY1[6]) );
  DFF_X1 \mY1_reg[5]  ( .D(rC5[5]), .CK(mCLK), .Q(mY1[5]) );
  DFF_X1 \rC5_reg[4]  ( .D(N283), .CK(mCLK), .Q(rC5[4]) );
  DFF_X1 \mY1_reg[4]  ( .D(rC5[4]), .CK(mCLK), .Q(mY1[4]) );
  DFF_X1 \mY1_reg[3]  ( .D(rC5[3]), .CK(mCLK), .Q(mY1[3]) );
  DFF_X1 \rC5_reg[2]  ( .D(N281), .CK(mCLK), .Q(rC5[2]) );
  DFF_X1 \mY1_reg[2]  ( .D(rC5[2]), .CK(mCLK), .Q(mY1[2]) );
  DFF_X1 \rC5_reg[1]  ( .D(N280), .CK(mCLK), .Q(rC5[1]) );
  DFF_X1 \mY1_reg[1]  ( .D(rC5[1]), .CK(mCLK), .Q(mY1[1]) );
  DFF_X1 \mY1_reg[0]  ( .D(rC5[0]), .CK(mCLK), .Q(mY1[0]) );
  DFF_X1 \rC7_reg[63]  ( .D(N470), .CK(mCLK), .Q(rC7[63]), .QN(n3116) );
  DFF_X1 \rC7_reg[62]  ( .D(N469), .CK(mCLK), .Q(rC7[62]), .QN(n3264) );
  DFF_X1 \rC7_reg[51]  ( .D(N458), .CK(mCLK), .Q(rC7[51]), .QN(n3250) );
  DFF_X1 \rC7_reg[50]  ( .D(N457), .CK(mCLK), .Q(rC7[50]), .QN(n3281) );
  DFF_X1 \rC7_reg[49]  ( .D(N456), .CK(mCLK), .Q(rC7[49]), .QN(n3096) );
  DFF_X1 \rC7_reg[48]  ( .D(N455), .CK(mCLK), .Q(rC7[48]), .QN(n3199) );
  DFF_X1 \rC7_reg[47]  ( .D(N454), .CK(mCLK), .Q(rC7[47]), .QN(n3269) );
  DFF_X1 \rC7_reg[46]  ( .D(N453), .CK(mCLK), .Q(rC7[46]), .QN(n3212) );
  DFF_X1 \rC7_reg[45]  ( .D(N452), .CK(mCLK), .Q(rC7[45]), .QN(n3251) );
  DFF_X1 \rC7_reg[44]  ( .D(N451), .CK(mCLK), .Q(rC7[44]), .QN(n3282) );
  DFF_X1 \rC7_reg[42]  ( .D(N449), .CK(mCLK), .Q(rC7[42]), .QN(n3200) );
  DFF_X1 \rC7_reg[41]  ( .D(N448), .CK(mCLK), .Q(rC7[41]), .QN(n3270) );
  DFF_X1 \rC7_reg[40]  ( .D(N447), .CK(mCLK), .Q(rC7[40]), .QN(n3205) );
  DFF_X1 \rC7_reg[39]  ( .D(N446), .CK(mCLK), .Q(rC7[39]), .QN(n3062) );
  DFF_X1 \rC7_reg[35]  ( .D(N442), .CK(mCLK), .Q(rC7[35]), .QN(n3273) );
  DFF_X1 \rC7_reg[34]  ( .D(N441), .CK(mCLK), .Q(rC7[34]), .QN(n3283) );
  DFF_X1 \rC7_reg[33]  ( .D(N440), .CK(mCLK), .Q(rC7[33]), .QN(n3089) );
  DFF_X1 \rC7_reg[32]  ( .D(N439), .CK(mCLK), .Q(rC7[32]), .QN(n3009) );
  DFF_X1 \rC7_reg[31]  ( .D(N438), .CK(mCLK), .Q(rC7[31]), .QN(n3126) );
  DFF_X1 \rC7_reg[30]  ( .D(N437), .CK(mCLK), .Q(rC7[30]), .QN(n3276) );
  DFF_X1 \rC7_reg[29]  ( .D(N436), .CK(mCLK), .Q(rC7[29]), .QN(n3119) );
  DFF_X1 \rC7_reg[13]  ( .D(N420), .CK(mCLK), .Q(rC7[13]), .QN(n3403) );
  DFF_X1 \rC7_reg[11]  ( .D(N418), .CK(mCLK), .Q(rC7[11]), .QN(n3686) );
  DFF_X1 \rC7_reg[10]  ( .D(N417), .CK(mCLK), .Q(rC7[10]), .QN(n3186) );
  DFF_X1 \rC7_reg[9]  ( .D(N416), .CK(mCLK), .Q(rC7[9]), .QN(n3064) );
  DFF_X1 \rC7_reg[2]  ( .D(N409), .CK(mCLK), .Q(rC7[2]), .QN(n3687) );
  DFF_X1 \rC6_reg[63]  ( .D(N406), .CK(mCLK), .Q(rC6[63]), .QN(n3192) );
  DFF_X1 \rC6_reg[62]  ( .D(N405), .CK(mCLK), .Q(rC6[62]), .QN(n3053) );
  DFF_X1 \rC6_reg[61]  ( .D(N404), .CK(mCLK), .Q(rC6[61]), .QN(n3038) );
  DFF_X1 \rC6_reg[60]  ( .D(N403), .CK(mCLK), .Q(rC6[60]), .QN(n3128) );
  DFF_X1 \rC6_reg[59]  ( .D(N402), .CK(mCLK), .Q(rC6[59]), .QN(n3203) );
  DFF_X1 \rC6_reg[58]  ( .D(N401), .CK(mCLK), .Q(rC6[58]), .QN(n3125) );
  DFF_X1 \rC6_reg[57]  ( .D(N400), .CK(mCLK), .Q(rC6[57]), .QN(n3024) );
  DFF_X1 \rC6_reg[56]  ( .D(N399), .CK(mCLK), .Q(rC6[56]), .QN(n3123) );
  DFF_X1 \rC6_reg[55]  ( .D(N398), .CK(mCLK), .Q(rC6[55]), .QN(n3213) );
  DFF_X1 \rC6_reg[54]  ( .D(N397), .CK(mCLK), .Q(rC6[54]), .QN(n3135) );
  DFF_X1 \rC6_reg[53]  ( .D(N396), .CK(mCLK), .Q(rC6[53]), .QN(n3280) );
  DFF_X1 \rC6_reg[52]  ( .D(N395), .CK(mCLK), .Q(rC6[52]), .QN(n3175) );
  DFF_X1 \rC6_reg[51]  ( .D(N394), .CK(mCLK), .Q(rC6[51]), .QN(n3160) );
  DFF_X1 \rC6_reg[50]  ( .D(N393), .CK(mCLK), .Q(rC6[50]), .QN(n3027) );
  DFF_X1 \rC6_reg[49]  ( .D(N392), .CK(mCLK), .Q(rC6[49]), .QN(n3173) );
  DFF_X1 \rC6_reg[48]  ( .D(N391), .CK(mCLK), .Q(rC6[48]), .QN(n3100) );
  DFF_X1 \rC6_reg[47]  ( .D(N390), .CK(mCLK), .Q(rC6[47]), .QN(n3035) );
  DFF_X1 \rC6_reg[46]  ( .D(N389), .CK(mCLK), .Q(rC6[46]), .QN(n3124) );
  DFF_X1 \rC6_reg[45]  ( .D(N388), .CK(mCLK), .Q(rC6[45]), .QN(n3161) );
  DFF_X1 \rC6_reg[44]  ( .D(N387), .CK(mCLK), .Q(rC6[44]), .QN(n3039) );
  DFF_X1 \rC6_reg[43]  ( .D(N386), .CK(mCLK), .Q(rC6[43]), .QN(n3174) );
  DFF_X1 \rC6_reg[42]  ( .D(N385), .CK(mCLK), .Q(rC6[42]), .QN(n3101) );
  DFF_X1 \rC6_reg[41]  ( .D(N384), .CK(mCLK), .Q(rC6[41]), .QN(n3036) );
  DFF_X1 \rC6_reg[40]  ( .D(N383), .CK(mCLK), .Q(rC6[40]), .QN(n3129) );
  DFF_X1 \rC6_reg[39]  ( .D(N382), .CK(mCLK), .Q(rC6[39]), .QN(n3265) );
  DFF_X1 \rC6_reg[38]  ( .D(N381), .CK(mCLK), .Q(rC6[38]), .QN(n3271) );
  DFF_X1 \rC6_reg[37]  ( .D(N380), .CK(mCLK), .Q(rC6[37]), .QN(n3219) );
  DFF_X1 \rC6_reg[36]  ( .D(N379), .CK(mCLK), .Q(rC6[36]), .QN(n3267) );
  DFF_X1 \rC6_reg[35]  ( .D(N378), .CK(mCLK), .Q(rC6[35]), .QN(n3060) );
  DFF_X1 \rC6_reg[34]  ( .D(N377), .CK(mCLK), .Q(rC6[34]), .QN(n3015) );
  DFF_X1 \rC6_reg[33]  ( .D(N376), .CK(mCLK), .Q(rC6[33]), .QN(n3179) );
  DFF_X1 \rC6_reg[32]  ( .D(N375), .CK(mCLK), .Q(rC6[32]), .QN(n3257) );
  DFF_X1 \rC6_reg[31]  ( .D(N374), .CK(mCLK), .Q(rC6[31]), .QN(n3214) );
  DFF_X1 \rC6_reg[30]  ( .D(N373), .CK(mCLK), .Q(rC6[30]), .QN(n3063) );
  DFF_X1 \rC6_reg[29]  ( .D(N372), .CK(mCLK), .Q(rC6[29]), .QN(n3208) );
  DFF_X1 \rC6_reg[28]  ( .D(N371), .CK(mCLK), .Q(rC6[28]), .QN(n3278) );
  DFF_X1 \rC6_reg[27]  ( .D(N370), .CK(mCLK), .Q(rC6[27]), .QN(n3148) );
  DFF_X1 \rC6_reg[26]  ( .D(N369), .CK(mCLK), .Q(rC6[26]), .QN(n3025) );
  DFF_X1 \rC6_reg[25]  ( .D(N368), .CK(mCLK), .Q(rC6[25]), .QN(n3071) );
  DFF_X1 \rC6_reg[24]  ( .D(N367), .CK(mCLK), .Q(rC6[24]), .QN(n3266) );
  DFF_X1 \rC6_reg[23]  ( .D(N366), .CK(mCLK), .Q(rC6[23]), .QN(n3061) );
  DFF_X1 \rC6_reg[22]  ( .D(N365), .CK(mCLK), .Q(rC6[22]), .QN(n3016) );
  DFF_X1 \rC6_reg[21]  ( .D(N364), .CK(mCLK), .Q(rC6[21]), .QN(n3117) );
  DFF_X1 \rC6_reg[20]  ( .D(N363), .CK(mCLK), .Q(rC6[20]), .QN(n3285) );
  DFF_X1 \rC6_reg[19]  ( .D(N362), .CK(mCLK), .Q(rC6[19]), .QN(n3132) );
  DFF_X1 \rC6_reg[18]  ( .D(N361), .CK(mCLK), .Q(rC6[18]), .QN(n3099) );
  DFF_X1 \rC6_reg[17]  ( .D(N360), .CK(mCLK), .Q(rC6[17]), .QN(n3046) );
  DFF_X1 \rC6_reg[16]  ( .D(N359), .CK(mCLK), .Q(rC6[16]), .QN(n3127) );
  DFF_X1 \rC6_reg[15]  ( .D(N358), .CK(mCLK), .Q(rC6[15]), .QN(n3258) );
  DFF_X1 \rC6_reg[14]  ( .D(N357), .CK(mCLK), .Q(rC6[14]), .QN(n3182) );
  DFF_X1 \rC6_reg[13]  ( .D(N356), .CK(mCLK), .Q(rC6[13]), .QN(n3284) );
  DFF_X1 \rC6_reg[12]  ( .D(N355), .CK(mCLK), .Q(rC6[12]), .QN(n3402) );
  DFF_X1 \rC6_reg[11]  ( .D(N354), .CK(mCLK), .Q(rC6[11]), .QN(n3678) );
  DFF_X1 \rC6_reg[10]  ( .D(N353), .CK(mCLK), .Q(rC6[10]), .QN(n3677) );
  DFF_X1 \rC6_reg[9]  ( .D(N352), .CK(mCLK), .Q(rC6[9]), .QN(n3277) );
  DFF_X1 \rC6_reg[8]  ( .D(N351), .CK(mCLK), .Q(rC6[8]), .QN(n3120) );
  DFF_X1 \rC6_reg[7]  ( .D(N350), .CK(mCLK), .Q(rC6[7]), .QN(n3095) );
  DFF_X1 \rC6_reg[6]  ( .D(N349), .CK(mCLK), .Q(rC6[6]), .QN(n3058) );
  DFF_X1 \rC6_reg[5]  ( .D(N348), .CK(mCLK), .Q(rC6[5]), .QN(n3674) );
  DFF_X1 \rC6_reg[4]  ( .D(N347), .CK(mCLK), .Q(rC6[4]), .QN(n3131) );
  DFF_X1 \rC6_reg[3]  ( .D(N346), .CK(mCLK), .Q(rC6[3]), .QN(n3679) );
  DFF_X1 \rC6_reg[2]  ( .D(N345), .CK(mCLK), .Q(rC6[2]), .QN(n3681) );
  DFF_X1 \rC6_reg[1]  ( .D(N344), .CK(mCLK), .Q(rC6[1]), .QN(n3676) );
  DFF_X1 \rC6_reg[0]  ( .D(N343), .CK(mCLK), .Q(rC6[0]), .QN(n3683) );
  DFF_X1 \mY3_reg[63]  ( .D(N664), .CK(mCLK), .Q(mY3[63]) );
  DFF_X1 \mY3_reg[7]  ( .D(N608), .CK(mCLK), .Q(mY3[7]) );
  DFF_X1 \mY3_reg[6]  ( .D(N607), .CK(mCLK), .Q(mY3[6]) );
  DFF_X1 \mY3_reg[5]  ( .D(N606), .CK(mCLK), .Q(mY3[5]) );
  DFF_X1 \mY2_reg[48]  ( .D(N585), .CK(mCLK), .Q(mY2[48]) );
  DFF_X1 \mY2_reg[23]  ( .D(N560), .CK(mCLK), .Q(mY2[23]) );
  DFF_X1 \mY2_reg[22]  ( .D(N559), .CK(mCLK), .Q(mY2[22]) );
  DFF_X1 \mY2_reg[21]  ( .D(N558), .CK(mCLK), .Q(mY2[21]) );
  DFF_X1 \mY2_reg[11]  ( .D(N548), .CK(mCLK), .Q(mY2[11]) );
  DFF_X1 \mY2_reg[10]  ( .D(N547), .CK(mCLK), .Q(mY2[10]) );
  DFF_X1 \mY2_reg[9]  ( .D(N546), .CK(mCLK), .Q(mY2[9]) );
  DFF_X1 \mY2_reg[8]  ( .D(N545), .CK(mCLK), .Q(mY2[8]) );
  DFF_X1 \mY2_reg[7]  ( .D(N544), .CK(mCLK), .Q(mY2[7]) );
  DFF_X1 \mY2_reg[6]  ( .D(N543), .CK(mCLK), .Q(mY2[6]) );
  DFF_X1 \mY2_reg[5]  ( .D(N542), .CK(mCLK), .Q(mY2[5]) );
  DFF_X1 \mY2_reg[4]  ( .D(N541), .CK(mCLK), .Q(mY2[4]) );
  DFF_X1 \mY2_reg[3]  ( .D(N540), .CK(mCLK), .Q(mY2[3]) );
  DFF_X1 \mY2_reg[2]  ( .D(N539), .CK(mCLK), .Q(mY2[2]) );
  DFF_X1 \mY2_reg[1]  ( .D(N538), .CK(mCLK), .Q(mY2[1]) );
  DFF_X1 \mY2_reg[0]  ( .D(N537), .CK(mCLK), .Q(mY2[0]) );
  DFF_X1 \rC8_reg[63]  ( .D(N534), .CK(mCLK), .Q(rC8[63]) );
  DFF_X1 \mY4_reg[63]  ( .D(rC8[63]), .CK(mCLK), .Q(mY4[63]) );
  DFF_X1 \rC8_reg[62]  ( .D(N533), .CK(mCLK), .Q(rC8[62]) );
  DFF_X1 \mY4_reg[62]  ( .D(rC8[62]), .CK(mCLK), .Q(mY4[62]) );
  DFF_X1 \rC8_reg[61]  ( .D(N532), .CK(mCLK), .Q(rC8[61]) );
  DFF_X1 \mY4_reg[61]  ( .D(rC8[61]), .CK(mCLK), .Q(mY4[61]) );
  DFF_X1 \rC8_reg[60]  ( .D(N531), .CK(mCLK), .Q(rC8[60]) );
  DFF_X1 \mY4_reg[60]  ( .D(rC8[60]), .CK(mCLK), .Q(mY4[60]) );
  DFF_X1 \rC8_reg[59]  ( .D(N530), .CK(mCLK), .Q(rC8[59]) );
  DFF_X1 \mY4_reg[59]  ( .D(rC8[59]), .CK(mCLK), .Q(mY4[59]) );
  DFF_X1 \mY4_reg[58]  ( .D(rC8[58]), .CK(mCLK), .Q(mY4[58]) );
  DFF_X1 \rC8_reg[57]  ( .D(N528), .CK(mCLK), .Q(rC8[57]) );
  DFF_X1 \mY4_reg[57]  ( .D(rC8[57]), .CK(mCLK), .Q(mY4[57]) );
  DFF_X1 \mY4_reg[56]  ( .D(rC8[56]), .CK(mCLK), .Q(mY4[56]) );
  DFF_X1 \rC8_reg[55]  ( .D(N526), .CK(mCLK), .Q(rC8[55]) );
  DFF_X1 \mY4_reg[55]  ( .D(rC8[55]), .CK(mCLK), .Q(mY4[55]) );
  DFF_X1 \rC8_reg[54]  ( .D(N525), .CK(mCLK), .Q(rC8[54]) );
  DFF_X1 \mY4_reg[54]  ( .D(rC8[54]), .CK(mCLK), .Q(mY4[54]) );
  DFF_X1 \rC8_reg[53]  ( .D(N524), .CK(mCLK), .Q(rC8[53]) );
  DFF_X1 \mY4_reg[53]  ( .D(rC8[53]), .CK(mCLK), .Q(mY4[53]) );
  DFF_X1 \rC8_reg[52]  ( .D(N523), .CK(mCLK), .Q(rC8[52]) );
  DFF_X1 \mY4_reg[52]  ( .D(rC8[52]), .CK(mCLK), .Q(mY4[52]) );
  DFF_X1 \rC8_reg[51]  ( .D(N522), .CK(mCLK), .Q(rC8[51]) );
  DFF_X1 \mY4_reg[51]  ( .D(rC8[51]), .CK(mCLK), .Q(mY4[51]) );
  DFF_X1 \rC8_reg[50]  ( .D(N521), .CK(mCLK), .Q(rC8[50]) );
  DFF_X1 \mY4_reg[50]  ( .D(rC8[50]), .CK(mCLK), .Q(mY4[50]) );
  DFF_X1 \rC8_reg[49]  ( .D(N520), .CK(mCLK), .Q(rC8[49]) );
  DFF_X1 \mY4_reg[49]  ( .D(rC8[49]), .CK(mCLK), .Q(mY4[49]) );
  DFF_X1 \rC8_reg[48]  ( .D(N519), .CK(mCLK), .Q(rC8[48]) );
  DFF_X1 \mY4_reg[48]  ( .D(rC8[48]), .CK(mCLK), .Q(mY4[48]) );
  DFF_X1 \rC8_reg[47]  ( .D(N518), .CK(mCLK), .Q(rC8[47]) );
  DFF_X1 \mY4_reg[47]  ( .D(rC8[47]), .CK(mCLK), .Q(mY4[47]) );
  DFF_X1 \rC8_reg[46]  ( .D(N517), .CK(mCLK), .Q(rC8[46]) );
  DFF_X1 \mY4_reg[46]  ( .D(rC8[46]), .CK(mCLK), .Q(mY4[46]) );
  DFF_X1 \rC8_reg[45]  ( .D(N516), .CK(mCLK), .Q(rC8[45]) );
  DFF_X1 \mY4_reg[45]  ( .D(rC8[45]), .CK(mCLK), .Q(mY4[45]) );
  DFF_X1 \rC8_reg[44]  ( .D(N515), .CK(mCLK), .Q(rC8[44]) );
  DFF_X1 \mY4_reg[44]  ( .D(rC8[44]), .CK(mCLK), .Q(mY4[44]) );
  DFF_X1 \rC8_reg[43]  ( .D(N514), .CK(mCLK), .Q(rC8[43]) );
  DFF_X1 \mY4_reg[43]  ( .D(rC8[43]), .CK(mCLK), .Q(mY4[43]) );
  DFF_X1 \rC8_reg[42]  ( .D(N513), .CK(mCLK), .Q(rC8[42]) );
  DFF_X1 \mY4_reg[42]  ( .D(rC8[42]), .CK(mCLK), .Q(mY4[42]) );
  DFF_X1 \rC8_reg[41]  ( .D(N512), .CK(mCLK), .Q(rC8[41]) );
  DFF_X1 \mY4_reg[41]  ( .D(rC8[41]), .CK(mCLK), .Q(mY4[41]) );
  DFF_X1 \rC8_reg[40]  ( .D(N511), .CK(mCLK), .Q(rC8[40]) );
  DFF_X1 \mY4_reg[40]  ( .D(rC8[40]), .CK(mCLK), .Q(mY4[40]) );
  DFF_X1 \rC8_reg[39]  ( .D(N510), .CK(mCLK), .Q(rC8[39]) );
  DFF_X1 \mY4_reg[39]  ( .D(rC8[39]), .CK(mCLK), .Q(mY4[39]) );
  DFF_X1 \mY4_reg[38]  ( .D(rC8[38]), .CK(mCLK), .Q(mY4[38]) );
  DFF_X1 \mY4_reg[37]  ( .D(rC8[37]), .CK(mCLK), .Q(mY4[37]) );
  DFF_X1 \rC8_reg[36]  ( .D(N507), .CK(mCLK), .Q(rC8[36]) );
  DFF_X1 \mY4_reg[36]  ( .D(rC8[36]), .CK(mCLK), .Q(mY4[36]) );
  DFF_X1 \mY4_reg[35]  ( .D(rC8[35]), .CK(mCLK), .Q(mY4[35]) );
  DFF_X1 \rC8_reg[34]  ( .D(N505), .CK(mCLK), .Q(rC8[34]) );
  DFF_X1 \mY4_reg[34]  ( .D(rC8[34]), .CK(mCLK), .Q(mY4[34]) );
  DFF_X1 \mY4_reg[33]  ( .D(rC8[33]), .CK(mCLK), .Q(mY4[33]) );
  DFF_X1 \rC8_reg[32]  ( .D(N503), .CK(mCLK), .Q(rC8[32]) );
  DFF_X1 \mY4_reg[32]  ( .D(rC8[32]), .CK(mCLK), .Q(mY4[32]) );
  DFF_X1 \rC8_reg[31]  ( .D(N502), .CK(mCLK), .Q(rC8[31]) );
  DFF_X1 \mY4_reg[31]  ( .D(rC8[31]), .CK(mCLK), .Q(mY4[31]) );
  DFF_X1 \rC8_reg[30]  ( .D(N501), .CK(mCLK), .Q(rC8[30]) );
  DFF_X1 \mY4_reg[30]  ( .D(rC8[30]), .CK(mCLK), .Q(mY4[30]) );
  DFF_X1 \rC8_reg[29]  ( .D(N500), .CK(mCLK), .Q(rC8[29]) );
  DFF_X1 \mY4_reg[29]  ( .D(rC8[29]), .CK(mCLK), .Q(mY4[29]) );
  DFF_X1 \rC8_reg[28]  ( .D(N499), .CK(mCLK), .Q(rC8[28]) );
  DFF_X1 \mY4_reg[28]  ( .D(rC8[28]), .CK(mCLK), .Q(mY4[28]) );
  DFF_X1 \rC8_reg[27]  ( .D(N498), .CK(mCLK), .Q(rC8[27]) );
  DFF_X1 \mY4_reg[27]  ( .D(rC8[27]), .CK(mCLK), .Q(mY4[27]) );
  DFF_X1 \rC8_reg[26]  ( .D(N497), .CK(mCLK), .Q(rC8[26]) );
  DFF_X1 \mY4_reg[26]  ( .D(rC8[26]), .CK(mCLK), .Q(mY4[26]) );
  DFF_X1 \rC8_reg[25]  ( .D(N496), .CK(mCLK), .Q(rC8[25]) );
  DFF_X1 \mY4_reg[25]  ( .D(rC8[25]), .CK(mCLK), .Q(mY4[25]) );
  DFF_X1 \rC8_reg[24]  ( .D(N495), .CK(mCLK), .Q(rC8[24]) );
  DFF_X1 \mY4_reg[24]  ( .D(rC8[24]), .CK(mCLK), .Q(mY4[24]) );
  DFF_X1 \rC8_reg[23]  ( .D(N494), .CK(mCLK), .Q(rC8[23]) );
  DFF_X1 \mY4_reg[23]  ( .D(rC8[23]), .CK(mCLK), .Q(mY4[23]) );
  DFF_X1 \rC8_reg[22]  ( .D(N493), .CK(mCLK), .Q(rC8[22]) );
  DFF_X1 \mY4_reg[22]  ( .D(rC8[22]), .CK(mCLK), .Q(mY4[22]) );
  DFF_X1 \rC8_reg[21]  ( .D(N492), .CK(mCLK), .Q(rC8[21]) );
  DFF_X1 \mY4_reg[21]  ( .D(rC8[21]), .CK(mCLK), .Q(mY4[21]) );
  DFF_X1 \rC8_reg[20]  ( .D(N491), .CK(mCLK), .Q(rC8[20]) );
  DFF_X1 \mY4_reg[20]  ( .D(rC8[20]), .CK(mCLK), .Q(mY4[20]) );
  DFF_X1 \rC8_reg[19]  ( .D(N490), .CK(mCLK), .Q(rC8[19]) );
  DFF_X1 \mY4_reg[19]  ( .D(rC8[19]), .CK(mCLK), .Q(mY4[19]) );
  DFF_X1 \rC8_reg[18]  ( .D(N489), .CK(mCLK), .Q(rC8[18]) );
  DFF_X1 \mY4_reg[18]  ( .D(rC8[18]), .CK(mCLK), .Q(mY4[18]) );
  DFF_X1 \rC8_reg[17]  ( .D(N488), .CK(mCLK), .Q(rC8[17]) );
  DFF_X1 \mY4_reg[17]  ( .D(rC8[17]), .CK(mCLK), .Q(mY4[17]) );
  DFF_X1 \rC8_reg[16]  ( .D(N487), .CK(mCLK), .Q(rC8[16]) );
  DFF_X1 \mY4_reg[16]  ( .D(rC8[16]), .CK(mCLK), .Q(mY4[16]) );
  DFF_X1 \rC8_reg[15]  ( .D(N486), .CK(mCLK), .Q(rC8[15]) );
  DFF_X1 \mY4_reg[15]  ( .D(rC8[15]), .CK(mCLK), .Q(mY4[15]) );
  DFF_X1 \rC8_reg[14]  ( .D(N485), .CK(mCLK), .Q(rC8[14]) );
  DFF_X1 \mY4_reg[14]  ( .D(rC8[14]), .CK(mCLK), .Q(mY4[14]) );
  DFF_X1 \rC8_reg[13]  ( .D(N484), .CK(mCLK), .Q(rC8[13]) );
  DFF_X1 \mY4_reg[13]  ( .D(rC8[13]), .CK(mCLK), .Q(mY4[13]) );
  DFF_X1 \rC8_reg[12]  ( .D(N483), .CK(mCLK), .Q(rC8[12]) );
  DFF_X1 \mY4_reg[12]  ( .D(rC8[12]), .CK(mCLK), .Q(mY4[12]) );
  DFF_X1 \rC8_reg[11]  ( .D(N482), .CK(mCLK), .Q(rC8[11]) );
  DFF_X1 \mY4_reg[11]  ( .D(rC8[11]), .CK(mCLK), .Q(mY4[11]) );
  DFF_X1 \rC8_reg[10]  ( .D(N481), .CK(mCLK), .Q(rC8[10]) );
  DFF_X1 \mY4_reg[10]  ( .D(rC8[10]), .CK(mCLK), .Q(mY4[10]) );
  DFF_X1 \rC8_reg[9]  ( .D(N480), .CK(mCLK), .Q(rC8[9]) );
  DFF_X1 \mY4_reg[9]  ( .D(rC8[9]), .CK(mCLK), .Q(mY4[9]) );
  DFF_X1 \rC8_reg[8]  ( .D(N479), .CK(mCLK), .Q(rC8[8]) );
  DFF_X1 \mY4_reg[8]  ( .D(rC8[8]), .CK(mCLK), .Q(mY4[8]) );
  DFF_X1 \rC8_reg[7]  ( .D(N478), .CK(mCLK), .Q(rC8[7]) );
  DFF_X1 \mY4_reg[7]  ( .D(rC8[7]), .CK(mCLK), .Q(mY4[7]) );
  DFF_X1 \rC8_reg[6]  ( .D(N477), .CK(mCLK), .Q(rC8[6]) );
  DFF_X1 \mY4_reg[6]  ( .D(rC8[6]), .CK(mCLK), .Q(mY4[6]) );
  DFF_X1 \rC8_reg[5]  ( .D(N476), .CK(mCLK), .Q(rC8[5]) );
  DFF_X1 \mY4_reg[5]  ( .D(rC8[5]), .CK(mCLK), .Q(mY4[5]) );
  DFF_X1 \rC8_reg[4]  ( .D(N475), .CK(mCLK), .Q(rC8[4]) );
  DFF_X1 \mY4_reg[4]  ( .D(rC8[4]), .CK(mCLK), .Q(mY4[4]) );
  DFF_X1 \rC8_reg[3]  ( .D(N474), .CK(mCLK), .Q(rC8[3]) );
  DFF_X1 \mY4_reg[3]  ( .D(rC8[3]), .CK(mCLK), .Q(mY4[3]) );
  DFF_X1 \rC8_reg[2]  ( .D(N473), .CK(mCLK), .Q(rC8[2]) );
  DFF_X1 \mY4_reg[2]  ( .D(rC8[2]), .CK(mCLK), .Q(mY4[2]) );
  DFF_X1 \rC8_reg[1]  ( .D(N472), .CK(mCLK), .Q(rC8[1]) );
  DFF_X1 \mY4_reg[1]  ( .D(rC8[1]), .CK(mCLK), .Q(mY4[1]) );
  DFF_X1 \rC8_reg[0]  ( .D(N471), .CK(mCLK), .Q(rC8[0]) );
  DFF_X1 \mY4_reg[0]  ( .D(rC8[0]), .CK(mCLK), .Q(mY4[0]) );
  NAND3_X1 U3023 ( .A1(n2593), .A2(n2448), .A3(n2594), .ZN(n2592) );
  NAND3_X1 U3024 ( .A1(n2603), .A2(n2602), .A3(n2601), .ZN(n2596) );
  NAND3_X1 U3025 ( .A1(n2609), .A2(n3120), .A3(rC7[8]), .ZN(n2608) );
  NAND3_X1 U3026 ( .A1(n3495), .A2(n3182), .A3(rC7[14]), .ZN(n2602) );
  OAI33_X1 U3027 ( .A1(n3016), .A2(rC7[22]), .A3(n2452), .B1(n3061), .B2(
        rC7[23]), .B3(n2630), .ZN(n2629) );
  OAI33_X1 U3028 ( .A1(n3015), .A2(rC7[34]), .A3(n2436), .B1(n3060), .B2(
        rC7[35]), .B3(n2635), .ZN(n2634) );
  OAI33_X1 U3029 ( .A1(n3020), .A2(rC2[49]), .A3(n2214), .B1(n3067), .B2(
        rC2[50]), .B3(n2658), .ZN(n2657) );
  OAI33_X1 U3030 ( .A1(n3184), .A2(rC2[25]), .A3(n2244), .B1(n3066), .B2(
        rC2[26]), .B3(n2679), .ZN(n2678) );
  OAI33_X1 U3031 ( .A1(n3115), .A2(rC4[22]), .A3(n2248), .B1(n3023), .B2(
        rC4[23]), .B3(n2686), .ZN(n2685) );
  OAI33_X1 U3032 ( .A1(n3112), .A2(rC4[16]), .A3(n2690), .B1(n2691), .B2(n2690), .B3(n2692), .ZN(n2689) );
  NAND3_X1 U3033 ( .A1(n3446), .A2(n2698), .A3(n2699), .ZN(n2697) );
  NAND3_X1 U3034 ( .A1(n2700), .A2(n3241), .A3(rC2[10]), .ZN(n2699) );
  OAI33_X1 U3035 ( .A1(n3114), .A2(rC4[46]), .A3(n2218), .B1(n3022), .B2(
        rC4[47]), .B3(n2729), .ZN(n2728) );
  NAND3_X1 U3036 ( .A1(n2732), .A2(n3207), .A3(rC4[61]), .ZN(n2731) );
  NAND3_X1 U3037 ( .A1(n2775), .A2(n2167), .A3(n2776), .ZN(n2774) );
  NAND3_X1 U3038 ( .A1(n2799), .A2(n3091), .A3(rC1[11]), .ZN(n2805) );
  OAI33_X1 U3039 ( .A1(n3019), .A2(rC1[49]), .A3(n2136), .B1(n3065), .B2(
        rC1[50]), .B3(n2817), .ZN(n2751) );
  OAI33_X1 U3040 ( .A1(n3113), .A2(rC3[46]), .A3(n2141), .B1(n3021), .B2(
        rC3[47]), .B3(n2824), .ZN(n2823) );
  NAND3_X1 U3041 ( .A1(n2827), .A2(n3206), .A3(rC3[61]), .ZN(n2826) );
  DFF_X1 \rC7_reg[12]  ( .D(N419), .CK(mCLK), .Q(rC7[12]), .QN(n3684) );
  DFF_X1 \mY2_reg[55]  ( .D(N592), .CK(mCLK), .Q(mY2[55]) );
  DFF_X1 \mY2_reg[56]  ( .D(N593), .CK(mCLK), .Q(mY2[56]) );
  DFF_X1 \mY2_reg[12]  ( .D(N549), .CK(mCLK), .Q(mY2[12]) );
  DFF_X1 \mY3_reg[11]  ( .D(N612), .CK(mCLK), .Q(mY3[11]) );
  DFF_X1 \mY3_reg[1]  ( .D(N602), .CK(mCLK), .Q(mY3[1]) );
  DFF_X1 \mY3_reg[10]  ( .D(N611), .CK(mCLK), .Q(mY3[10]) );
  DFF_X1 \mY3_reg[0]  ( .D(N601), .CK(mCLK), .Q(mY3[0]) );
  DFF_X1 \mY3_reg[2]  ( .D(N603), .CK(mCLK), .Q(mY3[2]) );
  DFF_X1 \mY3_reg[12]  ( .D(N613), .CK(mCLK), .Q(mY3[12]) );
  DFF_X1 \mY2_reg[27]  ( .D(N564), .CK(mCLK), .Q(mY2[27]) );
  DFF_X1 \mY2_reg[30]  ( .D(N567), .CK(mCLK), .Q(mY2[30]) );
  DFF_X1 \mY2_reg[24]  ( .D(N561), .CK(mCLK), .Q(mY2[24]) );
  DFF_X1 \mY2_reg[25]  ( .D(N562), .CK(mCLK), .Q(mY2[25]) );
  DFF_X1 \mY2_reg[26]  ( .D(N563), .CK(mCLK), .Q(mY2[26]) );
  DFF_X1 \mY2_reg[28]  ( .D(N565), .CK(mCLK), .Q(mY2[28]) );
  DFF_X1 \mY2_reg[45]  ( .D(N582), .CK(mCLK), .Q(mY2[45]) );
  DFF_X1 \mY2_reg[46]  ( .D(N583), .CK(mCLK), .Q(mY2[46]) );
  DFF_X1 \mY2_reg[47]  ( .D(N584), .CK(mCLK), .Q(mY2[47]) );
  DFF_X1 \mY2_reg[13]  ( .D(N550), .CK(mCLK), .Q(mY2[13]) );
  DFF_X1 \mY2_reg[14]  ( .D(N551), .CK(mCLK), .Q(mY2[14]) );
  DFF_X1 \mY2_reg[15]  ( .D(N552), .CK(mCLK), .Q(mY2[15]) );
  DFF_X1 \mY2_reg[16]  ( .D(N553), .CK(mCLK), .Q(mY2[16]) );
  DFF_X1 \mY2_reg[17]  ( .D(N554), .CK(mCLK), .Q(mY2[17]) );
  DFF_X1 \mY2_reg[18]  ( .D(N555), .CK(mCLK), .Q(mY2[18]) );
  DFF_X1 \mY2_reg[19]  ( .D(N556), .CK(mCLK), .Q(mY2[19]) );
  DFF_X1 \mY2_reg[20]  ( .D(N557), .CK(mCLK), .Q(mY2[20]) );
  DFF_X1 \mY2_reg[34]  ( .D(N571), .CK(mCLK), .Q(mY2[34]) );
  DFF_X1 \mY2_reg[35]  ( .D(N572), .CK(mCLK), .Q(mY2[35]) );
  DFF_X1 \mY2_reg[49]  ( .D(N586), .CK(mCLK), .Q(mY2[49]) );
  DFF_X1 \mY2_reg[50]  ( .D(N587), .CK(mCLK), .Q(mY2[50]) );
  DFF_X1 \mY2_reg[51]  ( .D(N588), .CK(mCLK), .Q(mY2[51]) );
  DFF_X1 \mY2_reg[52]  ( .D(N589), .CK(mCLK), .Q(mY2[52]) );
  DFF_X1 \mY2_reg[53]  ( .D(N590), .CK(mCLK), .Q(mY2[53]) );
  DFF_X1 \mY2_reg[54]  ( .D(N591), .CK(mCLK), .Q(mY2[54]) );
  DFF_X1 \mY3_reg[45]  ( .D(N646), .CK(mCLK), .Q(mY3[45]) );
  DFF_X1 \mY3_reg[47]  ( .D(N648), .CK(mCLK), .Q(mY3[47]) );
  DFF_X1 \mY3_reg[48]  ( .D(N649), .CK(mCLK), .Q(mY3[48]) );
  DFF_X1 \mY2_reg[29]  ( .D(N566), .CK(mCLK), .Q(mY2[29]) );
  DFF_X1 \mY2_reg[31]  ( .D(N568), .CK(mCLK), .Q(mY2[31]) );
  DFF_X1 \mY2_reg[32]  ( .D(N569), .CK(mCLK), .Q(mY2[32]) );
  DFF_X1 \mY2_reg[60]  ( .D(N597), .CK(mCLK), .Q(mY2[60]) );
  DFF_X1 \mY2_reg[61]  ( .D(N598), .CK(mCLK), .Q(mY2[61]) );
  DFF_X1 \mY2_reg[62]  ( .D(N599), .CK(mCLK), .Q(mY2[62]) );
  DFF_X1 \mY3_reg[4]  ( .D(N605), .CK(mCLK), .Q(mY3[4]) );
  DFF_X1 \mY3_reg[9]  ( .D(N610), .CK(mCLK), .Q(mY3[9]) );
  DFF_X1 \mY3_reg[13]  ( .D(N614), .CK(mCLK), .Q(mY3[13]) );
  DFF_X1 \mY3_reg[16]  ( .D(N617), .CK(mCLK), .Q(mY3[16]) );
  DFF_X1 \mY3_reg[17]  ( .D(N618), .CK(mCLK), .Q(mY3[17]) );
  DFF_X1 \mY3_reg[18]  ( .D(N619), .CK(mCLK), .Q(mY3[18]) );
  DFF_X1 \mY3_reg[19]  ( .D(N620), .CK(mCLK), .Q(mY3[19]) );
  DFF_X1 \mY3_reg[29]  ( .D(N630), .CK(mCLK), .Q(mY3[29]) );
  DFF_X1 \mY3_reg[30]  ( .D(N631), .CK(mCLK), .Q(mY3[30]) );
  DFF_X1 \mY3_reg[20]  ( .D(N621), .CK(mCLK), .Q(mY3[20]) );
  DFF_X1 \mY3_reg[23]  ( .D(N624), .CK(mCLK), .Q(mY3[23]) );
  DFF_X1 \mY3_reg[32]  ( .D(N633), .CK(mCLK), .Q(mY3[32]) );
  DFF_X1 \mY3_reg[33]  ( .D(N634), .CK(mCLK), .Q(mY3[33]) );
  DFF_X1 \mY3_reg[34]  ( .D(N635), .CK(mCLK), .Q(mY3[34]) );
  DFF_X1 \mY3_reg[35]  ( .D(N636), .CK(mCLK), .Q(mY3[35]) );
  DFF_X1 \mY3_reg[36]  ( .D(N637), .CK(mCLK), .Q(mY3[36]) );
  DFF_X1 \mY3_reg[37]  ( .D(N638), .CK(mCLK), .Q(mY3[37]) );
  DFF_X1 \mY3_reg[38]  ( .D(N639), .CK(mCLK), .Q(mY3[38]) );
  DFF_X1 \mY3_reg[39]  ( .D(N640), .CK(mCLK), .Q(mY3[39]) );
  DFF_X1 \mY3_reg[54]  ( .D(N655), .CK(mCLK), .Q(mY3[54]) );
  DFF_X1 \mY3_reg[55]  ( .D(N656), .CK(mCLK), .Q(mY3[55]) );
  DFF_X1 \mY2_reg[36]  ( .D(N573), .CK(mCLK), .Q(mY2[36]) );
  DFF_X1 \mY2_reg[39]  ( .D(N576), .CK(mCLK), .Q(mY2[39]) );
  DFF_X1 \mY2_reg[42]  ( .D(N579), .CK(mCLK), .Q(mY2[42]) );
  DFF_X1 \mY3_reg[44]  ( .D(N645), .CK(mCLK), .Q(mY3[44]) );
  DFF_X1 \mY3_reg[49]  ( .D(N650), .CK(mCLK), .Q(mY3[49]) );
  DFF_X1 \mY3_reg[50]  ( .D(N651), .CK(mCLK), .Q(mY3[50]) );
  DFF_X1 \mY3_reg[51]  ( .D(N652), .CK(mCLK), .Q(mY3[51]) );
  DFF_X1 \mY3_reg[52]  ( .D(N653), .CK(mCLK), .Q(mY3[52]) );
  DFF_X1 \mY3_reg[60]  ( .D(N661), .CK(mCLK), .Q(mY3[60]) );
  DFF_X1 \mY3_reg[61]  ( .D(N662), .CK(mCLK), .Q(mY3[61]) );
  DFF_X1 \mY3_reg[62]  ( .D(N663), .CK(mCLK), .Q(mY3[62]) );
  DFF_X1 \rC8_reg[56]  ( .D(N527), .CK(mCLK), .Q(rC8[56]) );
  DFF_X1 \rC8_reg[33]  ( .D(N504), .CK(mCLK), .Q(rC8[33]) );
  DFF_X1 \rC8_reg[58]  ( .D(N529), .CK(mCLK), .Q(rC8[58]) );
  DFF_X1 \rC8_reg[35]  ( .D(N506), .CK(mCLK), .Q(rC8[35]) );
  DFF_X1 \rC8_reg[37]  ( .D(N508), .CK(mCLK), .Q(rC8[37]) );
  DFF_X1 \rC8_reg[38]  ( .D(N509), .CK(mCLK), .Q(rC8[38]) );
  DFF_X2 \rC5_reg[10]  ( .D(N289), .CK(mCLK), .Q(rC5[10]) );
  DFF_X2 \rC7_reg[15]  ( .D(N422), .CK(mCLK), .Q(rC7[15]), .QN(n3008) );
  DFF_X2 \rC7_reg[18]  ( .D(N425), .CK(mCLK), .Q(rC7[18]), .QN(n3193) );
  DFF_X2 \rC7_reg[56]  ( .D(N463), .CK(mCLK), .Q(rC7[56]), .QN(n3215) );
  DFF_X2 \rC5_reg[44]  ( .D(N323), .CK(mCLK), .Q(rC5[44]) );
  DFF_X2 \rC5_reg[46]  ( .D(N325), .CK(mCLK), .Q(rC5[46]) );
  DFF_X2 \rC7_reg[58]  ( .D(N465), .CK(mCLK), .Q(rC7[58]), .QN(n3237) );
  DFF_X1 \rC7_reg[57]  ( .D(N464), .CK(mCLK), .Q(rC7[57]), .QN(n3275) );
  DFF_X2 \rC5_reg[20]  ( .D(N299), .CK(mCLK), .Q(rC5[20]) );
  DFF_X2 \rC5_reg[19]  ( .D(N298), .CK(mCLK), .Q(rC5[19]) );
  DFF_X2 \rC5_reg[34]  ( .D(N313), .CK(mCLK), .Q(rC5[34]) );
  DFF_X2 \mY3_reg[53]  ( .D(N654), .CK(mCLK), .Q(mY3[53]) );
  DFF_X2 \rC5_reg[51]  ( .D(N330), .CK(mCLK), .Q(rC5[51]) );
  DFF_X2 \rC5_reg[52]  ( .D(N331), .CK(mCLK), .Q(rC5[52]) );
  DFF_X2 \mY3_reg[41]  ( .D(N642), .CK(mCLK), .Q(mY3[41]) );
  DFF_X2 \mY2_reg[40]  ( .D(N577), .CK(mCLK), .Q(mY2[40]) );
  DFF_X1 \rC7_reg[3]  ( .D(N410), .CK(mCLK), .QN(n3685) );
  DFF_X2 \rC5_reg[63]  ( .D(N342), .CK(mCLK), .Q(rC5[63]) );
  DFF_X2 \rC7_reg[21]  ( .D(N428), .CK(mCLK), .Q(rC7[21]), .QN(n3194) );
  DFF_X1 \mY3_reg[3]  ( .D(N604), .CK(mCLK), .Q(mY3[3]) );
  DFF_X1 \mY3_reg[42]  ( .D(N643), .CK(mCLK), .Q(mY3[42]) );
  DFF_X1 \mY3_reg[31]  ( .D(N632), .CK(mCLK), .Q(mY3[31]) );
  DFF_X2 \mY3_reg[27]  ( .D(N628), .CK(mCLK), .Q(mY3[27]) );
  DFF_X2 \mY3_reg[59]  ( .D(N660), .CK(mCLK), .Q(mY3[59]) );
  DFF_X2 \mY3_reg[57]  ( .D(N658), .CK(mCLK), .Q(mY3[57]) );
  DFF_X1 \mY3_reg[40]  ( .D(N641), .CK(mCLK), .Q(mY3[40]) );
  DFF_X1 \mY2_reg[57]  ( .D(N594), .CK(mCLK), .Q(mY2[57]) );
  DFF_X1 \mY2_reg[59]  ( .D(N596), .CK(mCLK), .Q(mY2[59]) );
  DFF_X1 \mY2_reg[63]  ( .D(N600), .CK(mCLK), .Q(mY2[63]) );
  DFF_X1 \mY3_reg[56]  ( .D(N657), .CK(mCLK), .Q(mY3[56]) );
  DFF_X1 \mY3_reg[58]  ( .D(N659), .CK(mCLK), .Q(mY3[58]) );
  DFF_X1 \mY2_reg[37]  ( .D(N574), .CK(mCLK), .Q(mY2[37]) );
  DFF_X2 \mY3_reg[46]  ( .D(N647), .CK(mCLK), .Q(mY3[46]) );
  DFF_X1 \mY2_reg[43]  ( .D(N580), .CK(mCLK), .Q(mY2[43]) );
  DFF_X1 \mY3_reg[14]  ( .D(N615), .CK(mCLK), .Q(mY3[14]) );
  DFF_X1 \mY3_reg[28]  ( .D(N629), .CK(mCLK), .Q(mY3[28]) );
  DFF_X1 \mY3_reg[43]  ( .D(N644), .CK(mCLK), .Q(mY3[43]) );
  DFF_X1 \mY3_reg[21]  ( .D(N622), .CK(mCLK), .Q(mY3[21]) );
  DFF_X1 \mY3_reg[22]  ( .D(N623), .CK(mCLK), .Q(mY3[22]) );
  DFF_X1 \mY3_reg[24]  ( .D(N625), .CK(mCLK), .Q(mY3[24]) );
  DFF_X1 \mY3_reg[25]  ( .D(N626), .CK(mCLK), .Q(mY3[25]) );
  DFF_X1 \mY3_reg[26]  ( .D(N627), .CK(mCLK), .Q(mY3[26]) );
  DFF_X1 \mY3_reg[15]  ( .D(N616), .CK(mCLK), .Q(mY3[15]) );
  DFF_X1 \mY2_reg[38]  ( .D(N575), .CK(mCLK), .Q(mY2[38]) );
  DFF_X1 \mY2_reg[41]  ( .D(N578), .CK(mCLK), .Q(mY2[41]) );
  DFF_X1 \mY2_reg[33]  ( .D(N570), .CK(mCLK), .Q(mY2[33]) );
  DFF_X1 \mY2_reg[44]  ( .D(N581), .CK(mCLK), .Q(mY2[44]) );
  DFF_X1 \mY3_reg[8]  ( .D(N609), .CK(mCLK), .Q(mY3[8]) );
  DFF_X1 \rC7_reg[53]  ( .D(N460), .CK(mCLK), .Q(rC7[53]), .QN(n3026) );
  DFF_X1 \rC7_reg[8]  ( .D(N415), .CK(mCLK), .Q(rC7[8]), .QN(n3204) );
  DFF_X1 \rC5_reg[12]  ( .D(N291), .CK(mCLK), .Q(rC5[12]) );
  DFF_X1 \rC7_reg[7]  ( .D(N414), .CK(mCLK), .Q(rC7[7]), .QN(n3286) );
  DFF_X1 \rC5_reg[54]  ( .D(N333), .CK(mCLK), .Q(rC5[54]) );
  DFF_X1 \rC5_reg[9]  ( .D(N288), .CK(mCLK), .Q(rC5[9]) );
  DFF_X1 \rC5_reg[0]  ( .D(N279), .CK(mCLK), .Q(rC5[0]) );
  DFF_X1 \rC7_reg[52]  ( .D(N459), .CK(mCLK), .Q(rC7[52]), .QN(n3098) );
  DFF_X1 \rC5_reg[42]  ( .D(N321), .CK(mCLK), .Q(rC5[42]) );
  DFF_X1 \rC5_reg[59]  ( .D(N338), .CK(mCLK), .Q(rC5[59]) );
  DFF_X1 \rC7_reg[14]  ( .D(N421), .CK(mCLK), .Q(rC7[14]), .QN(n3087) );
  DFF_X1 \rC5_reg[57]  ( .D(N336), .CK(mCLK), .Q(rC5[57]) );
  DFF_X1 \rC7_reg[38]  ( .D(N445), .CK(mCLK), .Q(rC7[38]), .QN(n3037) );
  DFF_X1 \rC7_reg[24]  ( .D(N431), .CK(mCLK), .Q(rC7[24]), .QN(n3054) );
  DFF_X1 \rC7_reg[5]  ( .D(N412), .CK(mCLK), .Q(rC7[5]), .QN(n3259) );
  DFF_X1 \rC7_reg[22]  ( .D(N429), .CK(mCLK), .Q(rC7[22]), .QN(n3279) );
  DFF_X1 \rC7_reg[17]  ( .D(N424), .CK(mCLK), .Q(rC7[17]), .QN(n3268) );
  DFF_X1 \rC5_reg[47]  ( .D(N326), .CK(mCLK), .Q(rC5[47]) );
  DFF_X1 \rC7_reg[0]  ( .D(N407), .CK(mCLK), .Q(rC7[0]), .QN(n3347) );
  DFF_X1 \rC7_reg[36]  ( .D(N443), .CK(mCLK), .Q(rC7[36]), .QN(n3055) );
  DFF_X1 \rC5_reg[45]  ( .D(N324), .CK(mCLK), .Q(rC5[45]) );
  DFF_X1 \rC7_reg[43]  ( .D(N450), .CK(mCLK), .Q(rC7[43]), .QN(n3097) );
  DFF_X1 \rC5_reg[8]  ( .D(N287), .CK(mCLK), .Q(rC5[8]) );
  DFF_X1 \rC5_reg[56]  ( .D(N335), .CK(mCLK), .Q(rC5[56]) );
  DFF_X1 \rC5_reg[62]  ( .D(N341), .CK(mCLK), .Q(rC5[62]) );
  DFF_X1 \rC5_reg[61]  ( .D(N340), .CK(mCLK), .Q(rC5[61]) );
  DFF_X1 \rC7_reg[23]  ( .D(N430), .CK(mCLK), .Q(rC7[23]), .QN(n3272) );
  DFF_X1 \rC7_reg[25]  ( .D(N432), .CK(mCLK), .Q(rC7[25]), .QN(n3274) );
  DFF_X1 \rC7_reg[1]  ( .D(N408), .CK(mCLK), .Q(rC7[1]), .QN(n3345) );
  DFF_X1 \rC7_reg[61]  ( .D(N468), .CK(mCLK), .Q(rC7[61]), .QN(n3343) );
  DFF_X1 \rC7_reg[4]  ( .D(N411), .CK(mCLK), .Q(rC7[4]), .QN(n3254) );
  DFF_X1 \rC7_reg[16]  ( .D(N423), .CK(mCLK), .Q(rC7[16]), .QN(n3217) );
  DFF_X1 \rC7_reg[6]  ( .D(N413), .CK(mCLK), .Q(rC7[6]), .QN(n3191) );
  DFF_X1 \rC7_reg[59]  ( .D(N466), .CK(mCLK), .Q(rC7[59]), .QN(n3147) );
  DFF_X1 \rC7_reg[55]  ( .D(N462), .CK(mCLK), .Q(rC7[55]), .QN(n3133) );
  DFF_X1 \rC7_reg[28]  ( .D(N435), .CK(mCLK), .Q(rC7[28]), .QN(n3018) );
  DFF_X1 \rC5_reg[14]  ( .D(N293), .CK(mCLK), .Q(rC5[14]) );
  DFF_X1 \rC5_reg[15]  ( .D(N294), .CK(mCLK), .Q(rC5[15]) );
  DFF_X1 \rC5_reg[31]  ( .D(N310), .CK(mCLK), .Q(rC5[31]) );
  DFF_X1 \rC5_reg[43]  ( .D(N322), .CK(mCLK), .Q(rC5[43]) );
  DFF_X1 \rC7_reg[54]  ( .D(N461), .CK(mCLK), .Q(rC7[54]), .QN(n3216) );
  DFF_X1 \rC5_reg[7]  ( .D(N286), .CK(mCLK), .Q(rC5[7]) );
  DFF_X1 \rC5_reg[49]  ( .D(N328), .CK(mCLK), .Q(rC5[49]) );
  DFF_X2 \mY2_reg[58]  ( .D(N595), .CK(mCLK), .Q(mY2[58]) );
  DFF_X1 \rC5_reg[6]  ( .D(N285), .CK(mCLK), .Q(rC5[6]) );
  DFF_X1 \rC7_reg[26]  ( .D(N433), .CK(mCLK), .Q(rC7[26]), .QN(n3344) );
  DFF_X1 \rC5_reg[48]  ( .D(N327), .CK(mCLK), .Q(rC5[48]) );
  DFF_X1 \rC5_reg[58]  ( .D(N337), .CK(mCLK), .Q(rC5[58]) );
  DFF_X1 \rC7_reg[20]  ( .D(N427), .CK(mCLK), .QN(n3092) );
  DFF_X1 \rC5_reg[18]  ( .D(N297), .CK(mCLK), .Q(rC5[18]) );
  DFF_X1 \rC7_reg[37]  ( .D(N444), .CK(mCLK), .Q(rC7[37]), .QN(n3134) );
  DFF_X1 \rC7_reg[60]  ( .D(N467), .CK(mCLK), .Q(rC7[60]), .QN(n3218) );
  DFF_X1 \rC5_reg[3]  ( .D(N282), .CK(mCLK), .Q(rC5[3]) );
  DFF_X1 \rC5_reg[13]  ( .D(N292), .CK(mCLK), .Q(rC5[13]) );
  DFF_X1 \rC5_reg[53]  ( .D(N332), .CK(mCLK), .Q(rC5[53]) );
  DFF_X1 \rC7_reg[19]  ( .D(N426), .CK(mCLK), .Q(rC7[19]), .QN(n3255) );
  DFF_X1 \rC5_reg[60]  ( .D(N339), .CK(mCLK), .Q(rC5[60]) );
  DFF_X1 \rC7_reg[27]  ( .D(N434), .CK(mCLK), .Q(rC7[27]), .QN(n3249) );
  DFF_X1 \rC5_reg[55]  ( .D(N334), .CK(mCLK), .Q(rC5[55]) );
  DFF_X1 \rC5_reg[5]  ( .D(N284), .CK(mCLK), .Q(rC5[5]) );
  INV_X1 U3042 ( .A(n3624), .ZN(n2970) );
  BUF_X2 U3043 ( .A(n3456), .Z(n2979) );
  BUF_X1 U3044 ( .A(n3615), .Z(n2972) );
  BUF_X1 U3045 ( .A(n3448), .Z(n2978) );
  BUF_X1 U3046 ( .A(n3456), .Z(n3627) );
  BUF_X1 U3047 ( .A(n3748), .Z(n3667) );
  CLKBUF_X1 U3048 ( .A(n3625), .Z(n3630) );
  INV_X1 U3049 ( .A(n3741), .ZN(n2983) );
  INV_X1 U3050 ( .A(n3620), .ZN(n2984) );
  BUF_X1 U3051 ( .A(n3389), .Z(n2985) );
  BUF_X1 U3052 ( .A(n3389), .Z(n2986) );
  INV_X1 U3053 ( .A(n3743), .ZN(n2987) );
  BUF_X1 U3054 ( .A(n3620), .Z(n3743) );
  INV_X1 U3055 ( .A(n3791), .ZN(n3753) );
  INV_X1 U3056 ( .A(n3791), .ZN(n2989) );
  INV_X1 U3057 ( .A(n3791), .ZN(n2990) );
  INV_X1 U3058 ( .A(n3791), .ZN(n3755) );
  BUF_X1 U3059 ( .A(n3501), .Z(n2991) );
  BUF_X1 U3060 ( .A(n3501), .Z(n2992) );
  BUF_X1 U3061 ( .A(n3501), .Z(n2993) );
  BUF_X1 U3062 ( .A(n3788), .Z(n2994) );
  INV_X1 U3063 ( .A(n3778), .ZN(n2995) );
  BUF_X2 U3064 ( .A(n3787), .Z(n3778) );
  CLKBUF_X1 U3065 ( .A(n3751), .Z(n3501) );
  INV_X1 U3066 ( .A(n3786), .ZN(n3758) );
  NAND2_X1 U3067 ( .A1(n3525), .A2(n3524), .ZN(n2997) );
  NAND2_X1 U3068 ( .A1(n2592), .A2(n2998), .ZN(n2585) );
  INV_X1 U3069 ( .A(n2997), .ZN(n2998) );
  CLKBUF_X1 U3070 ( .A(n3681), .Z(n2999) );
  INV_X1 U3071 ( .A(n3681), .ZN(n3000) );
  BUF_X1 U3072 ( .A(n3611), .Z(n3470) );
  OR3_X1 U3073 ( .A1(n3682), .A2(n3688), .A3(n2620), .ZN(n3350) );
  AND2_X1 U3074 ( .A1(n3425), .A2(n3426), .ZN(n3351) );
  AND2_X1 U3075 ( .A1(n3516), .A2(n3517), .ZN(n3352) );
  AND2_X1 U3076 ( .A1(n3506), .A2(n3505), .ZN(n3353) );
  OR2_X1 U3077 ( .A1(n3690), .A2(n3689), .ZN(n3354) );
  OR2_X1 U3078 ( .A1(n3523), .A2(n3522), .ZN(n3355) );
  OR2_X1 U3079 ( .A1(n3521), .A2(n3520), .ZN(n3356) );
  BUF_X1 U3080 ( .A(n3475), .Z(n3664) );
  BUF_X2 U3081 ( .A(n3749), .Z(n3741) );
  BUF_X2 U3082 ( .A(n3491), .Z(n3641) );
  CLKBUF_X1 U3083 ( .A(n3625), .Z(n3626) );
  BUF_X2 U3084 ( .A(n3611), .Z(n3469) );
  BUF_X1 U3085 ( .A(n3741), .Z(n3639) );
  BUF_X1 U3086 ( .A(n3741), .Z(n3647) );
  BUF_X1 U3087 ( .A(n3750), .Z(n3476) );
  BUF_X2 U3088 ( .A(n3613), .Z(n3740) );
  BUF_X2 U3089 ( .A(n3746), .Z(n3742) );
  BUF_X1 U3090 ( .A(n3476), .Z(n3739) );
  BUF_X1 U3091 ( .A(n3623), .Z(n3738) );
  BUF_X1 U3092 ( .A(n3624), .Z(n3628) );
  BUF_X1 U3093 ( .A(n3624), .Z(n3629) );
  BUF_X1 U3094 ( .A(n3624), .Z(n3642) );
  BUF_X1 U3095 ( .A(n3620), .Z(n3736) );
  BUF_X1 U3096 ( .A(n3747), .Z(n3737) );
  CLKBUF_X3 U3097 ( .A(n3749), .Z(n3625) );
  BUF_X1 U3098 ( .A(n3456), .Z(n3643) );
  INV_X1 U3099 ( .A(n3382), .ZN(n3371) );
  INV_X1 U3100 ( .A(n3792), .ZN(n3372) );
  INV_X1 U3101 ( .A(n3792), .ZN(n3373) );
  INV_X1 U3102 ( .A(n3792), .ZN(n3754) );
  BUF_X2 U3103 ( .A(n3735), .Z(n3671) );
  INV_X1 U3104 ( .A(n3387), .ZN(n3375) );
  INV_X1 U3105 ( .A(n3376), .ZN(n3377) );
  INV_X1 U3106 ( .A(n3378), .ZN(n3379) );
  INV_X1 U3107 ( .A(n3786), .ZN(n3380) );
  BUF_X2 U3108 ( .A(n3787), .Z(n3772) );
  BUF_X2 U3109 ( .A(n3785), .Z(n3784) );
  INV_X1 U3110 ( .A(n3792), .ZN(n3752) );
  INV_X1 U3111 ( .A(n3382), .ZN(n3383) );
  BUF_X1 U3112 ( .A(n3793), .Z(n3785) );
  BUF_X1 U3113 ( .A(n3793), .Z(n3787) );
  INV_X1 U3114 ( .A(n3384), .ZN(n3385) );
  INV_X1 U3115 ( .A(n3786), .ZN(n3386) );
  INV_X1 U3116 ( .A(n3387), .ZN(n3388) );
  INV_X1 U3117 ( .A(n3751), .ZN(n3389) );
  BUF_X2 U3118 ( .A(n2639), .Z(n3751) );
  INV_X1 U3119 ( .A(n3786), .ZN(n3390) );
  INV_X1 U3120 ( .A(n3786), .ZN(n3391) );
  CLKBUF_X1 U3121 ( .A(n2696), .Z(n3392) );
  INV_X1 U3122 ( .A(n3822), .ZN(n3800) );
  INV_X2 U3123 ( .A(n3834), .ZN(n3804) );
  AOI221_X1 U3124 ( .B1(n3089), .B2(rC6[33]), .C1(n3009), .C2(rC6[32]), .A(
        n2577), .ZN(n3395) );
  OAI211_X1 U3125 ( .C1(rC2[12]), .C2(n3498), .A(n3396), .B(n3397), .ZN(n2705)
         );
  OAI21_X1 U3126 ( .B1(n2687), .B2(n3356), .A(n3398), .ZN(n3399) );
  INV_X1 U3127 ( .A(n2682), .ZN(n3398) );
  INV_X1 U3128 ( .A(n3399), .ZN(n2675) );
  AOI22_X1 U3129 ( .A1(n3400), .A2(rC1[3]), .B1(n3401), .B2(rC1[2]), .ZN(n2802) );
  AOI211_X1 U3130 ( .C1(n2746), .C2(n2745), .A(n2122), .B(n2747), .ZN(n2744)
         );
  AOI211_X1 U3131 ( .C1(n3402), .C2(rC7[12]), .A(rC7[11]), .B(n3678), .ZN(
        n2619) );
  OAI211_X1 U3132 ( .C1(n2474), .C2(n2622), .A(n3507), .B(n2623), .ZN(n2615)
         );
  OAI221_X1 U3133 ( .B1(n2271), .B2(n2713), .C1(rC2[3]), .C2(n3450), .A(n2714), 
        .ZN(n2708) );
  OAI22_X1 U3134 ( .A1(n3403), .A2(rC6[13]), .B1(n2610), .B2(n2611), .ZN(n2605) );
  BUF_X1 U3135 ( .A(n3833), .Z(n3828) );
  INV_X2 U3136 ( .A(n3785), .ZN(n3759) );
  INV_X2 U3137 ( .A(n3785), .ZN(n3760) );
  OAI211_X1 U3138 ( .C1(rC3[12]), .C2(n2183), .A(n2179), .B(n2805), .ZN(n3418)
         );
  AOI22_X1 U3139 ( .A1(n3416), .A2(rC1[15]), .B1(n3371), .B2(n3447), .ZN(n3421) );
  NAND2_X1 U3140 ( .A1(n2570), .A2(n3351), .ZN(n2563) );
  BUF_X1 U3141 ( .A(n3389), .Z(n3422) );
  NOR2_X1 U3142 ( .A1(n2648), .A2(n3354), .ZN(n2643) );
  BUF_X1 U3143 ( .A(n3827), .Z(n3617) );
  OR2_X1 U3144 ( .A1(n2568), .A2(n2569), .ZN(n3425) );
  OR2_X1 U3145 ( .A1(rC6[45]), .A2(n3251), .ZN(n3426) );
  BUF_X1 U3146 ( .A(n3790), .Z(n3427) );
  BUF_X1 U3147 ( .A(n3788), .Z(n3428) );
  BUF_X1 U3148 ( .A(n3389), .Z(n3429) );
  OAI22_X1 U3149 ( .A1(rC6[12]), .A2(n3684), .B1(rC6[11]), .B2(n3686), .ZN(
        n3431) );
  BUF_X1 U3150 ( .A(n3829), .Z(n3814) );
  BUF_X1 U3151 ( .A(n3823), .Z(n3826) );
  OAI22_X1 U3152 ( .A1(rC3[9]), .A2(n3419), .B1(n3385), .B2(n3375), .ZN(n3444)
         );
  INV_X1 U3153 ( .A(n3816), .ZN(n3445) );
  BUF_X1 U3154 ( .A(n3832), .Z(n3810) );
  CLKBUF_X1 U3155 ( .A(n2259), .Z(n3446) );
  INV_X1 U3156 ( .A(n3616), .ZN(n3448) );
  INV_X1 U3157 ( .A(n3816), .ZN(n3449) );
  BUF_X2 U3158 ( .A(n3831), .Z(n3816) );
  BUF_X1 U3159 ( .A(n3475), .Z(n3665) );
  CLKBUF_X1 U3160 ( .A(n3431), .Z(n3452) );
  BUF_X2 U3161 ( .A(n3834), .Z(n3609) );
  BUF_X1 U3162 ( .A(n3491), .Z(n3634) );
  BUF_X2 U3163 ( .A(n3831), .Z(n3808) );
  INV_X1 U3164 ( .A(n3816), .ZN(n3454) );
  CLKBUF_X1 U3165 ( .A(n3625), .Z(n3656) );
  BUF_X1 U3166 ( .A(n3750), .Z(n3456) );
  CLKBUF_X1 U3167 ( .A(n3741), .Z(n3654) );
  BUF_X2 U3168 ( .A(n3735), .Z(n3459) );
  INV_X1 U3169 ( .A(n3816), .ZN(n3460) );
  INV_X1 U3170 ( .A(n3816), .ZN(n3461) );
  BUF_X2 U3171 ( .A(n3832), .Z(n3817) );
  INV_X1 U3172 ( .A(n3462), .ZN(n3463) );
  BUF_X1 U3173 ( .A(n3827), .Z(n3468) );
  CLKBUF_X1 U3174 ( .A(n3486), .Z(n3471) );
  INV_X1 U3175 ( .A(n3748), .ZN(n3472) );
  BUF_X1 U3176 ( .A(n3749), .Z(n3748) );
  INV_X1 U3177 ( .A(n3741), .ZN(n3473) );
  INV_X1 U3178 ( .A(n3612), .ZN(n3475) );
  INV_X1 U3179 ( .A(n3625), .ZN(n3481) );
  INV_X1 U3180 ( .A(n3482), .ZN(n3483) );
  INV_X1 U3181 ( .A(n3486), .ZN(n3487) );
  OR2_X1 U3182 ( .A1(rC4[0]), .A2(n3455), .ZN(n3488) );
  OR2_X1 U3183 ( .A1(rC4[1]), .A2(n3480), .ZN(n3489) );
  NAND3_X1 U3184 ( .A1(n3488), .A2(n2715), .A3(n3489), .ZN(n2714) );
  NAND2_X1 U3185 ( .A1(n2562), .A2(n3352), .ZN(n2558) );
  INV_X1 U3186 ( .A(n3673), .ZN(n3491) );
  CLKBUF_X1 U3187 ( .A(n2640), .Z(n3673) );
  NAND2_X1 U3188 ( .A1(n2595), .A2(n3353), .ZN(n2593) );
  OR2_X1 U3189 ( .A1(rC6[4]), .A2(n3254), .ZN(n3493) );
  NAND2_X1 U3190 ( .A1(n3493), .A2(n2613), .ZN(n2616) );
  BUF_X1 U3191 ( .A(n3829), .Z(n3494) );
  AOI22_X1 U3192 ( .A1(n3008), .A2(rC6[15]), .B1(n3087), .B2(rC6[14]), .ZN(
        n3495) );
  NOR2_X1 U3193 ( .A1(n2627), .A2(n3350), .ZN(n2606) );
  INV_X2 U3194 ( .A(n3822), .ZN(n3795) );
  AOI22_X1 U3195 ( .A1(n3008), .A2(rC6[15]), .B1(n3087), .B2(rC6[14]), .ZN(
        n2604) );
  AOI22_X1 U3196 ( .A1(n3685), .A2(rC6[3]), .B1(rC6[2]), .B2(n3687), .ZN(n3496) );
  INV_X1 U3197 ( .A(n3751), .ZN(n3499) );
  CLKBUF_X1 U3198 ( .A(n3625), .Z(n3637) );
  CLKBUF_X1 U3199 ( .A(n3625), .Z(n3635) );
  INV_X1 U3200 ( .A(n3751), .ZN(n3792) );
  AND2_X1 U3201 ( .A1(n3502), .A2(n3513), .ZN(n2650) );
  NAND2_X1 U3202 ( .A1(n2655), .A2(n2654), .ZN(n3502) );
  NOR2_X1 U3203 ( .A1(n2744), .A2(n3355), .ZN(n2739) );
  OR2_X1 U3204 ( .A1(rC1[19]), .A2(n3256), .ZN(n3503) );
  OR2_X1 U3205 ( .A1(rC1[20]), .A2(n3093), .ZN(n3504) );
  NAND3_X1 U3206 ( .A1(n2777), .A2(n3504), .A3(n3503), .ZN(n2775) );
  OR2_X1 U3207 ( .A1(rC6[19]), .A2(n3255), .ZN(n3505) );
  OR2_X1 U3208 ( .A1(rC6[20]), .A2(n3092), .ZN(n3506) );
  OR2_X1 U3209 ( .A1(rC6[3]), .A2(n3685), .ZN(n3507) );
  AND3_X1 U3210 ( .A1(n3510), .A2(n3509), .A3(n3508), .ZN(n2552) );
  NAND2_X1 U3211 ( .A1(rC7[57]), .A2(n3024), .ZN(n3508) );
  NAND2_X1 U3212 ( .A1(n2413), .A2(n2553), .ZN(n3509) );
  OR3_X1 U3213 ( .A1(n2556), .A2(n2555), .A3(n2557), .ZN(n3510) );
  OR2_X2 U3214 ( .A1(n2771), .A2(n2166), .ZN(n3511) );
  OR2_X1 U3215 ( .A1(n2772), .A2(n2773), .ZN(n3512) );
  NAND3_X1 U3216 ( .A1(n2774), .A2(n3512), .A3(n3511), .ZN(n2768) );
  AOI221_X4 U3217 ( .B1(rC3[21]), .B2(n3130), .C1(rC3[22]), .C2(n3014), .A(
        n2811), .ZN(n2772) );
  NOR2_X1 U3218 ( .A1(n3598), .A2(n2657), .ZN(n3513) );
  OR2_X1 U3219 ( .A1(n2694), .A2(n2693), .ZN(n3514) );
  OR2_X1 U3220 ( .A1(n2695), .A2(n3392), .ZN(n3515) );
  NAND3_X1 U3221 ( .A1(n3514), .A2(n2697), .A3(n3515), .ZN(n2691) );
  OR2_X1 U3222 ( .A1(n2560), .A2(n2561), .ZN(n3516) );
  OR2_X1 U3223 ( .A1(rC6[51]), .A2(n3250), .ZN(n3517) );
  AND2_X1 U3224 ( .A1(rC3[3]), .A2(n3252), .ZN(n3518) );
  AND2_X1 U3225 ( .A1(n2802), .A2(n2803), .ZN(n3519) );
  NOR3_X1 U3226 ( .A1(n3518), .A2(n3519), .A3(n2192), .ZN(n2797) );
  AND2_X1 U3227 ( .A1(rC4[20]), .A2(n3253), .ZN(n3520) );
  AND2_X1 U3228 ( .A1(rC4[19]), .A2(n3094), .ZN(n3521) );
  OR2_X1 U3229 ( .A1(n2588), .A2(n2589), .ZN(n3524) );
  AND2_X1 U3230 ( .A1(n2740), .A2(n2741), .ZN(n3522) );
  AND2_X1 U3231 ( .A1(n2742), .A2(n2743), .ZN(n3523) );
  AOI221_X1 U3232 ( .B1(rC7[21]), .B2(n3117), .C1(rC7[22]), .C2(n3016), .A(
        n2452), .ZN(n2590) );
  OR2_X1 U3233 ( .A1(n2590), .A2(n2591), .ZN(n3525) );
  BUF_X1 U3234 ( .A(n3789), .Z(n3765) );
  BUF_X1 U3235 ( .A(n3389), .Z(n3766) );
  BUF_X1 U3236 ( .A(n3790), .Z(n3762) );
  BUF_X1 U3237 ( .A(n3790), .Z(n3763) );
  BUF_X1 U3238 ( .A(n3389), .Z(n3764) );
  BUF_X1 U3239 ( .A(n3789), .Z(n3768) );
  BUF_X1 U3240 ( .A(n3389), .Z(n3769) );
  BUF_X1 U3241 ( .A(n3789), .Z(n3767) );
  BUF_X1 U3242 ( .A(n3788), .Z(n3776) );
  BUF_X1 U3243 ( .A(n3389), .Z(n3777) );
  BUF_X1 U3244 ( .A(n3389), .Z(n3773) );
  BUF_X1 U3245 ( .A(n3389), .Z(n3774) );
  BUF_X1 U3246 ( .A(n3389), .Z(n3775) );
  BUF_X1 U3247 ( .A(n3792), .Z(n3771) );
  BUF_X1 U3248 ( .A(n3792), .Z(n3770) );
  INV_X1 U3249 ( .A(n3868), .ZN(n3837) );
  INV_X1 U3250 ( .A(n3723), .ZN(n3695) );
  INV_X1 U3251 ( .A(n3723), .ZN(n3694) );
  INV_X1 U3252 ( .A(n3723), .ZN(n3693) );
  INV_X1 U3253 ( .A(n3723), .ZN(n3692) );
  INV_X1 U3254 ( .A(n3868), .ZN(n3840) );
  INV_X1 U3255 ( .A(n3868), .ZN(n3839) );
  INV_X1 U3256 ( .A(n3868), .ZN(n3838) );
  INV_X1 U3257 ( .A(n3724), .ZN(n3697) );
  INV_X1 U3258 ( .A(n3724), .ZN(n3696) );
  INV_X1 U3259 ( .A(n3869), .ZN(n3842) );
  INV_X1 U3260 ( .A(n3869), .ZN(n3841) );
  INV_X1 U3261 ( .A(n3786), .ZN(n3757) );
  INV_X1 U3262 ( .A(n3786), .ZN(n3756) );
  BUF_X1 U3263 ( .A(n3614), .Z(n3813) );
  BUF_X1 U3264 ( .A(n3787), .Z(n3779) );
  BUF_X1 U3265 ( .A(n3787), .Z(n3780) );
  BUF_X1 U3266 ( .A(n3786), .Z(n3783) );
  BUF_X1 U3267 ( .A(n3786), .Z(n3781) );
  BUF_X1 U3268 ( .A(n3786), .Z(n3782) );
  BUF_X1 U3269 ( .A(n3499), .Z(n3789) );
  BUF_X1 U3270 ( .A(n3499), .Z(n3790) );
  BUF_X1 U3271 ( .A(n3499), .Z(n3788) );
  BUF_X1 U3272 ( .A(n3725), .Z(n3723) );
  BUF_X1 U3273 ( .A(n3870), .Z(n3868) );
  BUF_X1 U3274 ( .A(n3725), .Z(n3724) );
  BUF_X1 U3275 ( .A(n3870), .Z(n3869) );
  BUF_X1 U3276 ( .A(n3877), .Z(n3848) );
  BUF_X1 U3277 ( .A(n3878), .Z(n3845) );
  BUF_X1 U3278 ( .A(n3878), .Z(n3843) );
  BUF_X1 U3279 ( .A(n3878), .Z(n3844) );
  BUF_X1 U3280 ( .A(n3870), .Z(n3867) );
  BUF_X1 U3281 ( .A(n3871), .Z(n3864) );
  BUF_X1 U3282 ( .A(n3872), .Z(n3862) );
  BUF_X1 U3283 ( .A(n3726), .Z(n3721) );
  BUF_X1 U3284 ( .A(n3725), .Z(n3722) );
  BUF_X1 U3285 ( .A(n3726), .Z(n3719) );
  BUF_X1 U3286 ( .A(n3726), .Z(n3720) );
  BUF_X1 U3287 ( .A(n3727), .Z(n3717) );
  BUF_X1 U3288 ( .A(n3727), .Z(n3718) );
  BUF_X1 U3289 ( .A(n3728), .Z(n3714) );
  BUF_X1 U3290 ( .A(n3728), .Z(n3715) );
  BUF_X1 U3291 ( .A(n3727), .Z(n3716) );
  BUF_X1 U3292 ( .A(n3729), .Z(n3712) );
  BUF_X1 U3293 ( .A(n3728), .Z(n3713) );
  BUF_X1 U3294 ( .A(n3730), .Z(n3709) );
  BUF_X1 U3295 ( .A(n3729), .Z(n3710) );
  BUF_X1 U3296 ( .A(n3729), .Z(n3711) );
  BUF_X1 U3297 ( .A(n3730), .Z(n3707) );
  BUF_X1 U3298 ( .A(n3730), .Z(n3708) );
  BUF_X1 U3299 ( .A(n3731), .Z(n3705) );
  BUF_X1 U3300 ( .A(n3731), .Z(n3706) );
  BUF_X1 U3301 ( .A(n3732), .Z(n3702) );
  BUF_X1 U3302 ( .A(n3732), .Z(n3703) );
  BUF_X1 U3303 ( .A(n3731), .Z(n3704) );
  BUF_X1 U3304 ( .A(n3733), .Z(n3700) );
  BUF_X1 U3305 ( .A(n3732), .Z(n3701) );
  BUF_X1 U3306 ( .A(n3733), .Z(n3698) );
  BUF_X1 U3307 ( .A(n3733), .Z(n3699) );
  BUF_X1 U3308 ( .A(n3871), .Z(n3866) );
  BUF_X1 U3309 ( .A(n3871), .Z(n3865) );
  BUF_X1 U3310 ( .A(n3872), .Z(n3863) );
  BUF_X1 U3311 ( .A(n3873), .Z(n3859) );
  BUF_X1 U3312 ( .A(n3873), .Z(n3860) );
  BUF_X1 U3313 ( .A(n3872), .Z(n3861) );
  BUF_X1 U3314 ( .A(n3874), .Z(n3857) );
  BUF_X1 U3315 ( .A(n3873), .Z(n3858) );
  BUF_X1 U3316 ( .A(n3875), .Z(n3854) );
  BUF_X1 U3317 ( .A(n3874), .Z(n3855) );
  BUF_X1 U3318 ( .A(n3874), .Z(n3856) );
  BUF_X1 U3319 ( .A(n3875), .Z(n3852) );
  BUF_X1 U3320 ( .A(n3875), .Z(n3853) );
  BUF_X1 U3321 ( .A(n3876), .Z(n3849) );
  BUF_X1 U3322 ( .A(n3876), .Z(n3850) );
  BUF_X1 U3323 ( .A(n3876), .Z(n3851) );
  BUF_X1 U3324 ( .A(n3877), .Z(n3846) );
  BUF_X1 U3325 ( .A(n3877), .Z(n3847) );
  BUF_X2 U3326 ( .A(n3793), .Z(n3786) );
  BUF_X1 U3327 ( .A(n3750), .Z(n3746) );
  BUF_X1 U3328 ( .A(n3750), .Z(n3747) );
  BUF_X1 U3329 ( .A(n3734), .Z(n3725) );
  BUF_X1 U3330 ( .A(n3879), .Z(n3870) );
  BUF_X1 U3331 ( .A(n3873), .Z(n3878) );
  BUF_X1 U3332 ( .A(n3734), .Z(n3726) );
  BUF_X1 U3333 ( .A(n3734), .Z(n3727) );
  BUF_X1 U3334 ( .A(n3734), .Z(n3728) );
  BUF_X1 U3335 ( .A(n3725), .Z(n3729) );
  BUF_X1 U3336 ( .A(n3726), .Z(n3730) );
  BUF_X1 U3337 ( .A(n3728), .Z(n3731) );
  BUF_X1 U3338 ( .A(n3729), .Z(n3732) );
  BUF_X1 U3339 ( .A(n3730), .Z(n3733) );
  BUF_X1 U3340 ( .A(n3879), .Z(n3871) );
  BUF_X1 U3341 ( .A(n3879), .Z(n3872) );
  BUF_X1 U3342 ( .A(n3879), .Z(n3873) );
  BUF_X1 U3343 ( .A(n3870), .Z(n3874) );
  BUF_X1 U3344 ( .A(n3871), .Z(n3875) );
  BUF_X1 U3345 ( .A(n3874), .Z(n3876) );
  BUF_X1 U3346 ( .A(n3875), .Z(n3877) );
  OAI22_X1 U3347 ( .A1(n3648), .A2(n3298), .B1(n3049), .B2(n3670), .ZN(N441)
         );
  OAI22_X1 U3348 ( .A1(n3643), .A2(n3150), .B1(n3210), .B2(n3670), .ZN(N302)
         );
  OAI22_X1 U3349 ( .A1(n3637), .A2(n3149), .B1(n3209), .B2(n3670), .ZN(N314)
         );
  OAI22_X1 U3350 ( .A1(n3742), .A2(n3245), .B1(n3153), .B2(n3622), .ZN(N316)
         );
  OAI22_X1 U3351 ( .A1(n3634), .A2(n3247), .B1(n3151), .B2(n3622), .ZN(N417)
         );
  OAI22_X1 U3352 ( .A1(n3634), .A2(n3091), .B1(n3296), .B2(n3670), .ZN(N418)
         );
  OAI22_X1 U3353 ( .A1(n3633), .A2(n3211), .B1(n3118), .B2(n3670), .ZN(N420)
         );
  OAI22_X1 U3354 ( .A1(n3631), .A2(n3154), .B1(n3238), .B2(n3622), .ZN(N438)
         );
  OAI22_X1 U3355 ( .A1(n3740), .A2(n3043), .B1(n3299), .B2(n3622), .ZN(N439)
         );
  OAI22_X1 U3356 ( .A1(n3636), .A2(n3075), .B1(n3178), .B2(n3622), .ZN(N443)
         );
  OAI22_X1 U3357 ( .A1(n3667), .A2(n3028), .B1(n3330), .B2(n3670), .ZN(N447)
         );
  OAI22_X1 U3358 ( .A1(n3661), .A2(n3221), .B1(n3162), .B2(n3622), .ZN(N451)
         );
  OAI22_X1 U3359 ( .A1(n3666), .A2(n3232), .B1(n3113), .B2(n3670), .ZN(N453)
         );
  OAI22_X1 U3360 ( .A1(n3639), .A2(n3314), .B1(n3021), .B2(n3670), .ZN(N454)
         );
  OAI22_X1 U3361 ( .A1(n3628), .A2(n3102), .B1(n3187), .B2(n3670), .ZN(N455)
         );
  OAI22_X1 U3362 ( .A1(n3631), .A2(n3065), .B1(n3313), .B2(n3622), .ZN(N457)
         );
  OAI22_X1 U3363 ( .A1(n2979), .A2(n3320), .B1(n3056), .B2(n3670), .ZN(N458)
         );
  OAI22_X1 U3364 ( .A1(n3742), .A2(n3130), .B1(n3202), .B2(n3622), .ZN(N300)
         );
  OAI22_X1 U3365 ( .A1(n3654), .A2(n3014), .B1(n3329), .B2(n3622), .ZN(N301)
         );
  OAI22_X1 U3366 ( .A1(n3632), .A2(n3079), .B1(n3321), .B2(n3622), .ZN(N304)
         );
  OAI22_X1 U3367 ( .A1(n3629), .A2(n3235), .B1(n3168), .B2(n3670), .ZN(N305)
         );
  OAI22_X1 U3368 ( .A1(n3628), .A2(n3290), .B1(n3007), .B2(n3622), .ZN(N306)
         );
  OAI22_X1 U3369 ( .A1(n3640), .A2(n3331), .B1(n3029), .B2(n3622), .ZN(N307)
         );
  OAI22_X1 U3370 ( .A1(n2979), .A2(n3229), .B1(n3144), .B2(n3670), .ZN(N308)
         );
  OAI22_X1 U3371 ( .A1(n3627), .A2(n3289), .B1(n3069), .B2(n3622), .ZN(N318)
         );
  OAI22_X1 U3372 ( .A1(n3633), .A2(n3330), .B1(n3028), .B2(n3670), .ZN(N319)
         );
  OAI22_X1 U3373 ( .A1(n3630), .A2(n3209), .B1(n3149), .B2(n3671), .ZN(N442)
         );
  OAI22_X1 U3374 ( .A1(n3742), .A2(n3195), .B1(n3136), .B2(n3459), .ZN(N312)
         );
  OAI22_X1 U3375 ( .A1(n3740), .A2(n3374), .B1(n3419), .B2(n3459), .ZN(N416)
         );
  OAI22_X1 U3376 ( .A1(n3649), .A2(n3165), .B1(n3226), .B2(n3459), .ZN(N452)
         );
  OAI22_X1 U3377 ( .A1(n3638), .A2(n3049), .B1(n3298), .B2(n3459), .ZN(N313)
         );
  OAI22_X1 U3378 ( .A1(n3739), .A2(n3178), .B1(n3075), .B2(n3459), .ZN(N315)
         );
  AND2_X1 U3379 ( .A1(n2213), .A2(n2656), .ZN(n3598) );
  INV_X1 U3380 ( .A(n2587), .ZN(n2444) );
  INV_X1 U3381 ( .A(n2770), .ZN(n2161) );
  INV_X1 U3382 ( .A(n2749), .ZN(n2131) );
  INV_X1 U3383 ( .A(n2653), .ZN(n2209) );
  INV_X1 U3384 ( .A(n2561), .ZN(n2420) );
  INV_X1 U3385 ( .A(n2807), .ZN(n2166) );
  NAND2_X1 U3386 ( .A1(n3116), .A2(n3192), .ZN(N664) );
  NAND2_X1 U3387 ( .A1(n2276), .A2(n3338), .ZN(N470) );
  INV_X1 U3388 ( .A(n2821), .ZN(n2141) );
  INV_X1 U3389 ( .A(n2726), .ZN(n2218) );
  NAND2_X1 U3390 ( .A1(n3077), .A2(n3337), .ZN(N534) );
  OAI22_X1 U3391 ( .A1(n3845), .A2(n1975), .B1(n1911), .B2(n3836), .ZN(N88) );
  OAI22_X1 U3392 ( .A1(n3845), .A2(n1974), .B1(n1910), .B2(n3836), .ZN(N89) );
  OAI22_X1 U3393 ( .A1(n3846), .A2(n1973), .B1(n1909), .B2(n3836), .ZN(N90) );
  OAI22_X1 U3394 ( .A1(n3846), .A2(n1972), .B1(n1908), .B2(n3836), .ZN(N91) );
  OAI22_X1 U3395 ( .A1(n3846), .A2(n1971), .B1(n1907), .B2(n3836), .ZN(N92) );
  OAI22_X1 U3396 ( .A1(n3843), .A2(n1970), .B1(n1906), .B2(n3836), .ZN(N93) );
  OAI22_X1 U3397 ( .A1(n3843), .A2(n1969), .B1(n1905), .B2(n3836), .ZN(N94) );
  OAI22_X1 U3398 ( .A1(n3843), .A2(n1968), .B1(n1904), .B2(n3836), .ZN(N95) );
  OAI22_X1 U3399 ( .A1(n3843), .A2(n1967), .B1(n1903), .B2(n3836), .ZN(N96) );
  OAI22_X1 U3400 ( .A1(n3843), .A2(n1966), .B1(n1902), .B2(n3836), .ZN(N97) );
  OAI22_X1 U3401 ( .A1(n3844), .A2(n1965), .B1(n1901), .B2(n3836), .ZN(N98) );
  OAI22_X1 U3402 ( .A1(n3700), .A2(n2068), .B1(n2004), .B2(n3691), .ZN(N254)
         );
  OAI22_X1 U3403 ( .A1(n3701), .A2(n2067), .B1(n2003), .B2(n3691), .ZN(N255)
         );
  OAI22_X1 U3404 ( .A1(n3701), .A2(n2066), .B1(n2002), .B2(n3691), .ZN(N256)
         );
  OAI22_X1 U3405 ( .A1(n3701), .A2(n2065), .B1(n2001), .B2(n3691), .ZN(N257)
         );
  OAI22_X1 U3406 ( .A1(n3701), .A2(n2064), .B1(n2000), .B2(n3691), .ZN(N258)
         );
  OAI22_X1 U3407 ( .A1(n3698), .A2(n2063), .B1(n1999), .B2(n3691), .ZN(N259)
         );
  OAI22_X1 U3408 ( .A1(n3698), .A2(n2062), .B1(n1998), .B2(n3691), .ZN(N260)
         );
  OAI22_X1 U3409 ( .A1(n3698), .A2(n2061), .B1(n1997), .B2(n3691), .ZN(N261)
         );
  OAI22_X1 U3410 ( .A1(n3698), .A2(n2060), .B1(n1996), .B2(n3691), .ZN(N262)
         );
  OAI22_X1 U3411 ( .A1(n3698), .A2(n2059), .B1(n1995), .B2(n3691), .ZN(N263)
         );
  OAI22_X1 U3412 ( .A1(n3699), .A2(n2058), .B1(n1994), .B2(n3691), .ZN(N264)
         );
  OAI22_X1 U3413 ( .A1(n3699), .A2(n2057), .B1(n1993), .B2(n3691), .ZN(N265)
         );
  OAI22_X1 U3414 ( .A1(n3866), .A2(n1925), .B1(n1989), .B2(n3836), .ZN(N10) );
  OAI22_X1 U3415 ( .A1(n3721), .A2(n2055), .B1(n2832), .B2(n2119), .ZN(N139)
         );
  OAI22_X1 U3416 ( .A1(n3846), .A2(n1926), .B1(n2543), .B2(n1990), .ZN(N9) );
  OAI22_X1 U3417 ( .A1(n3866), .A2(n1963), .B1(n1899), .B2(n2543), .ZN(N100)
         );
  OAI22_X1 U3418 ( .A1(n3866), .A2(n1962), .B1(n1898), .B2(n2543), .ZN(N101)
         );
  OAI22_X1 U3419 ( .A1(n3866), .A2(n1961), .B1(n1897), .B2(n2543), .ZN(N102)
         );
  OAI22_X1 U3420 ( .A1(n3866), .A2(n1960), .B1(n1896), .B2(n2543), .ZN(N103)
         );
  OAI22_X1 U3421 ( .A1(n3867), .A2(n1959), .B1(n1895), .B2(n2543), .ZN(N104)
         );
  OAI22_X1 U3422 ( .A1(n3867), .A2(n1957), .B1(n1893), .B2(n2543), .ZN(N106)
         );
  OAI22_X1 U3423 ( .A1(n3721), .A2(n2054), .B1(n2118), .B2(n2832), .ZN(N140)
         );
  OAI22_X1 U3424 ( .A1(n3721), .A2(n2053), .B1(n2117), .B2(n2832), .ZN(N141)
         );
  OAI22_X1 U3425 ( .A1(n3721), .A2(n2052), .B1(n2116), .B2(n2832), .ZN(N142)
         );
  OAI22_X1 U3426 ( .A1(n3721), .A2(n2051), .B1(n2115), .B2(n2832), .ZN(N143)
         );
  OAI22_X1 U3427 ( .A1(n3722), .A2(n2050), .B1(n2114), .B2(n2832), .ZN(N144)
         );
  OAI22_X1 U3428 ( .A1(n3722), .A2(n2049), .B1(n2113), .B2(n2832), .ZN(N145)
         );
  OAI22_X1 U3429 ( .A1(n3847), .A2(n1990), .B1(n1926), .B2(n3838), .ZN(N73) );
  OAI22_X1 U3430 ( .A1(n3847), .A2(n1989), .B1(n1925), .B2(n3838), .ZN(N74) );
  OAI22_X1 U3431 ( .A1(n3847), .A2(n1988), .B1(n1924), .B2(n3838), .ZN(N75) );
  OAI22_X1 U3432 ( .A1(n3848), .A2(n1987), .B1(n1923), .B2(n3837), .ZN(N76) );
  OAI22_X1 U3433 ( .A1(n3848), .A2(n1986), .B1(n1922), .B2(n3837), .ZN(N77) );
  OAI22_X1 U3434 ( .A1(n3848), .A2(n1985), .B1(n1921), .B2(n3837), .ZN(N78) );
  OAI22_X1 U3435 ( .A1(n3848), .A2(n1984), .B1(n1920), .B2(n3837), .ZN(N79) );
  OAI22_X1 U3436 ( .A1(n3848), .A2(n1983), .B1(n1919), .B2(n3837), .ZN(N80) );
  OAI22_X1 U3437 ( .A1(n3849), .A2(n1982), .B1(n1918), .B2(n3837), .ZN(N81) );
  OAI22_X1 U3438 ( .A1(n3844), .A2(n1981), .B1(n1917), .B2(n3837), .ZN(N82) );
  OAI22_X1 U3439 ( .A1(n3844), .A2(n1980), .B1(n1916), .B2(n3837), .ZN(N83) );
  OAI22_X1 U3440 ( .A1(n3844), .A2(n1979), .B1(n1915), .B2(n3837), .ZN(N84) );
  OAI22_X1 U3441 ( .A1(n3845), .A2(n1978), .B1(n1914), .B2(n3837), .ZN(N85) );
  OAI22_X1 U3442 ( .A1(n3845), .A2(n1977), .B1(n1913), .B2(n3837), .ZN(N86) );
  OAI22_X1 U3443 ( .A1(n3845), .A2(n1976), .B1(n1912), .B2(n3837), .ZN(N87) );
  OAI22_X1 U3444 ( .A1(n3710), .A2(n2116), .B1(n2052), .B2(n3695), .ZN(N206)
         );
  OAI22_X1 U3445 ( .A1(n3710), .A2(n2115), .B1(n2051), .B2(n3695), .ZN(N207)
         );
  OAI22_X1 U3446 ( .A1(n3710), .A2(n2114), .B1(n2050), .B2(n3695), .ZN(N208)
         );
  OAI22_X1 U3447 ( .A1(n3711), .A2(n2113), .B1(n2049), .B2(n3695), .ZN(N209)
         );
  OAI22_X1 U3448 ( .A1(n3711), .A2(n2112), .B1(n2048), .B2(n3695), .ZN(N210)
         );
  OAI22_X1 U3449 ( .A1(n3706), .A2(n2111), .B1(n2047), .B2(n3695), .ZN(N211)
         );
  OAI22_X1 U3450 ( .A1(n3706), .A2(n2110), .B1(n2046), .B2(n3695), .ZN(N212)
         );
  OAI22_X1 U3451 ( .A1(n3707), .A2(n2109), .B1(n2045), .B2(n3695), .ZN(N213)
         );
  OAI22_X1 U3452 ( .A1(n3707), .A2(n2108), .B1(n2044), .B2(n3695), .ZN(N214)
         );
  OAI22_X1 U3453 ( .A1(n3707), .A2(n2107), .B1(n2043), .B2(n3695), .ZN(N215)
         );
  OAI22_X1 U3454 ( .A1(n3707), .A2(n2106), .B1(n2042), .B2(n3695), .ZN(N216)
         );
  OAI22_X1 U3455 ( .A1(n3707), .A2(n2105), .B1(n2041), .B2(n3695), .ZN(N217)
         );
  OAI22_X1 U3456 ( .A1(n3708), .A2(n2104), .B1(n2040), .B2(n3694), .ZN(N218)
         );
  OAI22_X1 U3457 ( .A1(n3708), .A2(n2103), .B1(n2039), .B2(n3694), .ZN(N219)
         );
  OAI22_X1 U3458 ( .A1(n3708), .A2(n2102), .B1(n2038), .B2(n3694), .ZN(N220)
         );
  OAI22_X1 U3459 ( .A1(n3708), .A2(n2101), .B1(n2037), .B2(n3694), .ZN(N221)
         );
  OAI22_X1 U3460 ( .A1(n3708), .A2(n2100), .B1(n2036), .B2(n3694), .ZN(N222)
         );
  OAI22_X1 U3461 ( .A1(n3704), .A2(n2099), .B1(n2035), .B2(n3694), .ZN(N223)
         );
  OAI22_X1 U3462 ( .A1(n3704), .A2(n2098), .B1(n2034), .B2(n3694), .ZN(N224)
         );
  OAI22_X1 U3463 ( .A1(n3704), .A2(n2097), .B1(n2033), .B2(n3694), .ZN(N225)
         );
  OAI22_X1 U3464 ( .A1(n3704), .A2(n2096), .B1(n2032), .B2(n3694), .ZN(N226)
         );
  OAI22_X1 U3465 ( .A1(n3705), .A2(n2095), .B1(n2031), .B2(n3694), .ZN(N227)
         );
  OAI22_X1 U3466 ( .A1(n3705), .A2(n2094), .B1(n2030), .B2(n3694), .ZN(N228)
         );
  OAI22_X1 U3467 ( .A1(n3705), .A2(n2093), .B1(n2029), .B2(n3694), .ZN(N229)
         );
  OAI22_X1 U3468 ( .A1(n3705), .A2(n2092), .B1(n2028), .B2(n3693), .ZN(N230)
         );
  OAI22_X1 U3469 ( .A1(n3705), .A2(n2091), .B1(n2027), .B2(n3693), .ZN(N231)
         );
  OAI22_X1 U3470 ( .A1(n3706), .A2(n2090), .B1(n2026), .B2(n3693), .ZN(N232)
         );
  OAI22_X1 U3471 ( .A1(n3706), .A2(n2089), .B1(n2025), .B2(n3693), .ZN(N233)
         );
  OAI22_X1 U3472 ( .A1(n3706), .A2(n2088), .B1(n2024), .B2(n3693), .ZN(N234)
         );
  OAI22_X1 U3473 ( .A1(n3701), .A2(n2087), .B1(n2023), .B2(n3693), .ZN(N235)
         );
  OAI22_X1 U3474 ( .A1(n3702), .A2(n2086), .B1(n2022), .B2(n3693), .ZN(N236)
         );
  OAI22_X1 U3475 ( .A1(n3702), .A2(n2085), .B1(n2021), .B2(n3693), .ZN(N237)
         );
  OAI22_X1 U3476 ( .A1(n3702), .A2(n2084), .B1(n2020), .B2(n3693), .ZN(N238)
         );
  OAI22_X1 U3477 ( .A1(n3702), .A2(n2083), .B1(n2019), .B2(n3693), .ZN(N239)
         );
  OAI22_X1 U3478 ( .A1(n3702), .A2(n2082), .B1(n2018), .B2(n3693), .ZN(N240)
         );
  OAI22_X1 U3479 ( .A1(n3703), .A2(n2081), .B1(n2017), .B2(n3693), .ZN(N241)
         );
  OAI22_X1 U3480 ( .A1(n3703), .A2(n2080), .B1(n2016), .B2(n3692), .ZN(N242)
         );
  OAI22_X1 U3481 ( .A1(n3703), .A2(n2079), .B1(n2015), .B2(n3692), .ZN(N243)
         );
  OAI22_X1 U3482 ( .A1(n3703), .A2(n2078), .B1(n2014), .B2(n3692), .ZN(N244)
         );
  OAI22_X1 U3483 ( .A1(n3703), .A2(n2077), .B1(n2013), .B2(n3692), .ZN(N245)
         );
  OAI22_X1 U3484 ( .A1(n3704), .A2(n2076), .B1(n2012), .B2(n3692), .ZN(N246)
         );
  OAI22_X1 U3485 ( .A1(n3699), .A2(n2075), .B1(n2011), .B2(n3692), .ZN(N247)
         );
  OAI22_X1 U3486 ( .A1(n3699), .A2(n2074), .B1(n2010), .B2(n3692), .ZN(N248)
         );
  OAI22_X1 U3487 ( .A1(n3699), .A2(n2073), .B1(n2009), .B2(n3692), .ZN(N249)
         );
  OAI22_X1 U3488 ( .A1(n3700), .A2(n2072), .B1(n2008), .B2(n3692), .ZN(N250)
         );
  OAI22_X1 U3489 ( .A1(n3700), .A2(n2071), .B1(n2007), .B2(n3692), .ZN(N251)
         );
  OAI22_X1 U3490 ( .A1(n3700), .A2(n2070), .B1(n2006), .B2(n3692), .ZN(N252)
         );
  OAI22_X1 U3491 ( .A1(n3700), .A2(n2069), .B1(n2005), .B2(n3692), .ZN(N253)
         );
  OAI22_X1 U3492 ( .A1(n3855), .A2(n1895), .B1(n1959), .B2(n3840), .ZN(N40) );
  OAI22_X1 U3493 ( .A1(n3855), .A2(n1894), .B1(n1958), .B2(n3840), .ZN(N41) );
  OAI22_X1 U3494 ( .A1(n3855), .A2(n1893), .B1(n1957), .B2(n3840), .ZN(N42) );
  OAI22_X1 U3495 ( .A1(n3855), .A2(n1892), .B1(n1956), .B2(n3840), .ZN(N43) );
  OAI22_X1 U3496 ( .A1(n3856), .A2(n1891), .B1(n1955), .B2(n3840), .ZN(N44) );
  OAI22_X1 U3497 ( .A1(n3856), .A2(n1890), .B1(n1954), .B2(n3840), .ZN(N45) );
  OAI22_X1 U3498 ( .A1(n3851), .A2(n1889), .B1(n1953), .B2(n3840), .ZN(N46) );
  OAI22_X1 U3499 ( .A1(n3851), .A2(n1888), .B1(n1952), .B2(n3840), .ZN(N47) );
  OAI22_X1 U3500 ( .A1(n3852), .A2(n1887), .B1(n1951), .B2(n3840), .ZN(N48) );
  OAI22_X1 U3501 ( .A1(n3852), .A2(n1886), .B1(n1950), .B2(n3840), .ZN(N49) );
  OAI22_X1 U3502 ( .A1(n3852), .A2(n1885), .B1(n1949), .B2(n3840), .ZN(N50) );
  OAI22_X1 U3503 ( .A1(n3852), .A2(n1884), .B1(n1948), .B2(n3840), .ZN(N51) );
  OAI22_X1 U3504 ( .A1(n3852), .A2(n1883), .B1(n1947), .B2(n3839), .ZN(N52) );
  OAI22_X1 U3505 ( .A1(n3853), .A2(n1882), .B1(n1946), .B2(n3839), .ZN(N53) );
  OAI22_X1 U3506 ( .A1(n3853), .A2(n1881), .B1(n1945), .B2(n3839), .ZN(N54) );
  OAI22_X1 U3507 ( .A1(n3853), .A2(n1880), .B1(n1944), .B2(n3839), .ZN(N55) );
  OAI22_X1 U3508 ( .A1(n3853), .A2(n1879), .B1(n1943), .B2(n3839), .ZN(N56) );
  OAI22_X1 U3509 ( .A1(n3853), .A2(n1878), .B1(n1942), .B2(n3839), .ZN(N57) );
  OAI22_X1 U3510 ( .A1(n3849), .A2(n1877), .B1(n1941), .B2(n3839), .ZN(N58) );
  OAI22_X1 U3511 ( .A1(n3849), .A2(n1876), .B1(n1940), .B2(n3839), .ZN(N59) );
  OAI22_X1 U3512 ( .A1(n3849), .A2(n1875), .B1(n1939), .B2(n3839), .ZN(N60) );
  OAI22_X1 U3513 ( .A1(n3849), .A2(n1874), .B1(n1938), .B2(n3839), .ZN(N61) );
  OAI22_X1 U3514 ( .A1(n3850), .A2(n1873), .B1(n1937), .B2(n3839), .ZN(N62) );
  OAI22_X1 U3515 ( .A1(n3850), .A2(n1872), .B1(n1936), .B2(n3839), .ZN(N63) );
  OAI22_X1 U3516 ( .A1(n3850), .A2(n1871), .B1(n1935), .B2(n3838), .ZN(N64) );
  OAI22_X1 U3517 ( .A1(n3850), .A2(n1870), .B1(n1934), .B2(n3838), .ZN(N65) );
  OAI22_X1 U3518 ( .A1(n3850), .A2(n1869), .B1(n1933), .B2(n3838), .ZN(N66) );
  OAI22_X1 U3519 ( .A1(n3851), .A2(n1868), .B1(n1932), .B2(n3838), .ZN(N67) );
  OAI22_X1 U3520 ( .A1(n3851), .A2(n1867), .B1(n1931), .B2(n3838), .ZN(N68) );
  OAI22_X1 U3521 ( .A1(n3851), .A2(n1866), .B1(n1930), .B2(n3838), .ZN(N69) );
  OAI22_X1 U3522 ( .A1(n3846), .A2(n1865), .B1(n1929), .B2(n3838), .ZN(N70) );
  OAI22_X1 U3523 ( .A1(n3847), .A2(n1864), .B1(n1928), .B2(n3838), .ZN(N71) );
  OAI22_X1 U3524 ( .A1(n3847), .A2(n1863), .B1(n1927), .B2(n3838), .ZN(N72) );
  OAI22_X1 U3525 ( .A1(n3844), .A2(n1964), .B1(n1900), .B2(n2543), .ZN(N99) );
  OAI22_X1 U3526 ( .A1(n3867), .A2(n1958), .B1(n1894), .B2(n3842), .ZN(N105)
         );
  OAI22_X1 U3527 ( .A1(n3867), .A2(n1956), .B1(n1892), .B2(n3842), .ZN(N107)
         );
  OAI22_X1 U3528 ( .A1(n3867), .A2(n1955), .B1(n1891), .B2(n3842), .ZN(N108)
         );
  OAI22_X1 U3529 ( .A1(n3868), .A2(n1954), .B1(n1890), .B2(n3842), .ZN(N109)
         );
  OAI22_X1 U3530 ( .A1(n3863), .A2(n1953), .B1(n1889), .B2(n3842), .ZN(N110)
         );
  OAI22_X1 U3531 ( .A1(n3863), .A2(n1952), .B1(n1888), .B2(n3842), .ZN(N111)
         );
  OAI22_X1 U3532 ( .A1(n3864), .A2(n1951), .B1(n1887), .B2(n3842), .ZN(N112)
         );
  OAI22_X1 U3533 ( .A1(n3864), .A2(n1950), .B1(n1886), .B2(n3842), .ZN(N113)
         );
  OAI22_X1 U3534 ( .A1(n3864), .A2(n1949), .B1(n1885), .B2(n3842), .ZN(N114)
         );
  OAI22_X1 U3535 ( .A1(n3864), .A2(n1948), .B1(n1884), .B2(n3842), .ZN(N115)
         );
  OAI22_X1 U3536 ( .A1(n3864), .A2(n1947), .B1(n1883), .B2(n3842), .ZN(N116)
         );
  OAI22_X1 U3537 ( .A1(n3865), .A2(n1946), .B1(n1882), .B2(n3841), .ZN(N117)
         );
  OAI22_X1 U3538 ( .A1(n3865), .A2(n1945), .B1(n1881), .B2(n3841), .ZN(N118)
         );
  OAI22_X1 U3539 ( .A1(n3865), .A2(n1944), .B1(n1880), .B2(n3841), .ZN(N119)
         );
  OAI22_X1 U3540 ( .A1(n3865), .A2(n1943), .B1(n1879), .B2(n3841), .ZN(N120)
         );
  OAI22_X1 U3541 ( .A1(n3861), .A2(n1942), .B1(n1878), .B2(n3841), .ZN(N121)
         );
  OAI22_X1 U3542 ( .A1(n3861), .A2(n1941), .B1(n1877), .B2(n3841), .ZN(N122)
         );
  OAI22_X1 U3543 ( .A1(n3861), .A2(n1940), .B1(n1876), .B2(n3841), .ZN(N123)
         );
  OAI22_X1 U3544 ( .A1(n3861), .A2(n1939), .B1(n1875), .B2(n3841), .ZN(N124)
         );
  OAI22_X1 U3545 ( .A1(n3862), .A2(n1938), .B1(n1874), .B2(n3841), .ZN(N125)
         );
  OAI22_X1 U3546 ( .A1(n3862), .A2(n1937), .B1(n1873), .B2(n3841), .ZN(N126)
         );
  OAI22_X1 U3547 ( .A1(n3862), .A2(n1936), .B1(n1872), .B2(n3841), .ZN(N127)
         );
  OAI22_X1 U3548 ( .A1(n3862), .A2(n1935), .B1(n1871), .B2(n3841), .ZN(N128)
         );
  OAI22_X1 U3549 ( .A1(n3862), .A2(n1934), .B1(n1870), .B2(n3837), .ZN(N129)
         );
  OAI22_X1 U3550 ( .A1(n3863), .A2(n1933), .B1(n1869), .B2(n3840), .ZN(N130)
         );
  OAI22_X1 U3551 ( .A1(n3863), .A2(n1932), .B1(n1868), .B2(n3839), .ZN(N131)
         );
  OAI22_X1 U3552 ( .A1(n3858), .A2(n1931), .B1(n1867), .B2(n3838), .ZN(N132)
         );
  OAI22_X1 U3553 ( .A1(n3859), .A2(n1930), .B1(n1866), .B2(n3836), .ZN(N133)
         );
  OAI22_X1 U3554 ( .A1(n3859), .A2(n1929), .B1(n1865), .B2(n3842), .ZN(N134)
         );
  OAI22_X1 U3555 ( .A1(n3859), .A2(n1928), .B1(n1864), .B2(n3841), .ZN(N135)
         );
  OAI22_X1 U3556 ( .A1(n3722), .A2(n2048), .B1(n2112), .B2(n3697), .ZN(N146)
         );
  OAI22_X1 U3557 ( .A1(n3722), .A2(n2047), .B1(n2111), .B2(n3697), .ZN(N147)
         );
  OAI22_X1 U3558 ( .A1(n3722), .A2(n2046), .B1(n2110), .B2(n3697), .ZN(N148)
         );
  OAI22_X1 U3559 ( .A1(n3723), .A2(n2045), .B1(n2109), .B2(n3697), .ZN(N149)
         );
  OAI22_X1 U3560 ( .A1(n3723), .A2(n2044), .B1(n2108), .B2(n3697), .ZN(N150)
         );
  OAI22_X1 U3561 ( .A1(n3718), .A2(n2043), .B1(n2107), .B2(n3697), .ZN(N151)
         );
  OAI22_X1 U3562 ( .A1(n3718), .A2(n2042), .B1(n2106), .B2(n3697), .ZN(N152)
         );
  OAI22_X1 U3563 ( .A1(n3719), .A2(n2041), .B1(n2105), .B2(n3697), .ZN(N153)
         );
  OAI22_X1 U3564 ( .A1(n3719), .A2(n2040), .B1(n2104), .B2(n3697), .ZN(N154)
         );
  OAI22_X1 U3565 ( .A1(n3719), .A2(n2039), .B1(n2103), .B2(n3697), .ZN(N155)
         );
  OAI22_X1 U3566 ( .A1(n3719), .A2(n2038), .B1(n2102), .B2(n3697), .ZN(N156)
         );
  OAI22_X1 U3567 ( .A1(n3719), .A2(n2037), .B1(n2101), .B2(n3697), .ZN(N157)
         );
  OAI22_X1 U3568 ( .A1(n3720), .A2(n2036), .B1(n2100), .B2(n3696), .ZN(N158)
         );
  OAI22_X1 U3569 ( .A1(n3720), .A2(n2035), .B1(n2099), .B2(n3696), .ZN(N159)
         );
  OAI22_X1 U3570 ( .A1(n3720), .A2(n2034), .B1(n2098), .B2(n3696), .ZN(N160)
         );
  OAI22_X1 U3571 ( .A1(n3720), .A2(n2033), .B1(n2097), .B2(n3696), .ZN(N161)
         );
  OAI22_X1 U3572 ( .A1(n3720), .A2(n2032), .B1(n2096), .B2(n3696), .ZN(N162)
         );
  OAI22_X1 U3573 ( .A1(n3716), .A2(n2031), .B1(n2095), .B2(n3696), .ZN(N163)
         );
  OAI22_X1 U3574 ( .A1(n3716), .A2(n2030), .B1(n2094), .B2(n3696), .ZN(N164)
         );
  OAI22_X1 U3575 ( .A1(n3716), .A2(n2029), .B1(n2093), .B2(n3696), .ZN(N165)
         );
  OAI22_X1 U3576 ( .A1(n3716), .A2(n2028), .B1(n2092), .B2(n3696), .ZN(N166)
         );
  OAI22_X1 U3577 ( .A1(n3717), .A2(n2027), .B1(n2091), .B2(n3696), .ZN(N167)
         );
  OAI22_X1 U3578 ( .A1(n3717), .A2(n2026), .B1(n2090), .B2(n3696), .ZN(N168)
         );
  OAI22_X1 U3579 ( .A1(n3717), .A2(n2025), .B1(n2089), .B2(n3696), .ZN(N169)
         );
  OAI22_X1 U3580 ( .A1(n3717), .A2(n2024), .B1(n2088), .B2(n3696), .ZN(N170)
         );
  OAI22_X1 U3581 ( .A1(n3717), .A2(n2023), .B1(n2087), .B2(n3695), .ZN(N171)
         );
  OAI22_X1 U3582 ( .A1(n3718), .A2(n2022), .B1(n2086), .B2(n3694), .ZN(N172)
         );
  OAI22_X1 U3583 ( .A1(n3718), .A2(n2021), .B1(n2085), .B2(n3693), .ZN(N173)
         );
  OAI22_X1 U3584 ( .A1(n3718), .A2(n2020), .B1(n2084), .B2(n3692), .ZN(N174)
         );
  OAI22_X1 U3585 ( .A1(n3713), .A2(n2019), .B1(n2083), .B2(n3691), .ZN(N175)
         );
  OAI22_X1 U3586 ( .A1(n3714), .A2(n2018), .B1(n2082), .B2(n3697), .ZN(N176)
         );
  OAI22_X1 U3587 ( .A1(n3714), .A2(n2017), .B1(n2081), .B2(n3696), .ZN(N177)
         );
  OAI22_X1 U3588 ( .A1(n3714), .A2(n2016), .B1(n2080), .B2(n3695), .ZN(N178)
         );
  OAI22_X1 U3589 ( .A1(n3714), .A2(n2015), .B1(n2079), .B2(n3694), .ZN(N179)
         );
  OAI22_X1 U3590 ( .A1(n3714), .A2(n2014), .B1(n2078), .B2(n3693), .ZN(N180)
         );
  OAI22_X1 U3591 ( .A1(n3715), .A2(n2013), .B1(n2077), .B2(n3692), .ZN(N181)
         );
  OAI22_X1 U3592 ( .A1(n3715), .A2(n2012), .B1(n2076), .B2(n3695), .ZN(N182)
         );
  OAI22_X1 U3593 ( .A1(n3715), .A2(n2011), .B1(n2075), .B2(n3694), .ZN(N183)
         );
  OAI22_X1 U3594 ( .A1(n3715), .A2(n2010), .B1(n2074), .B2(n3693), .ZN(N184)
         );
  OAI22_X1 U3595 ( .A1(n3715), .A2(n2009), .B1(n2073), .B2(n3692), .ZN(N185)
         );
  OAI22_X1 U3596 ( .A1(n3716), .A2(n2008), .B1(n2072), .B2(n3691), .ZN(N186)
         );
  OAI22_X1 U3597 ( .A1(n3711), .A2(n2007), .B1(n2071), .B2(n3697), .ZN(N187)
         );
  OAI22_X1 U3598 ( .A1(n3711), .A2(n2006), .B1(n2070), .B2(n3696), .ZN(N188)
         );
  OAI22_X1 U3599 ( .A1(n3711), .A2(n2005), .B1(n2069), .B2(n3691), .ZN(N189)
         );
  OAI22_X1 U3600 ( .A1(n3712), .A2(n2004), .B1(n2068), .B2(n3695), .ZN(N190)
         );
  OAI22_X1 U3601 ( .A1(n3712), .A2(n2003), .B1(n2067), .B2(n3694), .ZN(N191)
         );
  OAI22_X1 U3602 ( .A1(n3712), .A2(n2002), .B1(n2066), .B2(n3693), .ZN(N192)
         );
  OAI22_X1 U3603 ( .A1(n3712), .A2(n2001), .B1(n2065), .B2(n3692), .ZN(N193)
         );
  OAI22_X1 U3604 ( .A1(n3712), .A2(n2000), .B1(n2064), .B2(n2832), .ZN(N194)
         );
  OAI22_X1 U3605 ( .A1(n3713), .A2(n1999), .B1(n2063), .B2(n2832), .ZN(N195)
         );
  OAI22_X1 U3606 ( .A1(n3713), .A2(n1998), .B1(n2062), .B2(n2832), .ZN(N196)
         );
  OAI22_X1 U3607 ( .A1(n3713), .A2(n1997), .B1(n2061), .B2(n2832), .ZN(N197)
         );
  OAI22_X1 U3608 ( .A1(n3713), .A2(n1996), .B1(n2060), .B2(n3695), .ZN(N198)
         );
  OAI22_X1 U3609 ( .A1(n3709), .A2(n1995), .B1(n2059), .B2(n3694), .ZN(N199)
         );
  OAI22_X1 U3610 ( .A1(n3709), .A2(n1994), .B1(n2058), .B2(n3693), .ZN(N200)
         );
  OAI22_X1 U3611 ( .A1(n3709), .A2(n1993), .B1(n2057), .B2(n3692), .ZN(N201)
         );
  OAI22_X1 U3612 ( .A1(n3709), .A2(n1992), .B1(n2056), .B2(n3691), .ZN(N202)
         );
  OAI22_X1 U3613 ( .A1(n3709), .A2(n2119), .B1(n2055), .B2(n3697), .ZN(N203)
         );
  OAI22_X1 U3614 ( .A1(n3710), .A2(n2118), .B1(n2054), .B2(n3696), .ZN(N204)
         );
  OAI22_X1 U3615 ( .A1(n3710), .A2(n2117), .B1(n2053), .B2(n3697), .ZN(N205)
         );
  OAI22_X1 U3616 ( .A1(n3868), .A2(n1924), .B1(n1988), .B2(n3842), .ZN(N11) );
  OAI22_X1 U3617 ( .A1(n3865), .A2(n1923), .B1(n1987), .B2(n3841), .ZN(N12) );
  OAI22_X1 U3618 ( .A1(n3863), .A2(n1922), .B1(n1986), .B2(n3837), .ZN(N13) );
  OAI22_X1 U3619 ( .A1(n3859), .A2(n1921), .B1(n1985), .B2(n3840), .ZN(N14) );
  OAI22_X1 U3620 ( .A1(n3859), .A2(n1920), .B1(n1984), .B2(n3839), .ZN(N15) );
  OAI22_X1 U3621 ( .A1(n3860), .A2(n1919), .B1(n1983), .B2(n3838), .ZN(N16) );
  OAI22_X1 U3622 ( .A1(n3860), .A2(n1918), .B1(n1982), .B2(n3837), .ZN(N17) );
  OAI22_X1 U3623 ( .A1(n3860), .A2(n1917), .B1(n1981), .B2(n3840), .ZN(N18) );
  OAI22_X1 U3624 ( .A1(n3860), .A2(n1916), .B1(n1980), .B2(n3839), .ZN(N19) );
  OAI22_X1 U3625 ( .A1(n3860), .A2(n1915), .B1(n1979), .B2(n3838), .ZN(N20) );
  OAI22_X1 U3626 ( .A1(n3861), .A2(n1914), .B1(n1978), .B2(n3836), .ZN(N21) );
  OAI22_X1 U3627 ( .A1(n3856), .A2(n1913), .B1(n1977), .B2(n3842), .ZN(N22) );
  OAI22_X1 U3628 ( .A1(n3856), .A2(n1912), .B1(n1976), .B2(n3841), .ZN(N23) );
  OAI22_X1 U3629 ( .A1(n3856), .A2(n1911), .B1(n1975), .B2(n3836), .ZN(N24) );
  OAI22_X1 U3630 ( .A1(n3857), .A2(n1910), .B1(n1974), .B2(n3837), .ZN(N25) );
  OAI22_X1 U3631 ( .A1(n3857), .A2(n1909), .B1(n1973), .B2(n3840), .ZN(N26) );
  OAI22_X1 U3632 ( .A1(n3857), .A2(n1908), .B1(n1972), .B2(n3839), .ZN(N27) );
  OAI22_X1 U3633 ( .A1(n3857), .A2(n1907), .B1(n1971), .B2(n3838), .ZN(N28) );
  OAI22_X1 U3634 ( .A1(n3857), .A2(n1906), .B1(n1970), .B2(n2543), .ZN(N29) );
  OAI22_X1 U3635 ( .A1(n3858), .A2(n1905), .B1(n1969), .B2(n2543), .ZN(N30) );
  OAI22_X1 U3636 ( .A1(n3858), .A2(n1904), .B1(n1968), .B2(n2543), .ZN(N31) );
  OAI22_X1 U3637 ( .A1(n3858), .A2(n1903), .B1(n1967), .B2(n3837), .ZN(N32) );
  OAI22_X1 U3638 ( .A1(n3858), .A2(n1902), .B1(n1966), .B2(n3840), .ZN(N33) );
  OAI22_X1 U3639 ( .A1(n3854), .A2(n1901), .B1(n1965), .B2(n3839), .ZN(N34) );
  OAI22_X1 U3640 ( .A1(n3854), .A2(n1900), .B1(n1964), .B2(n3838), .ZN(N35) );
  OAI22_X1 U3641 ( .A1(n3854), .A2(n1899), .B1(n1963), .B2(n3836), .ZN(N36) );
  OAI22_X1 U3642 ( .A1(n3854), .A2(n1898), .B1(n1962), .B2(n3842), .ZN(N37) );
  OAI22_X1 U3643 ( .A1(n3854), .A2(n1897), .B1(n1961), .B2(n3841), .ZN(N38) );
  OAI22_X1 U3644 ( .A1(n3855), .A2(n1896), .B1(n1960), .B2(n3842), .ZN(N39) );
  NAND2_X1 U3645 ( .A1(n1927), .A2(n1863), .ZN(N136) );
  NAND2_X1 U3646 ( .A1(n2056), .A2(n1992), .ZN(N266) );
  INV_X1 U3647 ( .A(n2832), .ZN(n3734) );
  INV_X1 U3648 ( .A(n2543), .ZN(n3879) );
  OAI22_X1 U3649 ( .A1(rC2[16]), .A2(n3223), .B1(rC2[15]), .B2(n3464), .ZN(
        n2692) );
  OAI22_X1 U3650 ( .A1(rC2[18]), .A2(n3012), .B1(rC2[17]), .B2(n3085), .ZN(
        n2690) );
  OAI211_X1 U3651 ( .C1(rC4[25]), .C2(n3170), .A(n2680), .B(n2684), .ZN(n2682)
         );
  AOI21_X1 U3652 ( .B1(rC2[24]), .B2(n3059), .A(n2685), .ZN(n2684) );
  INV_X1 U3653 ( .A(n2681), .ZN(n2248) );
  NAND2_X1 U3654 ( .A1(n2617), .A2(n2604), .ZN(n2627) );
  INV_X1 U3655 ( .A(n2680), .ZN(n2244) );
  AOI221_X1 U3656 ( .B1(n3038), .B2(rC7[61]), .C1(n3053), .C2(rC7[62]), .A(
        n2551), .ZN(n2547) );
  AOI221_X1 U3657 ( .B1(n3044), .B2(rC1[56]), .C1(n3137), .C2(rC1[57]), .A(
        n2738), .ZN(n2742) );
  AOI221_X1 U3658 ( .B1(n3089), .B2(rC6[33]), .C1(n3009), .C2(rC6[32]), .A(
        n2577), .ZN(n2581) );
  AOI221_X1 U3659 ( .B1(n3043), .B2(rC1[32]), .C1(n3136), .C2(rC1[33]), .A(
        n2760), .ZN(n2764) );
  OAI22_X1 U3660 ( .A1(rC4[41]), .A2(n3041), .B1(rC4[40]), .B2(n3158), .ZN(
        n2662) );
  INV_X1 U3661 ( .A(n2722), .ZN(n2225) );
  AOI22_X1 U3662 ( .A1(rC1[40]), .A2(n3028), .B1(rC1[41]), .B2(n3143), .ZN(
        n2755) );
  INV_X1 U3663 ( .A(n2758), .ZN(n2148) );
  AOI211_X1 U3664 ( .C1(n3190), .C2(rC2[37]), .A(n2669), .B(n2232), .ZN(n2663)
         );
  INV_X1 U3665 ( .A(n2719), .ZN(n2232) );
  AOI211_X1 U3666 ( .C1(rC2[36]), .C2(n3177), .A(n2720), .B(n2721), .ZN(n2719)
         );
  AOI211_X1 U3667 ( .C1(rC4[36]), .C2(n3017), .A(n3088), .B(rC4[35]), .ZN(
        n2720) );
  OAI222_X1 U3668 ( .A1(rC7[54]), .A2(n3135), .B1(n2637), .B2(n2559), .C1(
        rC7[55]), .C2(n3213), .ZN(n2555) );
  AOI22_X1 U3669 ( .A1(rC6[52]), .A2(n3098), .B1(rC6[53]), .B2(n3026), .ZN(
        n2637) );
  INV_X1 U3670 ( .A(n2717), .ZN(n2240) );
  OAI221_X1 U3671 ( .B1(n3122), .B2(rC2[27]), .C1(n3244), .C2(rC2[28]), .A(
        n2672), .ZN(n2717) );
  OAI211_X1 U3672 ( .C1(rC1[18]), .C2(n3013), .A(n3084), .B(rC1[17]), .ZN(
        n2778) );
  NOR3_X1 U3673 ( .A1(n3052), .A2(rC3[16]), .A3(n2783), .ZN(n2782) );
  AOI221_X1 U3674 ( .B1(rC4[57]), .B2(n3196), .C1(rC4[58]), .C2(n3050), .A(
        n2736), .ZN(n2641) );
  AOI221_X1 U3675 ( .B1(rC3[57]), .B2(n3197), .C1(rC3[58]), .C2(n3051), .A(
        n2831), .ZN(n2737) );
  OAI22_X1 U3676 ( .A1(rC1[56]), .A2(n3044), .B1(rC1[55]), .B2(n3155), .ZN(
        n2743) );
  AOI222_X1 U3677 ( .A1(rC2[31]), .A2(n3104), .B1(n2672), .B2(n2673), .C1(
        rC2[30]), .C2(n3220), .ZN(n2666) );
  OAI22_X1 U3678 ( .A1(rC4[29]), .A2(n3042), .B1(rC4[28]), .B2(n3159), .ZN(
        n2673) );
  AOI222_X1 U3679 ( .A1(rC6[43]), .A2(n3097), .B1(n2574), .B2(n2575), .C1(
        rC6[42]), .C2(n3200), .ZN(n2573) );
  OAI22_X1 U3680 ( .A1(rC7[41]), .A2(n3036), .B1(rC7[40]), .B2(n3129), .ZN(
        n2575) );
  AOI222_X1 U3681 ( .A1(rC6[49]), .A2(n3096), .B1(n2566), .B2(n2567), .C1(
        rC6[48]), .C2(n3199), .ZN(n2565) );
  OAI22_X1 U3682 ( .A1(rC7[47]), .A2(n3035), .B1(rC7[46]), .B2(n3124), .ZN(
        n2567) );
  OAI221_X1 U3683 ( .B1(rC4[32]), .B2(n3086), .C1(rC4[33]), .C2(n3225), .A(
        n2663), .ZN(n2671) );
  OAI221_X1 U3684 ( .B1(rC3[44]), .B2(n3162), .C1(rC3[45]), .C2(n3226), .A(
        n2818), .ZN(n2754) );
  OAI22_X1 U3685 ( .A1(rC2[60]), .A2(n3010), .B1(rC2[59]), .B2(n3082), .ZN(
        n2736) );
  OAI22_X1 U3686 ( .A1(rC1[60]), .A2(n3011), .B1(rC1[59]), .B2(n3083), .ZN(
        n2831) );
  OAI22_X1 U3687 ( .A1(rC1[36]), .A2(n3075), .B1(rC1[35]), .B2(n3209), .ZN(
        n2816) );
  OAI22_X1 U3688 ( .A1(rC1[18]), .A2(n3013), .B1(rC1[17]), .B2(n3084), .ZN(
        n2783) );
  OAI22_X1 U3689 ( .A1(rC1[24]), .A2(n3076), .B1(rC1[23]), .B2(n3210), .ZN(
        n2811) );
  AOI21_X1 U3690 ( .B1(rC6[36]), .B2(n3055), .A(n2634), .ZN(n2633) );
  OAI22_X1 U3691 ( .A1(rC4[39]), .A2(n3224), .B1(rC4[38]), .B2(n3032), .ZN(
        n2669) );
  OAI22_X1 U3692 ( .A1(rC1[6]), .A2(n3248), .B1(rC1[5]), .B2(n3033), .ZN(n2801) );
  AOI21_X1 U3693 ( .B1(rC3[4]), .B2(n3185), .A(n2801), .ZN(n2796) );
  OAI22_X1 U3694 ( .A1(rC3[6]), .A2(n3167), .B1(n2800), .B2(n2801), .ZN(n2798)
         );
  OAI22_X1 U3695 ( .A1(rC1[44]), .A2(n3221), .B1(rC1[43]), .B2(n3068), .ZN(
        n2750) );
  INV_X1 U3696 ( .A(n2754), .ZN(n2135) );
  OAI222_X1 U3697 ( .A1(rC3[54]), .A2(n3073), .B1(n2748), .B2(n2131), .C1(
        rC3[55]), .C2(n3240), .ZN(n2747) );
  INV_X1 U3698 ( .A(n2742), .ZN(n2122) );
  AOI221_X1 U3699 ( .B1(n2818), .B2(n2819), .C1(rC3[51]), .C2(n3056), .A(n2820), .ZN(n2745) );
  OAI222_X1 U3700 ( .A1(rC4[54]), .A2(n3074), .B1(n2652), .B2(n2209), .C1(
        rC4[55]), .C2(n3239), .ZN(n2651) );
  INV_X1 U3701 ( .A(n2646), .ZN(n2198) );
  AOI221_X1 U3702 ( .B1(n2723), .B2(n2724), .C1(rC4[51]), .C2(n3057), .A(n2725), .ZN(n2649) );
  OAI221_X1 U3703 ( .B1(rC4[44]), .B2(n3163), .C1(rC4[45]), .C2(n3227), .A(
        n2723), .ZN(n2659) );
  OAI221_X1 U3704 ( .B1(n3121), .B2(rC2[39]), .C1(n3243), .C2(rC2[40]), .A(
        n2661), .ZN(n2722) );
  AOI221_X1 U3705 ( .B1(rC3[15]), .B2(n3370), .C1(rC3[16]), .C2(n3052), .A(
        n2783), .ZN(n2780) );
  OAI221_X1 U3706 ( .B1(rC1[45]), .B2(n3165), .C1(rC1[46]), .C2(n3232), .A(
        n2821), .ZN(n2819) );
  OAI221_X1 U3707 ( .B1(rC2[45]), .B2(n3166), .C1(rC2[46]), .C2(n3233), .A(
        n2726), .ZN(n2724) );
  AOI221_X1 U3708 ( .B1(rC3[33]), .B2(n3195), .C1(rC3[34]), .C2(n3049), .A(
        n2816), .ZN(n2759) );
  OAI222_X1 U3709 ( .A1(rC3[30]), .A2(n3072), .B1(n2812), .B2(n2161), .C1(
        rC3[31]), .C2(n3238), .ZN(n2761) );
  AOI22_X1 U3710 ( .A1(n2764), .A2(n2765), .B1(n2766), .B2(n2767), .ZN(n2763)
         );
  OAI222_X1 U3711 ( .A1(rC7[30]), .A2(n3063), .B1(n2632), .B2(n2444), .C1(
        rC7[31]), .C2(n3214), .ZN(n2578) );
  AOI221_X1 U3712 ( .B1(rC7[33]), .B2(n3179), .C1(rC7[34]), .C2(n3015), .A(
        n2436), .ZN(n2576) );
  AOI22_X1 U3713 ( .A1(n2581), .A2(n2582), .B1(n2583), .B2(n2584), .ZN(n2580)
         );
  AOI22_X1 U3714 ( .A1(rC7[43]), .A2(n3174), .B1(rC7[44]), .B2(n3039), .ZN(
        n2568) );
  INV_X1 U3715 ( .A(n2569), .ZN(n2427) );
  OAI22_X1 U3716 ( .A1(rC7[57]), .A2(n3024), .B1(rC7[56]), .B2(n3123), .ZN(
        n2557) );
  OAI22_X1 U3717 ( .A1(rC7[51]), .A2(n3160), .B1(rC7[50]), .B2(n3027), .ZN(
        n2561) );
  OAI22_X1 U3718 ( .A1(rC7[45]), .A2(n3161), .B1(rC7[44]), .B2(n3039), .ZN(
        n2569) );
  OAI22_X1 U3719 ( .A1(rC7[27]), .A2(n3148), .B1(rC7[26]), .B2(n3025), .ZN(
        n2589) );
  OAI22_X1 U3720 ( .A1(rC6[54]), .A2(n3216), .B1(rC6[53]), .B2(n3026), .ZN(
        n2559) );
  AOI22_X1 U3721 ( .A1(n3063), .A2(rC7[30]), .B1(n3208), .B2(rC7[29]), .ZN(
        n2587) );
  AOI22_X1 U3722 ( .A1(n3078), .A2(rC3[42]), .B1(n3228), .B2(rC3[41]), .ZN(
        n2758) );
  AOI22_X1 U3723 ( .A1(n3072), .A2(rC3[30]), .B1(n3229), .B2(rC3[29]), .ZN(
        n2770) );
  AOI22_X1 U3724 ( .A1(n3099), .A2(rC7[18]), .B1(n3046), .B2(rC7[17]), .ZN(
        n2599) );
  AOI22_X1 U3725 ( .A1(n3007), .A2(rC1[27]), .B1(n3168), .B2(rC1[26]), .ZN(
        n2807) );
  AOI22_X1 U3726 ( .A1(n3110), .A2(rC4[30]), .B1(n3042), .B2(rC4[29]), .ZN(
        n2672) );
  AOI22_X1 U3727 ( .A1(n3101), .A2(rC7[42]), .B1(n3036), .B2(rC7[41]), .ZN(
        n2574) );
  AOI22_X1 U3728 ( .A1(n3073), .A2(rC3[54]), .B1(n3230), .B2(rC3[53]), .ZN(
        n2749) );
  AOI22_X1 U3729 ( .A1(n3074), .A2(rC4[54]), .B1(n3231), .B2(rC4[53]), .ZN(
        n2653) );
  AOI22_X1 U3730 ( .A1(n3109), .A2(rC4[6]), .B1(n3047), .B2(rC4[5]), .ZN(n2711) );
  AOI22_X1 U3731 ( .A1(n3069), .A2(rC1[39]), .B1(n3040), .B2(rC1[38]), .ZN(
        n2766) );
  AOI22_X1 U3732 ( .A1(n3100), .A2(rC7[48]), .B1(n3035), .B2(rC7[47]), .ZN(
        n2566) );
  OAI221_X1 U3733 ( .B1(rC2[21]), .B2(n3034), .C1(rC2[22]), .C2(n3234), .A(
        n2681), .ZN(n2677) );
  OAI221_X1 U3734 ( .B1(rC2[33]), .B2(n3164), .C1(rC2[34]), .C2(n3048), .A(
        n2718), .ZN(n2664) );
  OAI221_X1 U3735 ( .B1(rC1[39]), .B2(n3069), .C1(rC1[40]), .C2(n3028), .A(
        n2758), .ZN(n2757) );
  OAI221_X1 U3736 ( .B1(rC6[39]), .B2(n3062), .C1(rC6[40]), .C2(n3205), .A(
        n2574), .ZN(n2572) );
  OAI221_X1 U3737 ( .B1(rC6[10]), .B2(n3186), .C1(rC6[9]), .C2(n3064), .A(
        n2608), .ZN(n2607) );
  AOI21_X1 U3738 ( .B1(n3021), .B2(rC3[47]), .A(n2824), .ZN(n2821) );
  AOI21_X1 U3739 ( .B1(n3022), .B2(rC4[47]), .A(n2729), .ZN(n2726) );
  AOI21_X1 U3740 ( .B1(n3023), .B2(rC4[23]), .A(n2686), .ZN(n2681) );
  OAI22_X1 U3741 ( .A1(rC7[17]), .A2(n3046), .B1(rC7[16]), .B2(n3127), .ZN(
        n2600) );
  OAI22_X1 U3742 ( .A1(rC6[32]), .A2(n3009), .B1(rC6[31]), .B2(n3126), .ZN(
        n2582) );
  OAI22_X1 U3743 ( .A1(rC4[5]), .A2(n3047), .B1(rC4[4]), .B2(n3152), .ZN(n2712) );
  OAI22_X1 U3744 ( .A1(rC1[32]), .A2(n3043), .B1(rC1[31]), .B2(n3154), .ZN(
        n2765) );
  OAI22_X1 U3745 ( .A1(rC6[38]), .A2(n3037), .B1(rC6[37]), .B2(n3134), .ZN(
        n2584) );
  OAI22_X1 U3746 ( .A1(rC1[38]), .A2(n3040), .B1(rC1[37]), .B2(n3153), .ZN(
        n2767) );
  AOI22_X1 U3747 ( .A1(n3017), .A2(rC4[36]), .B1(n3088), .B2(rC4[35]), .ZN(
        n2718) );
  AOI21_X1 U3748 ( .B1(n3066), .B2(rC2[26]), .A(n2679), .ZN(n2680) );
  AOI22_X1 U3749 ( .A1(n3181), .A2(rC4[42]), .B1(n3041), .B2(rC4[41]), .ZN(
        n2661) );
  OAI22_X1 U3750 ( .A1(rC7[61]), .A2(n3038), .B1(rC7[60]), .B2(n3128), .ZN(
        n2548) );
  NOR3_X1 U3751 ( .A1(n2793), .A2(rC3[10]), .A3(n3151), .ZN(n2790) );
  AOI22_X1 U3752 ( .A1(n3090), .A2(rC2[9]), .B1(n2266), .B2(rC2[8]), .ZN(n2702) );
  AOI22_X1 U3753 ( .A1(n3062), .A2(rC6[39]), .B1(n3037), .B2(rC6[38]), .ZN(
        n2583) );
  NOR3_X1 U3754 ( .A1(n3053), .A2(rC7[62]), .A3(n2551), .ZN(n2550) );
  OAI22_X1 U3755 ( .A1(rC6[56]), .A2(n3215), .B1(rC6[55]), .B2(n3133), .ZN(
        n2553) );
  INV_X1 U3756 ( .A(n2557), .ZN(n2413) );
  OAI211_X1 U3757 ( .C1(rC3[37]), .C2(n3245), .A(n2766), .B(n2813), .ZN(n2760)
         );
  AOI211_X1 U3758 ( .C1(rC1[36]), .C2(n3075), .A(n2814), .B(n2815), .ZN(n2813)
         );
  AOI211_X1 U3759 ( .C1(rC3[36]), .C2(n3178), .A(n3149), .B(rC3[35]), .ZN(
        n2814) );
  NOR3_X1 U3760 ( .A1(n3049), .A2(rC3[34]), .A3(n2816), .ZN(n2815) );
  OAI22_X1 U3761 ( .A1(n2668), .A2(n2669), .B1(n2670), .B2(n2671), .ZN(n2667)
         );
  AOI22_X1 U3762 ( .A1(rC4[37]), .A2(n3106), .B1(rC4[38]), .B2(n3032), .ZN(
        n2668) );
  AOI22_X1 U3763 ( .A1(rC4[31]), .A2(n3180), .B1(rC4[32]), .B2(n3086), .ZN(
        n2670) );
  OAI22_X1 U3764 ( .A1(rC1[2]), .A2(n2337), .B1(rC1[1]), .B2(n3157), .ZN(n2803) );
  OAI211_X1 U3765 ( .C1(rC7[25]), .C2(n3071), .A(n2449), .B(n2628), .ZN(n2591)
         );
  INV_X1 U3766 ( .A(n2589), .ZN(n2449) );
  OAI211_X1 U3767 ( .C1(rC3[25]), .C2(n3079), .A(n2807), .B(n2808), .ZN(n2773)
         );
  AOI211_X1 U3768 ( .C1(rC1[24]), .C2(n3076), .A(n2809), .B(n2810), .ZN(n2808)
         );
  AOI211_X1 U3769 ( .C1(rC3[24]), .C2(n3189), .A(n3150), .B(rC3[23]), .ZN(
        n2809) );
  NOR3_X1 U3770 ( .A1(n3014), .A2(rC3[22]), .A3(n2811), .ZN(n2810) );
  NOR2_X1 U3771 ( .A1(n3116), .A2(rC6[63]), .ZN(n2551) );
  AOI22_X1 U3772 ( .A1(rC6[28]), .A2(n3018), .B1(rC6[29]), .B2(n3119), .ZN(
        n2632) );
  AOI22_X1 U3773 ( .A1(rC1[28]), .A2(n3029), .B1(rC1[29]), .B2(n3144), .ZN(
        n2812) );
  AOI22_X1 U3774 ( .A1(rC1[52]), .A2(n3030), .B1(rC1[53]), .B2(n3145), .ZN(
        n2748) );
  AOI22_X1 U3775 ( .A1(rC2[52]), .A2(n3031), .B1(rC2[53]), .B2(n3146), .ZN(
        n2652) );
  AOI22_X1 U3776 ( .A1(rC1[4]), .A2(n3107), .B1(rC1[5]), .B2(n3033), .ZN(n2800) );
  OAI21_X1 U3777 ( .B1(rC1[11]), .B2(n3091), .A(n2799), .ZN(n2793) );
  AOI22_X1 U3778 ( .A1(n2711), .A2(n2712), .B1(rC2[6]), .B2(n3201), .ZN(n2710)
         );
  OAI21_X1 U3779 ( .B1(rC2[4]), .B2(n3236), .A(n2711), .ZN(n2709) );
  NAND4_X1 U3780 ( .A1(n2827), .A2(n2828), .A3(n2740), .A4(n2829), .ZN(n2738)
         );
  OAI211_X1 U3781 ( .C1(rC1[60]), .C2(n3011), .A(n3083), .B(rC1[59]), .ZN(
        n2828) );
  AOI221_X1 U3782 ( .B1(rC1[61]), .B2(n3141), .C1(rC1[60]), .C2(n3011), .A(
        n2830), .ZN(n2829) );
  NOR3_X1 U3783 ( .A1(n3051), .A2(rC3[58]), .A3(n2831), .ZN(n2830) );
  INV_X1 U3784 ( .A(n2636), .ZN(n2436) );
  AOI21_X1 U3785 ( .B1(n3060), .B2(rC7[35]), .A(n2635), .ZN(n2636) );
  INV_X1 U3786 ( .A(n2825), .ZN(n2136) );
  AOI21_X1 U3787 ( .B1(n3065), .B2(rC1[50]), .A(n2817), .ZN(n2825) );
  AOI22_X1 U3788 ( .A1(rC7[49]), .A2(n3173), .B1(rC7[50]), .B2(n3027), .ZN(
        n2560) );
  AOI221_X1 U3789 ( .B1(n2547), .B2(n2548), .C1(n2405), .C2(n2549), .A(n2550), 
        .ZN(n2546) );
  OAI211_X1 U3790 ( .C1(rC2[18]), .C2(n3012), .A(n3085), .B(rC2[17]), .ZN(
        n2716) );
  AOI22_X1 U3791 ( .A1(rC4[1]), .A2(n3480), .B1(n3487), .B2(n3381), .ZN(n2713)
         );
  AOI22_X1 U3792 ( .A1(rC2[20]), .A2(n3111), .B1(rC2[21]), .B2(n3034), .ZN(
        n2676) );
  NOR2_X1 U3793 ( .A1(n3102), .A2(rC1[48]), .ZN(n2824) );
  NOR2_X1 U3794 ( .A1(n3056), .A2(rC3[51]), .ZN(n2817) );
  NOR2_X1 U3795 ( .A1(n3055), .A2(rC6[36]), .ZN(n2635) );
  NOR2_X1 U3796 ( .A1(n3057), .A2(rC4[51]), .ZN(n2658) );
  NOR2_X1 U3797 ( .A1(n3103), .A2(rC2[48]), .ZN(n2729) );
  NOR2_X1 U3798 ( .A1(n3059), .A2(rC2[24]), .ZN(n2686) );
  NOR2_X1 U3799 ( .A1(n3176), .A2(rC4[27]), .ZN(n2679) );
  OAI221_X1 U3800 ( .B1(rC6[27]), .B2(n3249), .C1(rC6[28]), .C2(n3018), .A(
        n2587), .ZN(n2586) );
  AOI22_X1 U3801 ( .A1(rC7[25]), .A2(n3071), .B1(rC7[26]), .B2(n3025), .ZN(
        n2588) );
  OAI221_X1 U3802 ( .B1(rC1[27]), .B2(n3007), .C1(rC1[28]), .C2(n3029), .A(
        n2770), .ZN(n2769) );
  AOI22_X1 U3803 ( .A1(rC3[25]), .A2(n3079), .B1(rC3[26]), .B2(n3235), .ZN(
        n2771) );
  OAI21_X1 U3804 ( .B1(rC1[52]), .B2(n3030), .A(n2749), .ZN(n2820) );
  OAI21_X1 U3805 ( .B1(rC2[52]), .B2(n3031), .A(n2653), .ZN(n2725) );
  AOI211_X1 U3806 ( .C1(n3020), .C2(rC2[49]), .A(n2214), .B(n2727), .ZN(n2723)
         );
  OAI21_X1 U3807 ( .B1(n3188), .B2(rC4[48]), .A(n2217), .ZN(n2727) );
  INV_X1 U3808 ( .A(n2728), .ZN(n2217) );
  NAND4_X1 U3809 ( .A1(n2732), .A2(n2733), .A3(n2644), .A4(n2734), .ZN(n2642)
         );
  OAI211_X1 U3810 ( .C1(rC2[60]), .C2(n3010), .A(n3082), .B(rC2[59]), .ZN(
        n2733) );
  AOI221_X1 U3811 ( .B1(rC2[61]), .B2(n3140), .C1(rC2[60]), .C2(n3010), .A(
        n2735), .ZN(n2734) );
  NOR3_X1 U3812 ( .A1(n3050), .A2(rC4[58]), .A3(n2736), .ZN(n2735) );
  AOI211_X1 U3813 ( .C1(rC2[18]), .C2(n3012), .A(n2688), .B(n2689), .ZN(n2687)
         );
  OAI21_X1 U3814 ( .B1(rC4[19]), .B2(n3094), .A(n2716), .ZN(n2688) );
  AOI22_X1 U3815 ( .A1(rC6[20]), .A2(n3092), .B1(rC6[21]), .B2(n3194), .ZN(
        n2594) );
  INV_X1 U3816 ( .A(n2591), .ZN(n2448) );
  OAI21_X1 U3817 ( .B1(rC1[62]), .B2(n3080), .A(n2826), .ZN(n2741) );
  INV_X1 U3818 ( .A(rC3[63]), .ZN(n2276) );
  INV_X1 U3819 ( .A(rC4[8]), .ZN(n2266) );
  AOI211_X1 U3820 ( .C1(n3019), .C2(rC1[49]), .A(n2136), .B(n2822), .ZN(n2818)
         );
  OAI21_X1 U3821 ( .B1(n3187), .B2(rC3[48]), .A(n2140), .ZN(n2822) );
  INV_X1 U3822 ( .A(n2823), .ZN(n2140) );
  OAI21_X1 U3823 ( .B1(rC6[46]), .B2(n3212), .A(n2566), .ZN(n2564) );
  INV_X1 U3824 ( .A(rC1[12]), .ZN(n2183) );
  INV_X1 U3825 ( .A(rC3[2]), .ZN(n2337) );
  AOI22_X1 U3826 ( .A1(rC1[20]), .A2(n3093), .B1(rC1[21]), .B2(n3202), .ZN(
        n2776) );
  INV_X1 U3827 ( .A(n2773), .ZN(n2167) );
  AOI22_X1 U3828 ( .A1(n2599), .A2(n2600), .B1(rC6[18]), .B2(n3193), .ZN(n2598) );
  OAI221_X1 U3829 ( .B1(rC6[15]), .B2(n3008), .C1(rC6[16]), .C2(n3217), .A(
        n2599), .ZN(n2597) );
  AOI22_X1 U3830 ( .A1(n2702), .A2(n2703), .B1(rC4[10]), .B2(n3142), .ZN(n2701) );
  OAI22_X1 U3831 ( .A1(rC2[8]), .A2(n2266), .B1(rC2[7]), .B2(n3169), .ZN(n2703) );
  NAND2_X1 U3832 ( .A1(rC1[63]), .A2(n2276), .ZN(n2740) );
  NAND2_X1 U3833 ( .A1(rC1[62]), .A2(n3080), .ZN(n2827) );
  NAND2_X1 U3834 ( .A1(rC3[12]), .A2(n3417), .ZN(n2799) );
  NAND2_X1 U3835 ( .A1(rC6[13]), .A2(n3403), .ZN(n2617) );
  NAND2_X1 U3836 ( .A1(rC2[62]), .A2(n3081), .ZN(n2732) );
  INV_X1 U3837 ( .A(n2638), .ZN(n2405) );
  OAI221_X1 U3838 ( .B1(rC6[59]), .B2(n3147), .C1(rC6[60]), .C2(n3218), .A(
        n2547), .ZN(n2638) );
  AND3_X1 U3839 ( .A1(rC2[34]), .A2(n3048), .A3(n2718), .ZN(n2721) );
  INV_X1 U3840 ( .A(n2631), .ZN(n2452) );
  AOI21_X1 U3841 ( .B1(n3061), .B2(rC7[23]), .A(n2630), .ZN(n2631) );
  INV_X1 U3842 ( .A(rC3[3]), .ZN(n2336) );
  INV_X1 U3843 ( .A(n2730), .ZN(n2214) );
  AOI21_X1 U3844 ( .B1(n3067), .B2(rC2[50]), .A(n2658), .ZN(n2730) );
  INV_X1 U3845 ( .A(rC3[12]), .ZN(n2327) );
  INV_X1 U3846 ( .A(rC4[11]), .ZN(n2263) );
  INV_X1 U3847 ( .A(n3383), .ZN(n2181) );
  INV_X1 U3848 ( .A(n3483), .ZN(n2260) );
  INV_X1 U3849 ( .A(n3385), .ZN(n2331) );
  OAI221_X1 U3850 ( .B1(mX4[2]), .B2(n2053), .C1(mX4[1]), .C2(n2054), .A(n2896), .ZN(n2895) );
  OAI211_X1 U3851 ( .C1(mX3[1]), .C2(n2118), .A(n2119), .B(mX3[0]), .ZN(n2896)
         );
  OAI221_X1 U3852 ( .B1(mX2[2]), .B2(n1924), .C1(mX2[1]), .C2(n1925), .A(n2960), .ZN(n2959) );
  OAI211_X1 U3853 ( .C1(mX1[1]), .C2(n1989), .A(n1990), .B(mX1[0]), .ZN(n2960)
         );
  OAI221_X1 U3854 ( .B1(mX4[6]), .B2(n2049), .C1(mX4[5]), .C2(n2050), .A(n2892), .ZN(n2891) );
  OAI221_X1 U3855 ( .B1(mX3[5]), .B2(n2114), .C1(mX3[4]), .C2(n2115), .A(n2893), .ZN(n2892) );
  OAI221_X1 U3856 ( .B1(mX4[4]), .B2(n2051), .C1(mX4[3]), .C2(n2052), .A(n2894), .ZN(n2893) );
  OAI221_X1 U3857 ( .B1(mX3[3]), .B2(n2116), .C1(mX3[2]), .C2(n2117), .A(n2895), .ZN(n2894) );
  OAI221_X1 U3858 ( .B1(mX2[6]), .B2(n1920), .C1(mX2[5]), .C2(n1921), .A(n2956), .ZN(n2955) );
  OAI221_X1 U3859 ( .B1(mX1[5]), .B2(n1985), .C1(mX1[4]), .C2(n1986), .A(n2957), .ZN(n2956) );
  OAI221_X1 U3860 ( .B1(mX2[4]), .B2(n1922), .C1(mX2[3]), .C2(n1923), .A(n2958), .ZN(n2957) );
  OAI221_X1 U3861 ( .B1(mX1[3]), .B2(n1987), .C1(mX1[2]), .C2(n1988), .A(n2959), .ZN(n2958) );
  OAI221_X1 U3862 ( .B1(mX4[9]), .B2(n2046), .C1(mX4[10]), .C2(n2045), .A(
        n2888), .ZN(n2887) );
  OAI221_X1 U3863 ( .B1(mX3[9]), .B2(n2110), .C1(mX3[8]), .C2(n2111), .A(n2889), .ZN(n2888) );
  OAI221_X1 U3864 ( .B1(mX4[8]), .B2(n2047), .C1(mX4[7]), .C2(n2048), .A(n2890), .ZN(n2889) );
  OAI221_X1 U3865 ( .B1(mX3[7]), .B2(n2112), .C1(mX3[6]), .C2(n2113), .A(n2891), .ZN(n2890) );
  OAI221_X1 U3866 ( .B1(mX2[9]), .B2(n1917), .C1(mX2[10]), .C2(n1916), .A(
        n2952), .ZN(n2951) );
  OAI221_X1 U3867 ( .B1(mX1[9]), .B2(n1981), .C1(mX1[8]), .C2(n1982), .A(n2953), .ZN(n2952) );
  OAI221_X1 U3868 ( .B1(mX2[8]), .B2(n1918), .C1(mX2[7]), .C2(n1919), .A(n2954), .ZN(n2953) );
  OAI221_X1 U3869 ( .B1(mX1[7]), .B2(n1983), .C1(mX1[6]), .C2(n1984), .A(n2955), .ZN(n2954) );
  OAI221_X1 U3870 ( .B1(mX4[14]), .B2(n2041), .C1(mX4[13]), .C2(n2042), .A(
        n2884), .ZN(n2883) );
  OAI221_X1 U3871 ( .B1(mX3[13]), .B2(n2106), .C1(mX3[12]), .C2(n2107), .A(
        n2885), .ZN(n2884) );
  OAI221_X1 U3872 ( .B1(mX4[12]), .B2(n2043), .C1(mX4[11]), .C2(n2044), .A(
        n2886), .ZN(n2885) );
  OAI221_X1 U3873 ( .B1(mX3[11]), .B2(n2108), .C1(mX3[10]), .C2(n2109), .A(
        n2887), .ZN(n2886) );
  OAI221_X1 U3874 ( .B1(mX2[14]), .B2(n1912), .C1(mX2[13]), .C2(n1913), .A(
        n2948), .ZN(n2947) );
  OAI221_X1 U3875 ( .B1(mX1[13]), .B2(n1977), .C1(mX1[12]), .C2(n1978), .A(
        n2949), .ZN(n2948) );
  OAI221_X1 U3876 ( .B1(mX2[12]), .B2(n1914), .C1(mX2[11]), .C2(n1915), .A(
        n2950), .ZN(n2949) );
  OAI221_X1 U3877 ( .B1(mX1[11]), .B2(n1979), .C1(mX1[10]), .C2(n1980), .A(
        n2951), .ZN(n2950) );
  OAI221_X1 U3878 ( .B1(mX4[18]), .B2(n2037), .C1(mX4[17]), .C2(n2038), .A(
        n2880), .ZN(n2879) );
  OAI221_X1 U3879 ( .B1(mX3[17]), .B2(n2102), .C1(mX3[16]), .C2(n2103), .A(
        n2881), .ZN(n2880) );
  OAI221_X1 U3880 ( .B1(mX4[16]), .B2(n2039), .C1(mX4[15]), .C2(n2040), .A(
        n2882), .ZN(n2881) );
  OAI221_X1 U3881 ( .B1(mX3[15]), .B2(n2104), .C1(mX3[14]), .C2(n2105), .A(
        n2883), .ZN(n2882) );
  OAI221_X1 U3882 ( .B1(mX2[18]), .B2(n1908), .C1(mX2[17]), .C2(n1909), .A(
        n2944), .ZN(n2943) );
  OAI221_X1 U3883 ( .B1(mX1[17]), .B2(n1973), .C1(mX1[16]), .C2(n1974), .A(
        n2945), .ZN(n2944) );
  OAI221_X1 U3884 ( .B1(mX2[16]), .B2(n1910), .C1(mX2[15]), .C2(n1911), .A(
        n2946), .ZN(n2945) );
  OAI221_X1 U3885 ( .B1(mX1[15]), .B2(n1975), .C1(mX1[14]), .C2(n1976), .A(
        n2947), .ZN(n2946) );
  OAI221_X1 U3886 ( .B1(mX4[22]), .B2(n2033), .C1(mX4[21]), .C2(n2034), .A(
        n2876), .ZN(n2875) );
  OAI221_X1 U3887 ( .B1(mX3[21]), .B2(n2098), .C1(mX3[20]), .C2(n2099), .A(
        n2877), .ZN(n2876) );
  OAI221_X1 U3888 ( .B1(mX4[20]), .B2(n2035), .C1(mX4[19]), .C2(n2036), .A(
        n2878), .ZN(n2877) );
  OAI221_X1 U3889 ( .B1(mX3[19]), .B2(n2100), .C1(mX3[18]), .C2(n2101), .A(
        n2879), .ZN(n2878) );
  OAI221_X1 U3890 ( .B1(mX2[22]), .B2(n1904), .C1(mX2[21]), .C2(n1905), .A(
        n2940), .ZN(n2939) );
  OAI221_X1 U3891 ( .B1(mX1[21]), .B2(n1969), .C1(mX1[20]), .C2(n1970), .A(
        n2941), .ZN(n2940) );
  OAI221_X1 U3892 ( .B1(mX2[20]), .B2(n1906), .C1(mX2[19]), .C2(n1907), .A(
        n2942), .ZN(n2941) );
  OAI221_X1 U3893 ( .B1(mX1[19]), .B2(n1971), .C1(mX1[18]), .C2(n1972), .A(
        n2943), .ZN(n2942) );
  OAI221_X1 U3894 ( .B1(mX4[26]), .B2(n2029), .C1(mX4[25]), .C2(n2030), .A(
        n2872), .ZN(n2871) );
  OAI221_X1 U3895 ( .B1(mX3[25]), .B2(n2094), .C1(mX3[24]), .C2(n2095), .A(
        n2873), .ZN(n2872) );
  OAI221_X1 U3896 ( .B1(mX4[24]), .B2(n2031), .C1(mX4[23]), .C2(n2032), .A(
        n2874), .ZN(n2873) );
  OAI221_X1 U3897 ( .B1(mX3[23]), .B2(n2096), .C1(mX3[22]), .C2(n2097), .A(
        n2875), .ZN(n2874) );
  OAI221_X1 U3898 ( .B1(mX2[26]), .B2(n1900), .C1(mX2[25]), .C2(n1901), .A(
        n2936), .ZN(n2935) );
  OAI221_X1 U3899 ( .B1(mX1[25]), .B2(n1965), .C1(mX1[24]), .C2(n1966), .A(
        n2937), .ZN(n2936) );
  OAI221_X1 U3900 ( .B1(mX2[24]), .B2(n1902), .C1(mX2[23]), .C2(n1903), .A(
        n2938), .ZN(n2937) );
  OAI221_X1 U3901 ( .B1(mX1[23]), .B2(n1967), .C1(mX1[22]), .C2(n1968), .A(
        n2939), .ZN(n2938) );
  OAI221_X1 U3902 ( .B1(mX4[30]), .B2(n2025), .C1(mX4[29]), .C2(n2026), .A(
        n2868), .ZN(n2867) );
  OAI221_X1 U3903 ( .B1(mX3[29]), .B2(n2090), .C1(mX3[28]), .C2(n2091), .A(
        n2869), .ZN(n2868) );
  OAI221_X1 U3904 ( .B1(mX4[28]), .B2(n2027), .C1(mX4[27]), .C2(n2028), .A(
        n2870), .ZN(n2869) );
  OAI221_X1 U3905 ( .B1(mX3[27]), .B2(n2092), .C1(mX3[26]), .C2(n2093), .A(
        n2871), .ZN(n2870) );
  OAI221_X1 U3906 ( .B1(mX2[30]), .B2(n1896), .C1(mX2[29]), .C2(n1897), .A(
        n2932), .ZN(n2931) );
  OAI221_X1 U3907 ( .B1(mX1[29]), .B2(n1961), .C1(mX1[28]), .C2(n1962), .A(
        n2933), .ZN(n2932) );
  OAI221_X1 U3908 ( .B1(mX2[28]), .B2(n1898), .C1(mX2[27]), .C2(n1899), .A(
        n2934), .ZN(n2933) );
  OAI221_X1 U3909 ( .B1(mX1[27]), .B2(n1963), .C1(mX1[26]), .C2(n1964), .A(
        n2935), .ZN(n2934) );
  OAI221_X1 U3910 ( .B1(mX4[34]), .B2(n2021), .C1(mX4[33]), .C2(n2022), .A(
        n2864), .ZN(n2863) );
  OAI221_X1 U3911 ( .B1(mX3[33]), .B2(n2086), .C1(mX3[32]), .C2(n2087), .A(
        n2865), .ZN(n2864) );
  OAI221_X1 U3912 ( .B1(mX4[32]), .B2(n2023), .C1(mX4[31]), .C2(n2024), .A(
        n2866), .ZN(n2865) );
  OAI221_X1 U3913 ( .B1(mX3[31]), .B2(n2088), .C1(mX3[30]), .C2(n2089), .A(
        n2867), .ZN(n2866) );
  OAI221_X1 U3914 ( .B1(mX2[34]), .B2(n1892), .C1(mX2[33]), .C2(n1893), .A(
        n2928), .ZN(n2927) );
  OAI221_X1 U3915 ( .B1(mX1[33]), .B2(n1957), .C1(mX1[32]), .C2(n1958), .A(
        n2929), .ZN(n2928) );
  OAI221_X1 U3916 ( .B1(mX2[32]), .B2(n1894), .C1(mX2[31]), .C2(n1895), .A(
        n2930), .ZN(n2929) );
  OAI221_X1 U3917 ( .B1(mX1[31]), .B2(n1959), .C1(mX1[30]), .C2(n1960), .A(
        n2931), .ZN(n2930) );
  OAI221_X1 U3918 ( .B1(mX4[38]), .B2(n2017), .C1(mX4[37]), .C2(n2018), .A(
        n2860), .ZN(n2859) );
  OAI221_X1 U3919 ( .B1(mX3[37]), .B2(n2082), .C1(mX3[36]), .C2(n2083), .A(
        n2861), .ZN(n2860) );
  OAI221_X1 U3920 ( .B1(mX4[36]), .B2(n2019), .C1(mX4[35]), .C2(n2020), .A(
        n2862), .ZN(n2861) );
  OAI221_X1 U3921 ( .B1(mX3[35]), .B2(n2084), .C1(mX3[34]), .C2(n2085), .A(
        n2863), .ZN(n2862) );
  OAI221_X1 U3922 ( .B1(mX2[38]), .B2(n1888), .C1(mX2[37]), .C2(n1889), .A(
        n2924), .ZN(n2923) );
  OAI221_X1 U3923 ( .B1(mX1[37]), .B2(n1953), .C1(mX1[36]), .C2(n1954), .A(
        n2925), .ZN(n2924) );
  OAI221_X1 U3924 ( .B1(mX2[36]), .B2(n1890), .C1(mX2[35]), .C2(n1891), .A(
        n2926), .ZN(n2925) );
  OAI221_X1 U3925 ( .B1(mX1[35]), .B2(n1955), .C1(mX1[34]), .C2(n1956), .A(
        n2927), .ZN(n2926) );
  OAI221_X1 U3926 ( .B1(mX4[42]), .B2(n2013), .C1(mX4[41]), .C2(n2014), .A(
        n2856), .ZN(n2855) );
  OAI221_X1 U3927 ( .B1(mX3[41]), .B2(n2078), .C1(mX3[40]), .C2(n2079), .A(
        n2857), .ZN(n2856) );
  OAI221_X1 U3928 ( .B1(mX4[40]), .B2(n2015), .C1(mX4[39]), .C2(n2016), .A(
        n2858), .ZN(n2857) );
  OAI221_X1 U3929 ( .B1(mX3[39]), .B2(n2080), .C1(mX3[38]), .C2(n2081), .A(
        n2859), .ZN(n2858) );
  OAI221_X1 U3930 ( .B1(mX2[42]), .B2(n1884), .C1(mX2[41]), .C2(n1885), .A(
        n2920), .ZN(n2919) );
  OAI221_X1 U3931 ( .B1(mX1[41]), .B2(n1949), .C1(mX1[40]), .C2(n1950), .A(
        n2921), .ZN(n2920) );
  OAI221_X1 U3932 ( .B1(mX2[40]), .B2(n1886), .C1(mX2[39]), .C2(n1887), .A(
        n2922), .ZN(n2921) );
  OAI221_X1 U3933 ( .B1(mX1[39]), .B2(n1951), .C1(mX1[38]), .C2(n1952), .A(
        n2923), .ZN(n2922) );
  OAI221_X1 U3934 ( .B1(mX4[46]), .B2(n2009), .C1(mX4[45]), .C2(n2010), .A(
        n2852), .ZN(n2851) );
  OAI221_X1 U3935 ( .B1(mX3[45]), .B2(n2074), .C1(mX3[44]), .C2(n2075), .A(
        n2853), .ZN(n2852) );
  OAI221_X1 U3936 ( .B1(mX4[44]), .B2(n2011), .C1(mX4[43]), .C2(n2012), .A(
        n2854), .ZN(n2853) );
  OAI221_X1 U3937 ( .B1(mX3[43]), .B2(n2076), .C1(mX3[42]), .C2(n2077), .A(
        n2855), .ZN(n2854) );
  OAI221_X1 U3938 ( .B1(mX2[46]), .B2(n1880), .C1(mX2[45]), .C2(n1881), .A(
        n2916), .ZN(n2915) );
  OAI221_X1 U3939 ( .B1(mX1[45]), .B2(n1945), .C1(mX1[44]), .C2(n1946), .A(
        n2917), .ZN(n2916) );
  OAI221_X1 U3940 ( .B1(mX2[44]), .B2(n1882), .C1(mX2[43]), .C2(n1883), .A(
        n2918), .ZN(n2917) );
  OAI221_X1 U3941 ( .B1(mX1[43]), .B2(n1947), .C1(mX1[42]), .C2(n1948), .A(
        n2919), .ZN(n2918) );
  OAI221_X1 U3942 ( .B1(mX4[50]), .B2(n2005), .C1(mX4[49]), .C2(n2006), .A(
        n2848), .ZN(n2847) );
  OAI221_X1 U3943 ( .B1(mX3[49]), .B2(n2070), .C1(mX3[48]), .C2(n2071), .A(
        n2849), .ZN(n2848) );
  OAI221_X1 U3944 ( .B1(mX4[48]), .B2(n2007), .C1(mX4[47]), .C2(n2008), .A(
        n2850), .ZN(n2849) );
  OAI221_X1 U3945 ( .B1(mX3[47]), .B2(n2072), .C1(mX3[46]), .C2(n2073), .A(
        n2851), .ZN(n2850) );
  OAI221_X1 U3946 ( .B1(mX2[50]), .B2(n1876), .C1(mX2[49]), .C2(n1877), .A(
        n2912), .ZN(n2911) );
  OAI221_X1 U3947 ( .B1(mX1[49]), .B2(n1941), .C1(mX1[48]), .C2(n1942), .A(
        n2913), .ZN(n2912) );
  OAI221_X1 U3948 ( .B1(mX2[48]), .B2(n1878), .C1(mX2[47]), .C2(n1879), .A(
        n2914), .ZN(n2913) );
  OAI221_X1 U3949 ( .B1(mX1[47]), .B2(n1943), .C1(mX1[46]), .C2(n1944), .A(
        n2915), .ZN(n2914) );
  OAI221_X1 U3950 ( .B1(mX4[54]), .B2(n2001), .C1(mX4[53]), .C2(n2002), .A(
        n2844), .ZN(n2843) );
  OAI221_X1 U3951 ( .B1(mX3[53]), .B2(n2066), .C1(mX3[52]), .C2(n2067), .A(
        n2845), .ZN(n2844) );
  OAI221_X1 U3952 ( .B1(mX4[52]), .B2(n2003), .C1(mX4[51]), .C2(n2004), .A(
        n2846), .ZN(n2845) );
  OAI221_X1 U3953 ( .B1(mX3[51]), .B2(n2068), .C1(mX3[50]), .C2(n2069), .A(
        n2847), .ZN(n2846) );
  OAI221_X1 U3954 ( .B1(mX2[54]), .B2(n1872), .C1(mX2[53]), .C2(n1873), .A(
        n2908), .ZN(n2907) );
  OAI221_X1 U3955 ( .B1(mX1[53]), .B2(n1937), .C1(mX1[52]), .C2(n1938), .A(
        n2909), .ZN(n2908) );
  OAI221_X1 U3956 ( .B1(mX2[52]), .B2(n1874), .C1(mX2[51]), .C2(n1875), .A(
        n2910), .ZN(n2909) );
  OAI221_X1 U3957 ( .B1(mX1[51]), .B2(n1939), .C1(mX1[50]), .C2(n1940), .A(
        n2911), .ZN(n2910) );
  OAI221_X1 U3958 ( .B1(mX4[58]), .B2(n1997), .C1(mX4[57]), .C2(n1998), .A(
        n2840), .ZN(n2839) );
  OAI221_X1 U3959 ( .B1(mX3[57]), .B2(n2062), .C1(mX3[56]), .C2(n2063), .A(
        n2841), .ZN(n2840) );
  OAI221_X1 U3960 ( .B1(mX4[56]), .B2(n1999), .C1(mX4[55]), .C2(n2000), .A(
        n2842), .ZN(n2841) );
  OAI221_X1 U3961 ( .B1(mX3[55]), .B2(n2064), .C1(mX3[54]), .C2(n2065), .A(
        n2843), .ZN(n2842) );
  OAI221_X1 U3962 ( .B1(mX2[58]), .B2(n1868), .C1(mX2[57]), .C2(n1869), .A(
        n2904), .ZN(n2903) );
  OAI221_X1 U3963 ( .B1(mX1[57]), .B2(n1933), .C1(mX1[56]), .C2(n1934), .A(
        n2905), .ZN(n2904) );
  OAI221_X1 U3964 ( .B1(mX2[56]), .B2(n1870), .C1(mX2[55]), .C2(n1871), .A(
        n2906), .ZN(n2905) );
  OAI221_X1 U3965 ( .B1(mX1[55]), .B2(n1935), .C1(mX1[54]), .C2(n1936), .A(
        n2907), .ZN(n2906) );
  OAI21_X1 U3966 ( .B1(mX4[61]), .B2(n1994), .A(n2836), .ZN(n2835) );
  OAI221_X1 U3967 ( .B1(mX3[61]), .B2(n2058), .C1(mX3[60]), .C2(n2059), .A(
        n2837), .ZN(n2836) );
  OAI221_X1 U3968 ( .B1(mX4[60]), .B2(n1995), .C1(mX4[59]), .C2(n1996), .A(
        n2838), .ZN(n2837) );
  OAI221_X1 U3969 ( .B1(mX3[59]), .B2(n2060), .C1(mX3[58]), .C2(n2061), .A(
        n2839), .ZN(n2838) );
  OAI21_X1 U3970 ( .B1(mX2[61]), .B2(n1865), .A(n2900), .ZN(n2899) );
  OAI221_X1 U3971 ( .B1(mX1[61]), .B2(n1929), .C1(mX1[60]), .C2(n1930), .A(
        n2901), .ZN(n2900) );
  OAI221_X1 U3972 ( .B1(mX2[60]), .B2(n1866), .C1(mX2[59]), .C2(n1867), .A(
        n2902), .ZN(n2901) );
  OAI221_X1 U3973 ( .B1(mX1[59]), .B2(n1931), .C1(mX1[58]), .C2(n1932), .A(
        n2903), .ZN(n2902) );
  INV_X1 U3974 ( .A(mX3[63]), .ZN(n1992) );
  INV_X1 U3975 ( .A(mX1[63]), .ZN(n1863) );
  INV_X1 U3976 ( .A(mX4[0]), .ZN(n2119) );
  INV_X1 U3977 ( .A(mX2[0]), .ZN(n1990) );
  INV_X1 U3978 ( .A(mX3[61]), .ZN(n1994) );
  INV_X1 U3979 ( .A(mX1[61]), .ZN(n1865) );
  INV_X1 U3980 ( .A(mX4[62]), .ZN(n2057) );
  INV_X1 U3981 ( .A(mX2[62]), .ZN(n1928) );
  INV_X1 U3982 ( .A(mX3[1]), .ZN(n2054) );
  INV_X1 U3983 ( .A(mX1[1]), .ZN(n1925) );
  INV_X1 U3984 ( .A(mX4[2]), .ZN(n2117) );
  INV_X1 U3985 ( .A(mX2[2]), .ZN(n1988) );
  INV_X1 U3986 ( .A(mX3[3]), .ZN(n2052) );
  INV_X1 U3987 ( .A(mX1[3]), .ZN(n1923) );
  INV_X1 U3988 ( .A(mX4[4]), .ZN(n2115) );
  INV_X1 U3989 ( .A(mX2[4]), .ZN(n1986) );
  INV_X1 U3990 ( .A(mX3[5]), .ZN(n2050) );
  INV_X1 U3991 ( .A(mX1[5]), .ZN(n1921) );
  INV_X1 U3992 ( .A(mX4[6]), .ZN(n2113) );
  INV_X1 U3993 ( .A(mX2[6]), .ZN(n1984) );
  INV_X1 U3994 ( .A(mX3[7]), .ZN(n2048) );
  INV_X1 U3995 ( .A(mX1[7]), .ZN(n1919) );
  INV_X1 U3996 ( .A(mX4[8]), .ZN(n2111) );
  INV_X1 U3997 ( .A(mX2[8]), .ZN(n1982) );
  INV_X1 U3998 ( .A(mX3[10]), .ZN(n2045) );
  INV_X1 U3999 ( .A(mX1[10]), .ZN(n1916) );
  INV_X1 U4000 ( .A(mX4[10]), .ZN(n2109) );
  INV_X1 U4001 ( .A(mX2[10]), .ZN(n1980) );
  INV_X1 U4002 ( .A(mX3[11]), .ZN(n2044) );
  INV_X1 U4003 ( .A(mX1[11]), .ZN(n1915) );
  INV_X1 U4004 ( .A(mX4[12]), .ZN(n2107) );
  INV_X1 U4005 ( .A(mX2[12]), .ZN(n1978) );
  INV_X1 U4006 ( .A(mX3[13]), .ZN(n2042) );
  INV_X1 U4007 ( .A(mX1[13]), .ZN(n1913) );
  INV_X1 U4008 ( .A(mX4[14]), .ZN(n2105) );
  INV_X1 U4009 ( .A(mX2[14]), .ZN(n1976) );
  INV_X1 U4010 ( .A(mX3[15]), .ZN(n2040) );
  INV_X1 U4011 ( .A(mX1[15]), .ZN(n1911) );
  INV_X1 U4012 ( .A(mX4[16]), .ZN(n2103) );
  INV_X1 U4013 ( .A(mX2[16]), .ZN(n1974) );
  INV_X1 U4014 ( .A(mX3[17]), .ZN(n2038) );
  INV_X1 U4015 ( .A(mX1[17]), .ZN(n1909) );
  INV_X1 U4016 ( .A(mX4[18]), .ZN(n2101) );
  INV_X1 U4017 ( .A(mX2[18]), .ZN(n1972) );
  INV_X1 U4018 ( .A(mX3[19]), .ZN(n2036) );
  INV_X1 U4019 ( .A(mX1[19]), .ZN(n1907) );
  INV_X1 U4020 ( .A(mX4[20]), .ZN(n2099) );
  INV_X1 U4021 ( .A(mX2[20]), .ZN(n1970) );
  INV_X1 U4022 ( .A(mX3[21]), .ZN(n2034) );
  INV_X1 U4023 ( .A(mX1[21]), .ZN(n1905) );
  INV_X1 U4024 ( .A(mX4[22]), .ZN(n2097) );
  INV_X1 U4025 ( .A(mX2[22]), .ZN(n1968) );
  INV_X1 U4026 ( .A(mX3[23]), .ZN(n2032) );
  INV_X1 U4027 ( .A(mX1[23]), .ZN(n1903) );
  INV_X1 U4028 ( .A(mX4[24]), .ZN(n2095) );
  INV_X1 U4029 ( .A(mX2[24]), .ZN(n1966) );
  INV_X1 U4030 ( .A(mX3[25]), .ZN(n2030) );
  INV_X1 U4031 ( .A(mX1[25]), .ZN(n1901) );
  INV_X1 U4032 ( .A(mX4[26]), .ZN(n2093) );
  INV_X1 U4033 ( .A(mX2[26]), .ZN(n1964) );
  INV_X1 U4034 ( .A(mX3[27]), .ZN(n2028) );
  INV_X1 U4035 ( .A(mX1[27]), .ZN(n1899) );
  INV_X1 U4036 ( .A(mX4[28]), .ZN(n2091) );
  INV_X1 U4037 ( .A(mX2[28]), .ZN(n1962) );
  INV_X1 U4038 ( .A(mX3[29]), .ZN(n2026) );
  INV_X1 U4039 ( .A(mX1[29]), .ZN(n1897) );
  INV_X1 U4040 ( .A(mX4[30]), .ZN(n2089) );
  INV_X1 U4041 ( .A(mX2[30]), .ZN(n1960) );
  INV_X1 U4042 ( .A(mX3[31]), .ZN(n2024) );
  INV_X1 U4043 ( .A(mX1[31]), .ZN(n1895) );
  INV_X1 U4044 ( .A(mX4[32]), .ZN(n2087) );
  INV_X1 U4045 ( .A(mX2[32]), .ZN(n1958) );
  INV_X1 U4046 ( .A(mX3[33]), .ZN(n2022) );
  INV_X1 U4047 ( .A(mX1[33]), .ZN(n1893) );
  INV_X1 U4048 ( .A(mX4[34]), .ZN(n2085) );
  INV_X1 U4049 ( .A(mX2[34]), .ZN(n1956) );
  INV_X1 U4050 ( .A(mX3[35]), .ZN(n2020) );
  INV_X1 U4051 ( .A(mX1[35]), .ZN(n1891) );
  INV_X1 U4052 ( .A(mX4[36]), .ZN(n2083) );
  INV_X1 U4053 ( .A(mX2[36]), .ZN(n1954) );
  INV_X1 U4054 ( .A(mX3[37]), .ZN(n2018) );
  INV_X1 U4055 ( .A(mX1[37]), .ZN(n1889) );
  INV_X1 U4056 ( .A(mX4[38]), .ZN(n2081) );
  INV_X1 U4057 ( .A(mX2[38]), .ZN(n1952) );
  INV_X1 U4058 ( .A(mX3[39]), .ZN(n2016) );
  INV_X1 U4059 ( .A(mX1[39]), .ZN(n1887) );
  INV_X1 U4060 ( .A(mX4[40]), .ZN(n2079) );
  INV_X1 U4061 ( .A(mX2[40]), .ZN(n1950) );
  INV_X1 U4062 ( .A(mX3[41]), .ZN(n2014) );
  INV_X1 U4063 ( .A(mX1[41]), .ZN(n1885) );
  INV_X1 U4064 ( .A(mX4[42]), .ZN(n2077) );
  INV_X1 U4065 ( .A(mX2[42]), .ZN(n1948) );
  INV_X1 U4066 ( .A(mX3[43]), .ZN(n2012) );
  INV_X1 U4067 ( .A(mX1[43]), .ZN(n1883) );
  INV_X1 U4068 ( .A(mX4[44]), .ZN(n2075) );
  INV_X1 U4069 ( .A(mX2[44]), .ZN(n1946) );
  INV_X1 U4070 ( .A(mX3[45]), .ZN(n2010) );
  INV_X1 U4071 ( .A(mX1[45]), .ZN(n1881) );
  INV_X1 U4072 ( .A(mX4[46]), .ZN(n2073) );
  INV_X1 U4073 ( .A(mX2[46]), .ZN(n1944) );
  INV_X1 U4074 ( .A(mX3[47]), .ZN(n2008) );
  INV_X1 U4075 ( .A(mX1[47]), .ZN(n1879) );
  INV_X1 U4076 ( .A(mX4[48]), .ZN(n2071) );
  INV_X1 U4077 ( .A(mX2[48]), .ZN(n1942) );
  INV_X1 U4078 ( .A(mX3[49]), .ZN(n2006) );
  INV_X1 U4079 ( .A(mX1[49]), .ZN(n1877) );
  INV_X1 U4080 ( .A(mX4[50]), .ZN(n2069) );
  INV_X1 U4081 ( .A(mX2[50]), .ZN(n1940) );
  INV_X1 U4082 ( .A(mX3[51]), .ZN(n2004) );
  INV_X1 U4083 ( .A(mX1[51]), .ZN(n1875) );
  INV_X1 U4084 ( .A(mX4[52]), .ZN(n2067) );
  INV_X1 U4085 ( .A(mX2[52]), .ZN(n1938) );
  INV_X1 U4086 ( .A(mX3[53]), .ZN(n2002) );
  INV_X1 U4087 ( .A(mX1[53]), .ZN(n1873) );
  INV_X1 U4088 ( .A(mX4[54]), .ZN(n2065) );
  INV_X1 U4089 ( .A(mX2[54]), .ZN(n1936) );
  INV_X1 U4090 ( .A(mX3[55]), .ZN(n2000) );
  INV_X1 U4091 ( .A(mX1[55]), .ZN(n1871) );
  INV_X1 U4092 ( .A(mX4[56]), .ZN(n2063) );
  INV_X1 U4093 ( .A(mX2[56]), .ZN(n1934) );
  INV_X1 U4094 ( .A(mX3[57]), .ZN(n1998) );
  INV_X1 U4095 ( .A(mX1[57]), .ZN(n1869) );
  INV_X1 U4096 ( .A(mX4[58]), .ZN(n2061) );
  INV_X1 U4097 ( .A(mX2[58]), .ZN(n1932) );
  INV_X1 U4098 ( .A(mX3[59]), .ZN(n1996) );
  INV_X1 U4099 ( .A(mX1[59]), .ZN(n1867) );
  INV_X1 U4100 ( .A(mX4[60]), .ZN(n2059) );
  INV_X1 U4101 ( .A(mX2[60]), .ZN(n1930) );
  INV_X1 U4102 ( .A(mX4[1]), .ZN(n2118) );
  INV_X1 U4103 ( .A(mX2[1]), .ZN(n1989) );
  INV_X1 U4104 ( .A(mX3[2]), .ZN(n2053) );
  INV_X1 U4105 ( .A(mX1[2]), .ZN(n1924) );
  INV_X1 U4106 ( .A(mX4[3]), .ZN(n2116) );
  INV_X1 U4107 ( .A(mX2[3]), .ZN(n1987) );
  INV_X1 U4108 ( .A(mX3[4]), .ZN(n2051) );
  INV_X1 U4109 ( .A(mX1[4]), .ZN(n1922) );
  INV_X1 U4110 ( .A(mX4[5]), .ZN(n2114) );
  INV_X1 U4111 ( .A(mX2[5]), .ZN(n1985) );
  INV_X1 U4112 ( .A(mX3[6]), .ZN(n2049) );
  INV_X1 U4113 ( .A(mX1[6]), .ZN(n1920) );
  INV_X1 U4114 ( .A(mX4[7]), .ZN(n2112) );
  INV_X1 U4115 ( .A(mX2[7]), .ZN(n1983) );
  INV_X1 U4116 ( .A(mX3[8]), .ZN(n2047) );
  INV_X1 U4117 ( .A(mX1[8]), .ZN(n1918) );
  INV_X1 U4118 ( .A(mX4[9]), .ZN(n2110) );
  INV_X1 U4119 ( .A(mX2[9]), .ZN(n1981) );
  INV_X1 U4120 ( .A(mX3[9]), .ZN(n2046) );
  INV_X1 U4121 ( .A(mX1[9]), .ZN(n1917) );
  INV_X1 U4122 ( .A(mX4[11]), .ZN(n2108) );
  INV_X1 U4123 ( .A(mX2[11]), .ZN(n1979) );
  INV_X1 U4124 ( .A(mX3[12]), .ZN(n2043) );
  INV_X1 U4125 ( .A(mX1[12]), .ZN(n1914) );
  INV_X1 U4126 ( .A(mX4[13]), .ZN(n2106) );
  INV_X1 U4127 ( .A(mX2[13]), .ZN(n1977) );
  INV_X1 U4128 ( .A(mX3[14]), .ZN(n2041) );
  INV_X1 U4129 ( .A(mX1[14]), .ZN(n1912) );
  INV_X1 U4130 ( .A(mX4[15]), .ZN(n2104) );
  INV_X1 U4131 ( .A(mX2[15]), .ZN(n1975) );
  INV_X1 U4132 ( .A(mX3[16]), .ZN(n2039) );
  INV_X1 U4133 ( .A(mX1[16]), .ZN(n1910) );
  INV_X1 U4134 ( .A(mX4[17]), .ZN(n2102) );
  INV_X1 U4135 ( .A(mX2[17]), .ZN(n1973) );
  INV_X1 U4136 ( .A(mX3[18]), .ZN(n2037) );
  INV_X1 U4137 ( .A(mX1[18]), .ZN(n1908) );
  INV_X1 U4138 ( .A(mX4[19]), .ZN(n2100) );
  INV_X1 U4139 ( .A(mX2[19]), .ZN(n1971) );
  INV_X1 U4140 ( .A(mX3[20]), .ZN(n2035) );
  INV_X1 U4141 ( .A(mX1[20]), .ZN(n1906) );
  INV_X1 U4142 ( .A(mX4[21]), .ZN(n2098) );
  INV_X1 U4143 ( .A(mX2[21]), .ZN(n1969) );
  INV_X1 U4144 ( .A(mX3[22]), .ZN(n2033) );
  INV_X1 U4145 ( .A(mX1[22]), .ZN(n1904) );
  INV_X1 U4146 ( .A(mX4[23]), .ZN(n2096) );
  INV_X1 U4147 ( .A(mX2[23]), .ZN(n1967) );
  INV_X1 U4148 ( .A(mX3[24]), .ZN(n2031) );
  INV_X1 U4149 ( .A(mX1[24]), .ZN(n1902) );
  INV_X1 U4150 ( .A(mX4[25]), .ZN(n2094) );
  INV_X1 U4151 ( .A(mX2[25]), .ZN(n1965) );
  INV_X1 U4152 ( .A(mX3[26]), .ZN(n2029) );
  INV_X1 U4153 ( .A(mX1[26]), .ZN(n1900) );
  INV_X1 U4154 ( .A(mX4[27]), .ZN(n2092) );
  INV_X1 U4155 ( .A(mX2[27]), .ZN(n1963) );
  INV_X1 U4156 ( .A(mX3[28]), .ZN(n2027) );
  INV_X1 U4157 ( .A(mX1[28]), .ZN(n1898) );
  INV_X1 U4158 ( .A(mX4[29]), .ZN(n2090) );
  INV_X1 U4159 ( .A(mX2[29]), .ZN(n1961) );
  INV_X1 U4160 ( .A(mX3[30]), .ZN(n2025) );
  INV_X1 U4161 ( .A(mX1[30]), .ZN(n1896) );
  INV_X1 U4162 ( .A(mX4[31]), .ZN(n2088) );
  INV_X1 U4163 ( .A(mX2[31]), .ZN(n1959) );
  INV_X1 U4164 ( .A(mX3[32]), .ZN(n2023) );
  INV_X1 U4165 ( .A(mX1[32]), .ZN(n1894) );
  INV_X1 U4166 ( .A(mX4[33]), .ZN(n2086) );
  INV_X1 U4167 ( .A(mX2[33]), .ZN(n1957) );
  INV_X1 U4168 ( .A(mX3[34]), .ZN(n2021) );
  INV_X1 U4169 ( .A(mX1[34]), .ZN(n1892) );
  INV_X1 U4170 ( .A(mX4[35]), .ZN(n2084) );
  INV_X1 U4171 ( .A(mX2[35]), .ZN(n1955) );
  INV_X1 U4172 ( .A(mX3[36]), .ZN(n2019) );
  INV_X1 U4173 ( .A(mX1[36]), .ZN(n1890) );
  INV_X1 U4174 ( .A(mX4[37]), .ZN(n2082) );
  INV_X1 U4175 ( .A(mX2[37]), .ZN(n1953) );
  INV_X1 U4176 ( .A(mX3[38]), .ZN(n2017) );
  INV_X1 U4177 ( .A(mX1[38]), .ZN(n1888) );
  INV_X1 U4178 ( .A(mX4[39]), .ZN(n2080) );
  INV_X1 U4179 ( .A(mX2[39]), .ZN(n1951) );
  INV_X1 U4180 ( .A(mX3[40]), .ZN(n2015) );
  INV_X1 U4181 ( .A(mX1[40]), .ZN(n1886) );
  INV_X1 U4182 ( .A(mX4[41]), .ZN(n2078) );
  INV_X1 U4183 ( .A(mX2[41]), .ZN(n1949) );
  INV_X1 U4184 ( .A(mX3[42]), .ZN(n2013) );
  INV_X1 U4185 ( .A(mX1[42]), .ZN(n1884) );
  INV_X1 U4186 ( .A(mX4[43]), .ZN(n2076) );
  INV_X1 U4187 ( .A(mX2[43]), .ZN(n1947) );
  INV_X1 U4188 ( .A(mX3[44]), .ZN(n2011) );
  INV_X1 U4189 ( .A(mX1[44]), .ZN(n1882) );
  INV_X1 U4190 ( .A(mX4[45]), .ZN(n2074) );
  INV_X1 U4191 ( .A(mX2[45]), .ZN(n1945) );
  INV_X1 U4192 ( .A(mX3[46]), .ZN(n2009) );
  INV_X1 U4193 ( .A(mX1[46]), .ZN(n1880) );
  INV_X1 U4194 ( .A(mX4[47]), .ZN(n2072) );
  INV_X1 U4195 ( .A(mX2[47]), .ZN(n1943) );
  INV_X1 U4196 ( .A(mX3[48]), .ZN(n2007) );
  INV_X1 U4197 ( .A(mX1[48]), .ZN(n1878) );
  INV_X1 U4198 ( .A(mX4[49]), .ZN(n2070) );
  INV_X1 U4199 ( .A(mX2[49]), .ZN(n1941) );
  INV_X1 U4200 ( .A(mX3[50]), .ZN(n2005) );
  INV_X1 U4201 ( .A(mX1[50]), .ZN(n1876) );
  INV_X1 U4202 ( .A(mX4[51]), .ZN(n2068) );
  INV_X1 U4203 ( .A(mX2[51]), .ZN(n1939) );
  INV_X1 U4204 ( .A(mX3[52]), .ZN(n2003) );
  INV_X1 U4205 ( .A(mX1[52]), .ZN(n1874) );
  INV_X1 U4206 ( .A(mX4[53]), .ZN(n2066) );
  INV_X1 U4207 ( .A(mX2[53]), .ZN(n1937) );
  INV_X1 U4208 ( .A(mX3[54]), .ZN(n2001) );
  INV_X1 U4209 ( .A(mX1[54]), .ZN(n1872) );
  INV_X1 U4210 ( .A(mX4[55]), .ZN(n2064) );
  INV_X1 U4211 ( .A(mX2[55]), .ZN(n1935) );
  INV_X1 U4212 ( .A(mX3[56]), .ZN(n1999) );
  INV_X1 U4213 ( .A(mX1[56]), .ZN(n1870) );
  INV_X1 U4214 ( .A(mX4[57]), .ZN(n2062) );
  INV_X1 U4215 ( .A(mX2[57]), .ZN(n1933) );
  INV_X1 U4216 ( .A(mX3[58]), .ZN(n1997) );
  INV_X1 U4217 ( .A(mX1[58]), .ZN(n1868) );
  INV_X1 U4218 ( .A(mX4[59]), .ZN(n2060) );
  INV_X1 U4219 ( .A(mX2[59]), .ZN(n1931) );
  INV_X1 U4220 ( .A(mX3[60]), .ZN(n1995) );
  INV_X1 U4221 ( .A(mX1[60]), .ZN(n1866) );
  INV_X1 U4222 ( .A(mX4[61]), .ZN(n2058) );
  INV_X1 U4223 ( .A(mX2[61]), .ZN(n1929) );
  INV_X1 U4224 ( .A(mX3[62]), .ZN(n1993) );
  INV_X1 U4225 ( .A(mX1[62]), .ZN(n1864) );
  INV_X1 U4226 ( .A(mX4[63]), .ZN(n2056) );
  INV_X1 U4227 ( .A(mX2[63]), .ZN(n1927) );
  OAI21_X1 U4228 ( .B1(mX3[63]), .B2(n2056), .A(n2833), .ZN(n2832) );
  OAI221_X1 U4229 ( .B1(mX4[62]), .B2(n1993), .C1(mX4[63]), .C2(n1992), .A(
        n2834), .ZN(n2833) );
  OAI21_X1 U4230 ( .B1(mX3[62]), .B2(n2057), .A(n2835), .ZN(n2834) );
  OAI21_X1 U4231 ( .B1(mX1[63]), .B2(n1927), .A(n2897), .ZN(n2543) );
  OAI221_X1 U4232 ( .B1(mX2[62]), .B2(n1864), .C1(mX2[63]), .C2(n1863), .A(
        n2898), .ZN(n2897) );
  OAI21_X1 U4233 ( .B1(mX1[62]), .B2(n1928), .A(n2899), .ZN(n2898) );
  INV_X1 U4234 ( .A(mX3[0]), .ZN(n2055) );
  INV_X1 U4235 ( .A(mX1[0]), .ZN(n1926) );
  BUF_X1 U4236 ( .A(n3824), .Z(n3830) );
  BUF_X1 U4237 ( .A(n3830), .Z(n3806) );
  INV_X1 U4238 ( .A(n3621), .ZN(n3610) );
  CLKBUF_X1 U4239 ( .A(n2640), .Z(n3611) );
  OAI22_X1 U4240 ( .A1(n3625), .A2(n3312), .B1(n3671), .B2(n3078), .ZN(N449)
         );
  OAI22_X1 U4241 ( .A1(n3635), .A2(n3299), .B1(n3043), .B2(n3671), .ZN(N311)
         );
  OAI22_X1 U4242 ( .A1(n3664), .A2(n3304), .B1(n3671), .B2(n2337), .ZN(N281)
         );
  OAI22_X1 U4243 ( .A1(n3628), .A2(n3346), .B1(n3040), .B2(n3470), .ZN(N317)
         );
  OAI22_X1 U4244 ( .A1(n3640), .A2(n3069), .B1(n3289), .B2(n3469), .ZN(N446)
         );
  OAI22_X1 U4245 ( .A1(n3643), .A2(n3080), .B1(n3328), .B2(n3470), .ZN(N469)
         );
  OAI22_X1 U4246 ( .A1(n3631), .A2(n3189), .B1(n3076), .B2(n3469), .ZN(N303)
         );
  OAI22_X1 U4247 ( .A1(n3647), .A2(n3143), .B1(n3228), .B2(n2972), .ZN(N448)
         );
  OAI22_X1 U4248 ( .A1(n3629), .A2(n3019), .B1(n3172), .B2(n2972), .ZN(N456)
         );
  OAI22_X1 U4249 ( .A1(n3625), .A2(n3324), .B1(n3072), .B2(n3481), .ZN(N437)
         );
  CLKBUF_X1 U4250 ( .A(n2640), .Z(n3672) );
  BUF_X1 U4251 ( .A(n3825), .Z(n3815) );
  CLKBUF_X1 U4252 ( .A(n2640), .Z(n3612) );
  BUF_X1 U4253 ( .A(n3822), .Z(n3811) );
  BUF_X2 U4254 ( .A(n3832), .Z(n3818) );
  BUF_X1 U4255 ( .A(n3614), .Z(n3812) );
  INV_X1 U4256 ( .A(n3831), .ZN(n3805) );
  INV_X1 U4257 ( .A(n3612), .ZN(n3613) );
  OAI22_X1 U4258 ( .A1(n3632), .A2(n3228), .B1(n3143), .B2(n3670), .ZN(N320)
         );
  OAI22_X1 U4259 ( .A1(n3641), .A2(n3072), .B1(n3324), .B2(n3622), .ZN(N309)
         );
  OAI22_X1 U4260 ( .A1(n3626), .A2(n3144), .B1(n3229), .B2(n3670), .ZN(N436)
         );
  BUF_X1 U4261 ( .A(n3835), .Z(n3614) );
  CLKBUF_X1 U4262 ( .A(n2640), .Z(n3615) );
  CLKBUF_X1 U4263 ( .A(n2640), .Z(n3616) );
  BUF_X1 U4264 ( .A(n3833), .Z(n3825) );
  BUF_X1 U4265 ( .A(n3833), .Z(n3827) );
  INV_X1 U4266 ( .A(n3822), .ZN(n3618) );
  INV_X1 U4267 ( .A(n3831), .ZN(n3619) );
  INV_X1 U4268 ( .A(n3672), .ZN(n3620) );
  CLKBUF_X1 U4269 ( .A(n2640), .Z(n3735) );
  BUF_X1 U4270 ( .A(n3825), .Z(n3807) );
  OAI22_X1 U4271 ( .A1(rC7[59]), .A2(n3203), .B1(rC7[58]), .B2(n3125), .ZN(
        n2549) );
  OAI22_X1 U4272 ( .A1(n3647), .A2(n3136), .B1(n3195), .B2(n3622), .ZN(N440)
         );
  INV_X1 U4273 ( .A(n3834), .ZN(n3621) );
  INV_X1 U4274 ( .A(n3794), .ZN(n3832) );
  INV_X1 U4275 ( .A(n3794), .ZN(n3831) );
  BUF_X2 U4276 ( .A(n3835), .Z(n3823) );
  INV_X1 U4277 ( .A(n3794), .ZN(n3834) );
  INV_X1 U4278 ( .A(n3614), .ZN(n3796) );
  BUF_X1 U4279 ( .A(n3614), .Z(n3821) );
  BUF_X1 U4280 ( .A(n3823), .Z(n3820) );
  BUF_X1 U4281 ( .A(n3824), .Z(n3829) );
  OAI22_X1 U4282 ( .A1(n3343), .A2(n3619), .B1(n3808), .B2(n3038), .ZN(N662)
         );
  OAI22_X1 U4283 ( .A1(n3147), .A2(n3618), .B1(n3610), .B2(n3203), .ZN(N660)
         );
  OAI22_X1 U4284 ( .A1(n3237), .A2(n3795), .B1(n3617), .B2(n3125), .ZN(N659)
         );
  OAI22_X1 U4285 ( .A1(n3275), .A2(n3619), .B1(n3610), .B2(n3024), .ZN(N658)
         );
  OAI22_X1 U4286 ( .A1(n3098), .A2(n3796), .B1(n3810), .B2(n3175), .ZN(N653)
         );
  OAI22_X1 U4287 ( .A1(n3058), .A2(n3805), .B1(n3821), .B2(n3191), .ZN(N543)
         );
  OAI22_X1 U4288 ( .A1(n3095), .A2(n3804), .B1(n3821), .B2(n3286), .ZN(N544)
         );
  OAI22_X1 U4289 ( .A1(n3131), .A2(n3805), .B1(n3826), .B2(n3254), .ZN(N541)
         );
  BUF_X1 U4290 ( .A(n3830), .Z(n3809) );
  BUF_X4 U4291 ( .A(n2640), .Z(n3622) );
  OAI22_X1 U4292 ( .A1(n3642), .A2(n3242), .B1(n2984), .B2(n3157), .ZN(N280)
         );
  OAI22_X1 U4293 ( .A1(n3120), .A2(n3804), .B1(n3821), .B2(n3204), .ZN(N545)
         );
  AOI22_X1 U4294 ( .A1(n3064), .A2(rC6[9]), .B1(n3204), .B2(rC6[8]), .ZN(n2609) );
  INV_X1 U4295 ( .A(n3794), .ZN(n3833) );
  OAI22_X1 U4296 ( .A1(n3087), .A2(n3799), .B1(n3806), .B2(n3182), .ZN(N615)
         );
  OAI22_X1 U4297 ( .A1(n3063), .A2(n3445), .B1(n3817), .B2(n3276), .ZN(N567)
         );
  OAI22_X1 U4298 ( .A1(n3099), .A2(n3795), .B1(n3609), .B2(n3193), .ZN(N555)
         );
  OAI22_X1 U4299 ( .A1(n3186), .A2(n3803), .B1(n3813), .B2(n3677), .ZN(N611)
         );
  OAI211_X1 U4300 ( .C1(rC7[37]), .C2(n3219), .A(n2583), .B(n2633), .ZN(n2577)
         );
  OAI22_X1 U4301 ( .A1(n3133), .A2(n3796), .B1(n3819), .B2(n3213), .ZN(N656)
         );
  INV_X1 U4302 ( .A(n3616), .ZN(n3623) );
  AND3_X1 U4303 ( .A1(rC7[7]), .A2(n3095), .A3(n2609), .ZN(n2625) );
  INV_X1 U4304 ( .A(n3615), .ZN(n3624) );
  AOI21_X1 U4305 ( .B1(rC6[24]), .B2(n3054), .A(n2629), .ZN(n2628) );
  NOR2_X1 U4306 ( .A1(n3054), .A2(rC6[24]), .ZN(n2630) );
  BUF_X1 U4307 ( .A(n3835), .Z(n3824) );
  OAI22_X1 U4308 ( .A1(n3127), .A2(n3795), .B1(n3819), .B2(n3217), .ZN(N553)
         );
  OAI22_X1 U4309 ( .A1(n3215), .A2(n3798), .B1(n3610), .B2(n3123), .ZN(N657)
         );
  OAI22_X1 U4310 ( .A1(n3686), .A2(n3803), .B1(n3808), .B2(n3678), .ZN(N612)
         );
  OAI22_X1 U4311 ( .A1(n3216), .A2(n3795), .B1(n3808), .B2(n3135), .ZN(N655)
         );
  OAI22_X1 U4312 ( .A1(n3258), .A2(n3795), .B1(n3819), .B2(n3008), .ZN(N552)
         );
  OAI22_X1 U4313 ( .A1(n3632), .A2(n3137), .B1(n3197), .B2(n3459), .ZN(N464)
         );
  OAI22_X1 U4314 ( .A1(n3182), .A2(n3804), .B1(n3821), .B2(n3087), .ZN(N551)
         );
  OAI22_X1 U4315 ( .A1(n3649), .A2(n3044), .B1(n3302), .B2(n2984), .ZN(N463)
         );
  OAI22_X1 U4316 ( .A1(n3805), .A2(n3347), .B1(n3812), .B2(n3683), .ZN(N601)
         );
  OAI22_X1 U4317 ( .A1(n3278), .A2(n3797), .B1(n3018), .B2(n3816), .ZN(N565)
         );
  OAI22_X1 U4318 ( .A1(n3403), .A2(n3797), .B1(n3820), .B2(n3284), .ZN(N614)
         );
  OAI22_X1 U4319 ( .A1(n3641), .A2(n3145), .B1(n3230), .B2(n3671), .ZN(N460)
         );
  OAI22_X1 U4320 ( .A1(n3740), .A2(n3030), .B1(n3287), .B2(n3670), .ZN(N459)
         );
  OAI22_X1 U4321 ( .A1(n3208), .A2(n3797), .B1(n3817), .B2(n3119), .ZN(N566)
         );
  OAI22_X1 U4322 ( .A1(n3148), .A2(n3799), .B1(n3828), .B2(n3249), .ZN(N564)
         );
  OAI22_X1 U4323 ( .A1(n3218), .A2(n3795), .B1(n3807), .B2(n3128), .ZN(N661)
         );
  OAI22_X1 U4324 ( .A1(n3795), .A2(n3046), .B1(n3818), .B2(n3268), .ZN(N554)
         );
  OAI22_X1 U4325 ( .A1(n3664), .A2(n3155), .B1(n3240), .B2(n3459), .ZN(N462)
         );
  OAI22_X1 U4326 ( .A1(n3642), .A2(n3029), .B1(n3331), .B2(n3459), .ZN(N435)
         );
  OAI22_X1 U4327 ( .A1(n3026), .A2(n3618), .B1(n3828), .B2(n3280), .ZN(N654)
         );
  OAI22_X1 U4328 ( .A1(n3668), .A2(n3305), .B1(n3051), .B2(n3470), .ZN(N465)
         );
  OAI22_X1 U4329 ( .A1(n3284), .A2(n3804), .B1(n3820), .B2(n3403), .ZN(N550)
         );
  OAI22_X1 U4330 ( .A1(n3650), .A2(n3252), .B1(n2336), .B2(n3469), .ZN(N282)
         );
  OAI22_X1 U4331 ( .A1(n3638), .A2(n3083), .B1(n3293), .B2(n3670), .ZN(N466)
         );
  OAI22_X1 U4332 ( .A1(n3634), .A2(n3139), .B1(n2984), .B2(n3348), .ZN(N279)
         );
  OAI22_X1 U4333 ( .A1(n3740), .A2(n3078), .B1(n3312), .B2(n3670), .ZN(N321)
         );
  OAI22_X1 U4334 ( .A1(n2978), .A2(n3185), .B1(n3459), .B2(n3107), .ZN(N283)
         );
  OAI22_X1 U4335 ( .A1(n2979), .A2(n3068), .B1(n3291), .B2(n3670), .ZN(N450)
         );
  OAI22_X1 U4336 ( .A1(n3641), .A2(n3334), .B1(n3033), .B2(n2972), .ZN(N284)
         );
  OAI22_X1 U4337 ( .A1(n3654), .A2(n2327), .B1(n2183), .B2(n3671), .ZN(N419)
         );
  OAI22_X1 U4338 ( .A1(n3657), .A2(n3011), .B1(n3262), .B2(n3470), .ZN(N467)
         );
  OAI22_X1 U4339 ( .A1(n3740), .A2(n3141), .B1(n3206), .B2(n3670), .ZN(N468)
         );
  OAI22_X1 U4340 ( .A1(n3634), .A2(n3167), .B1(n3469), .B2(n3248), .ZN(N285)
         );
  OAI22_X1 U4341 ( .A1(n3641), .A2(n3325), .B1(n3472), .B2(n3073), .ZN(N461)
         );
  OAI22_X1 U4342 ( .A1(n3642), .A2(n3040), .B1(n3473), .B2(n3346), .ZN(N445)
         );
  OAI211_X1 U4343 ( .C1(n2708), .C2(n2709), .A(n2699), .B(n2710), .ZN(n2693)
         );
  OAI211_X1 U4344 ( .C1(rC2[9]), .C2(n3090), .A(n2700), .B(n2701), .ZN(n2698)
         );
  INV_X1 U4345 ( .A(n2704), .ZN(n2259) );
  OAI22_X1 U4346 ( .A1(n3627), .A2(n3153), .B1(n3245), .B2(n3469), .ZN(N444)
         );
  OAI22_X1 U4347 ( .A1(n3780), .A2(n3041), .B1(n3308), .B2(n3390), .ZN(N384)
         );
  OAI22_X1 U4348 ( .A1(n3422), .A2(n3181), .B1(n3105), .B2(n3761), .ZN(N385)
         );
  OAI22_X1 U4349 ( .A1(n3763), .A2(n3010), .B1(n3261), .B2(n3754), .ZN(N531)
         );
  OAI22_X1 U4350 ( .A1(n3428), .A2(n3158), .B1(n3243), .B2(n3380), .ZN(N383)
         );
  OAI22_X1 U4351 ( .A1(n3774), .A2(n3177), .B1(n3017), .B2(n3754), .ZN(N507)
         );
  INV_X1 U4352 ( .A(n2544), .ZN(n3835) );
  OAI22_X1 U4353 ( .A1(n3776), .A2(n3224), .B1(n3121), .B2(n3380), .ZN(N382)
         );
  OAI22_X1 U4354 ( .A1(n2986), .A2(n3333), .B1(n3032), .B2(n3373), .ZN(N509)
         );
  OAI22_X1 U4355 ( .A1(n3763), .A2(n3081), .B1(n3327), .B2(n3752), .ZN(N533)
         );
  OAI22_X1 U4356 ( .A1(n3422), .A2(n3190), .B1(n3106), .B2(n3372), .ZN(N508)
         );
  OAI22_X1 U4357 ( .A1(n3427), .A2(n3140), .B1(n3207), .B2(n3752), .ZN(N532)
         );
  OAI22_X1 U4358 ( .A1(n3776), .A2(n3032), .B1(n3333), .B2(n3756), .ZN(N381)
         );
  OAI22_X1 U4359 ( .A1(n3427), .A2(n3082), .B1(n3292), .B2(n3372), .ZN(N530)
         );
  OAI22_X1 U4360 ( .A1(n3777), .A2(n3319), .B1(n3088), .B2(n3372), .ZN(N506)
         );
  OAI22_X1 U4361 ( .A1(n3776), .A2(n3106), .B1(n3190), .B2(n3391), .ZN(N380)
         );
  OAI22_X1 U4362 ( .A1(n3783), .A2(n3455), .B1(n3391), .B2(n3349), .ZN(N343)
         );
  OAI22_X1 U4363 ( .A1(n3784), .A2(n3109), .B1(n3201), .B2(n3390), .ZN(N349)
         );
  OAI22_X1 U4364 ( .A1(n3784), .A2(n3047), .B1(n3311), .B2(n3391), .ZN(N348)
         );
  OAI22_X1 U4365 ( .A1(n3783), .A2(n3152), .B1(n3236), .B2(n3386), .ZN(N347)
         );
  OAI22_X1 U4366 ( .A1(n3783), .A2(n3332), .B1(n3450), .B2(n2990), .ZN(N346)
         );
  OAI22_X1 U4367 ( .A1(n3783), .A2(n3381), .B1(n3758), .B2(n3471), .ZN(N345)
         );
  OAI22_X1 U4368 ( .A1(n3783), .A2(n3480), .B1(n3339), .B2(n3756), .ZN(N344)
         );
  OAI22_X1 U4369 ( .A1(n3777), .A2(n3017), .B1(n3177), .B2(n3386), .ZN(N379)
         );
  OAI22_X1 U4370 ( .A1(n3772), .A2(n3300), .B1(n3050), .B2(n3372), .ZN(N529)
         );
  OAI22_X1 U4371 ( .A1(n3428), .A2(n3048), .B1(n3342), .B2(n3752), .ZN(N505)
         );
  OAI22_X1 U4372 ( .A1(n3780), .A2(n3088), .B1(n3319), .B2(n3757), .ZN(N378)
         );
  OAI22_X1 U4373 ( .A1(n3781), .A2(n3138), .B1(n3196), .B2(n3373), .ZN(N528)
         );
  OAI22_X1 U4374 ( .A1(n3773), .A2(n3164), .B1(n3225), .B2(n3752), .ZN(N504)
         );
  OAI22_X1 U4375 ( .A1(n3780), .A2(n3342), .B1(n3048), .B2(n3761), .ZN(N377)
         );
  OAI22_X1 U4376 ( .A1(n3780), .A2(n3225), .B1(n3758), .B2(n3164), .ZN(N376)
         );
  OAI22_X1 U4377 ( .A1(n3781), .A2(n3260), .B1(n3012), .B2(n3760), .ZN(N361)
         );
  OAI22_X1 U4378 ( .A1(n3781), .A2(n3295), .B1(n3085), .B2(n3760), .ZN(N360)
         );
  OAI22_X1 U4379 ( .A1(n3781), .A2(n3112), .B1(n3223), .B2(n3760), .ZN(N359)
         );
  OAI22_X1 U4380 ( .A1(n3781), .A2(n3497), .B1(n3464), .B2(n3760), .ZN(N358)
         );
  OAI22_X1 U4381 ( .A1(n3780), .A2(n3108), .B1(n3760), .B2(n3198), .ZN(N356)
         );
  OAI22_X1 U4382 ( .A1(n3784), .A2(n3490), .B1(n3760), .B2(n2263), .ZN(N354)
         );
  OAI22_X1 U4383 ( .A1(n2994), .A2(n3142), .B1(n3760), .B2(n3241), .ZN(N353)
         );
  OAI22_X1 U4384 ( .A1(n3784), .A2(n3322), .B1(n3760), .B2(n3090), .ZN(N352)
         );
  OAI22_X1 U4385 ( .A1(n3784), .A2(n3310), .B1(n3760), .B2(n2266), .ZN(N351)
         );
  OAI22_X1 U4386 ( .A1(n3784), .A2(n3246), .B1(n3760), .B2(n3169), .ZN(N350)
         );
  OAI22_X1 U4387 ( .A1(n3762), .A2(n3045), .B1(n3301), .B2(n3758), .ZN(N527)
         );
  OAI22_X1 U4388 ( .A1(n3779), .A2(n3086), .B1(n3335), .B2(n3761), .ZN(N375)
         );
  AOI221_X1 U4389 ( .B1(n2675), .B2(n2676), .C1(n3398), .C2(n2677), .A(n2678), 
        .ZN(n2674) );
  OAI22_X1 U4390 ( .A1(n2985), .A2(n3156), .B1(n3239), .B2(n3386), .ZN(N526)
         );
  BUF_X1 U4391 ( .A(n3448), .Z(n3631) );
  BUF_X1 U4392 ( .A(n3623), .Z(n3632) );
  BUF_X1 U4393 ( .A(n3448), .Z(n3633) );
  BUF_X1 U4394 ( .A(n3623), .Z(n3636) );
  BUF_X1 U4395 ( .A(n3625), .Z(n3638) );
  BUF_X1 U4396 ( .A(n3475), .Z(n3640) );
  BUF_X1 U4397 ( .A(n3746), .Z(n3644) );
  BUF_X1 U4398 ( .A(n3748), .Z(n3645) );
  BUF_X1 U4399 ( .A(n3746), .Z(n3646) );
  BUF_X1 U4400 ( .A(n3625), .Z(n3648) );
  BUF_X1 U4401 ( .A(n3747), .Z(n3649) );
  BUF_X1 U4402 ( .A(n3476), .Z(n3650) );
  BUF_X1 U4403 ( .A(n3743), .Z(n3651) );
  BUF_X1 U4404 ( .A(n3748), .Z(n3652) );
  BUF_X1 U4405 ( .A(n3741), .Z(n3653) );
  BUF_X1 U4406 ( .A(n3744), .Z(n3655) );
  BUF_X1 U4407 ( .A(n3623), .Z(n3657) );
  BUF_X1 U4408 ( .A(n3745), .Z(n3658) );
  BUF_X1 U4409 ( .A(n3737), .Z(n3659) );
  BUF_X1 U4410 ( .A(n3476), .Z(n3660) );
  BUF_X1 U4411 ( .A(n3476), .Z(n3661) );
  BUF_X1 U4412 ( .A(n3738), .Z(n3662) );
  BUF_X1 U4413 ( .A(n3736), .Z(n3663) );
  BUF_X1 U4414 ( .A(n3736), .Z(n3666) );
  BUF_X1 U4415 ( .A(n3625), .Z(n3668) );
  BUF_X1 U4416 ( .A(n3745), .Z(n3669) );
  BUF_X4 U4417 ( .A(n2640), .Z(n3670) );
  OAI221_X4 U4418 ( .B1(n2737), .B2(n2738), .C1(rC1[63]), .C2(n2276), .A(n2739), .ZN(n2640) );
  INV_X1 U4419 ( .A(n2640), .ZN(n3750) );
  INV_X1 U4420 ( .A(n2640), .ZN(n3749) );
  BUF_X1 U4421 ( .A(n3613), .Z(n3744) );
  BUF_X1 U4422 ( .A(n3491), .Z(n3745) );
  OAI22_X1 U4423 ( .A1(n3646), .A2(n3007), .B1(n3290), .B2(n3671), .ZN(N434)
         );
  OAI211_X1 U4424 ( .C1(rC3[12]), .C2(n2183), .A(n2179), .B(n2805), .ZN(n2789)
         );
  OAI22_X1 U4425 ( .A1(n3644), .A2(n3340), .B1(n3093), .B2(n3473), .ZN(N299)
         );
  AOI22_X1 U4426 ( .A1(rC3[7]), .A2(n3420), .B1(rC3[8]), .B2(n3606), .ZN(n2794) );
  OAI22_X1 U4427 ( .A1(n3665), .A2(n3073), .B1(n3325), .B2(n3671), .ZN(N333)
         );
  OAI22_X1 U4428 ( .A1(n3629), .A2(n3230), .B1(n3145), .B2(n3671), .ZN(N332)
         );
  OAI22_X1 U4429 ( .A1(n3663), .A2(n3287), .B1(n3030), .B2(n2983), .ZN(N331)
         );
  OAI22_X1 U4430 ( .A1(n3736), .A2(n3056), .B1(n3320), .B2(n2970), .ZN(N330)
         );
  OAI22_X1 U4431 ( .A1(n3641), .A2(n3313), .B1(n3065), .B2(n3671), .ZN(N329)
         );
  OAI22_X1 U4432 ( .A1(n3649), .A2(n3172), .B1(n3019), .B2(n3622), .ZN(N328)
         );
  OAI22_X1 U4433 ( .A1(n3652), .A2(n3187), .B1(n3102), .B2(n3469), .ZN(N327)
         );
  OAI22_X1 U4434 ( .A1(n3639), .A2(n3021), .B1(n3314), .B2(n3622), .ZN(N326)
         );
  OAI22_X1 U4435 ( .A1(n3739), .A2(n3113), .B1(n3232), .B2(n2984), .ZN(N325)
         );
  OAI22_X1 U4436 ( .A1(n3649), .A2(n3226), .B1(n3165), .B2(n3670), .ZN(N324)
         );
  OAI22_X1 U4437 ( .A1(n3648), .A2(n3162), .B1(n3221), .B2(n2984), .ZN(N323)
         );
  OAI22_X1 U4438 ( .A1(n3653), .A2(n3291), .B1(n3068), .B2(n3459), .ZN(N322)
         );
  INV_X1 U4439 ( .A(n2804), .ZN(n2192) );
  OAI22_X1 U4440 ( .A1(n3650), .A2(n3238), .B1(n3154), .B2(n3670), .ZN(N310)
         );
  OAI22_X1 U4441 ( .A1(n3781), .A2(n3463), .B1(n2260), .B2(n3760), .ZN(N357)
         );
  OAI22_X1 U4442 ( .A1(n3769), .A2(n3074), .B1(n3326), .B2(n3391), .ZN(N397)
         );
  OAI22_X1 U4443 ( .A1(n3775), .A2(n3231), .B1(n3146), .B2(n3757), .ZN(N396)
         );
  OAI22_X1 U4444 ( .A1(n3772), .A2(n3288), .B1(n3031), .B2(n3386), .ZN(N395)
         );
  OAI22_X1 U4445 ( .A1(n3772), .A2(n3057), .B1(n3323), .B2(n3380), .ZN(N394)
         );
  OAI22_X1 U4446 ( .A1(n3774), .A2(n3315), .B1(n3067), .B2(n3390), .ZN(N393)
         );
  OAI22_X1 U4447 ( .A1(n3774), .A2(n3307), .B1(n3020), .B2(n2993), .ZN(N392)
         );
  OAI22_X1 U4448 ( .A1(n3775), .A2(n3188), .B1(n3103), .B2(n3390), .ZN(N391)
         );
  OAI22_X1 U4449 ( .A1(n3778), .A2(n3022), .B1(n3316), .B2(n3757), .ZN(N390)
         );
  OAI22_X1 U4450 ( .A1(n3429), .A2(n3114), .B1(n3233), .B2(n3761), .ZN(N389)
         );
  OAI22_X1 U4451 ( .A1(n3775), .A2(n3227), .B1(n3758), .B2(n3166), .ZN(N388)
         );
  OAI22_X1 U4452 ( .A1(n3766), .A2(n3163), .B1(n3222), .B2(n3756), .ZN(N387)
         );
  OAI22_X1 U4453 ( .A1(n3766), .A2(n3297), .B1(n3070), .B2(n3756), .ZN(N386)
         );
  OAI211_X1 U4454 ( .C1(rC4[7]), .C2(n3246), .A(n2259), .B(n2702), .ZN(n2694)
         );
  AOI22_X1 U4455 ( .A1(rC4[13]), .A2(n3108), .B1(n3483), .B2(n3500), .ZN(n2695) );
  BUF_X2 U4456 ( .A(n2544), .Z(n3794) );
  OAI22_X1 U4457 ( .A1(n2999), .A2(n3805), .B1(n3826), .B2(n3687), .ZN(N539)
         );
  OAI22_X1 U4458 ( .A1(n3779), .A2(n3180), .B1(n3104), .B2(n3761), .ZN(N374)
         );
  OAI22_X1 U4459 ( .A1(n3779), .A2(n3110), .B1(n3220), .B2(n3759), .ZN(N373)
         );
  OAI22_X1 U4460 ( .A1(n3779), .A2(n3042), .B1(n3309), .B2(n3759), .ZN(N372)
         );
  OAI22_X1 U4461 ( .A1(n3779), .A2(n3159), .B1(n3244), .B2(n3759), .ZN(N371)
         );
  OAI22_X1 U4462 ( .A1(n3778), .A2(n3176), .B1(n3122), .B2(n3759), .ZN(N370)
         );
  OAI22_X1 U4463 ( .A1(n3778), .A2(n3317), .B1(n3066), .B2(n3759), .ZN(N369)
         );
  OAI22_X1 U4464 ( .A1(n3778), .A2(n3170), .B1(n3184), .B2(n3759), .ZN(N368)
         );
  OAI22_X1 U4465 ( .A1(n3778), .A2(n3303), .B1(n3059), .B2(n3373), .ZN(N367)
         );
  OAI22_X1 U4466 ( .A1(n3782), .A2(n3023), .B1(n3318), .B2(n3759), .ZN(N366)
         );
  OAI22_X1 U4467 ( .A1(n3782), .A2(n3115), .B1(n3234), .B2(n3759), .ZN(N365)
         );
  OAI22_X1 U4468 ( .A1(n3782), .A2(n3336), .B1(n3034), .B2(n3759), .ZN(N364)
         );
  OAI22_X1 U4469 ( .A1(n3782), .A2(n3253), .B1(n3111), .B2(n3759), .ZN(N363)
         );
  OAI22_X1 U4470 ( .A1(n3782), .A2(n3094), .B1(n3341), .B2(n3759), .ZN(N362)
         );
  INV_X1 U4471 ( .A(n3679), .ZN(n3675) );
  OAI22_X1 U4472 ( .A1(n3674), .A2(n3805), .B1(n3821), .B2(n3259), .ZN(N542)
         );
  OAI22_X1 U4473 ( .A1(n3780), .A2(n3478), .B1(n3756), .B2(n3498), .ZN(N355)
         );
  OAI22_X1 U4474 ( .A1(n3784), .A2(n3471), .B1(n3381), .B2(n3757), .ZN(N473)
         );
  OAI22_X1 U4475 ( .A1(n3784), .A2(n3339), .B1(n3480), .B2(n3380), .ZN(N472)
         );
  OAI22_X1 U4476 ( .A1(n3770), .A2(n3337), .B1(n3077), .B2(n3390), .ZN(N406)
         );
  OAI22_X1 U4477 ( .A1(n3770), .A2(n3327), .B1(n3081), .B2(n3391), .ZN(N405)
         );
  OAI22_X1 U4478 ( .A1(n3771), .A2(n3207), .B1(n3140), .B2(n3380), .ZN(N404)
         );
  OAI22_X1 U4479 ( .A1(n3770), .A2(n3261), .B1(n3010), .B2(n3757), .ZN(N403)
         );
  OAI22_X1 U4480 ( .A1(n3777), .A2(n3292), .B1(n3758), .B2(n3082), .ZN(N402)
         );
  OAI22_X1 U4481 ( .A1(n2986), .A2(n3050), .B1(n3758), .B2(n3300), .ZN(N401)
         );
  OAI22_X1 U4482 ( .A1(n3766), .A2(n3196), .B1(n3138), .B2(n3386), .ZN(N400)
         );
  OAI22_X1 U4483 ( .A1(n3769), .A2(n3301), .B1(n3045), .B2(n3757), .ZN(N399)
         );
  OAI22_X1 U4484 ( .A1(n3772), .A2(n3239), .B1(n3156), .B2(n3386), .ZN(N398)
         );
  OAI22_X1 U4485 ( .A1(n3771), .A2(n3349), .B1(n3455), .B2(n3390), .ZN(N471)
         );
  AOI21_X1 U4486 ( .B1(n3490), .B2(rC4[11]), .A(n2707), .ZN(n2700) );
  OAI22_X1 U4487 ( .A1(n3765), .A2(n3326), .B1(n3074), .B2(n3380), .ZN(N525)
         );
  AOI22_X1 U4488 ( .A1(n3450), .A2(rC2[3]), .B1(n3486), .B2(rC2[2]), .ZN(n2715) );
  INV_X1 U4489 ( .A(n2715), .ZN(n2271) );
  OAI22_X1 U4490 ( .A1(n3429), .A2(n3146), .B1(n3231), .B2(n3756), .ZN(N524)
         );
  OAI22_X1 U4491 ( .A1(rC4[15]), .A2(n3497), .B1(rC4[14]), .B2(n3500), .ZN(
        n2696) );
  OAI22_X1 U4492 ( .A1(n3676), .A2(n3805), .B1(n3820), .B2(n3345), .ZN(N538)
         );
  AOI22_X1 U4493 ( .A1(n3058), .A2(rC7[6]), .B1(n3674), .B2(rC7[5]), .ZN(n3680) );
  OAI22_X1 U4494 ( .A1(n3651), .A2(n3379), .B1(n2181), .B2(n3670), .ZN(N421)
         );
  OAI22_X1 U4495 ( .A1(n3383), .A2(n3447), .B1(rC1[13]), .B2(n3211), .ZN(n2785) );
  AOI22_X1 U4496 ( .A1(n3416), .A2(rC1[15]), .B1(n3447), .B2(rC1[14]), .ZN(
        n2784) );
  AOI211_X1 U4497 ( .C1(n3402), .C2(rC7[12]), .A(rC7[11]), .B(n3678), .ZN(
        n3682) );
  AOI22_X1 U4498 ( .A1(n3058), .A2(rC7[6]), .B1(n3674), .B2(rC7[5]), .ZN(n2613) );
  OAI211_X1 U4499 ( .C1(rC4[12]), .C2(n3478), .A(n2705), .B(n2706), .ZN(n2704)
         );
  AOI21_X1 U4500 ( .B1(rC2[13]), .B2(n3198), .A(n2696), .ZN(n2706) );
  NOR2_X1 U4501 ( .A1(rC2[12]), .A2(n3498), .ZN(n2707) );
  OAI22_X1 U4502 ( .A1(n3428), .A2(n3031), .B1(n3288), .B2(n3391), .ZN(N523)
         );
  OAI22_X1 U4503 ( .A1(n3679), .A2(n3805), .B1(n3820), .B2(n3685), .ZN(N540)
         );
  OAI211_X1 U4504 ( .C1(rC7[7]), .C2(n3095), .A(n2609), .B(n2612), .ZN(n2611)
         );
  AOI22_X1 U4505 ( .A1(n3680), .A2(n2614), .B1(rC6[6]), .B2(n3191), .ZN(n2612)
         );
  OAI22_X1 U4506 ( .A1(rC7[5]), .A2(n3674), .B1(rC7[4]), .B2(n3131), .ZN(n2614) );
  INV_X1 U4507 ( .A(n2806), .ZN(n2179) );
  OAI21_X1 U4508 ( .B1(n3118), .B2(rC3[13]), .A(n2784), .ZN(n2806) );
  OAI22_X1 U4509 ( .A1(n3064), .A2(n3803), .B1(n3819), .B2(n3277), .ZN(N610)
         );
  OAI22_X1 U4510 ( .A1(n3025), .A2(n3797), .B1(n3826), .B2(n3344), .ZN(N563)
         );
  OAI22_X1 U4511 ( .A1(n3655), .A2(n3171), .B1(n2987), .B2(n3256), .ZN(N298)
         );
  OAI22_X1 U4512 ( .A1(n3677), .A2(n3804), .B1(n3812), .B2(n3186), .ZN(N547)
         );
  OAI22_X1 U4513 ( .A1(n3277), .A2(n3804), .B1(n3819), .B2(n3064), .ZN(N546)
         );
  OAI22_X1 U4514 ( .A1(n3678), .A2(n3804), .B1(n3808), .B2(n3686), .ZN(N548)
         );
  OAI22_X1 U4515 ( .A1(n3204), .A2(n3449), .B1(n3818), .B2(n3120), .ZN(N609)
         );
  OAI22_X1 U4516 ( .A1(n3071), .A2(n3619), .B1(n3828), .B2(n3274), .ZN(N562)
         );
  OAI22_X1 U4517 ( .A1(n3250), .A2(n3618), .B1(n3808), .B2(n3160), .ZN(N652)
         );
  OAI22_X1 U4518 ( .A1(n3286), .A2(n3799), .B1(n3811), .B2(n3095), .ZN(N608)
         );
  OAI22_X1 U4519 ( .A1(n3266), .A2(n3619), .B1(n3609), .B2(n3054), .ZN(N561)
         );
  OAI221_X1 U4520 ( .B1(n3139), .B2(rC3[0]), .C1(n3242), .C2(rC3[1]), .A(n2802), .ZN(n2804) );
  OAI22_X1 U4521 ( .A1(n3281), .A2(n3618), .B1(n3494), .B2(n3027), .ZN(N651)
         );
  OAI22_X1 U4522 ( .A1(n3096), .A2(n3795), .B1(n3807), .B2(n3173), .ZN(N650)
         );
  OAI22_X1 U4523 ( .A1(n3199), .A2(n3799), .B1(n3812), .B2(n3100), .ZN(N649)
         );
  OAI22_X1 U4524 ( .A1(n3269), .A2(n3797), .B1(n3818), .B2(n3035), .ZN(N648)
         );
  OAI22_X1 U4525 ( .A1(n3212), .A2(n3618), .B1(n3810), .B2(n3124), .ZN(N647)
         );
  OAI22_X1 U4526 ( .A1(n3251), .A2(n3795), .B1(n3817), .B2(n3161), .ZN(N646)
         );
  OAI22_X1 U4527 ( .A1(n3282), .A2(n3621), .B1(n3494), .B2(n3039), .ZN(N645)
         );
  OAI22_X1 U4528 ( .A1(n3097), .A2(n3799), .B1(n3828), .B2(n3174), .ZN(N644)
         );
  OAI22_X1 U4529 ( .A1(n3200), .A2(n3796), .B1(n3609), .B2(n3101), .ZN(N643)
         );
  OAI22_X1 U4530 ( .A1(n3270), .A2(n3618), .B1(n3806), .B2(n3036), .ZN(N642)
         );
  OAI22_X1 U4531 ( .A1(n3205), .A2(n3795), .B1(n3828), .B2(n3129), .ZN(N641)
         );
  OAI22_X1 U4532 ( .A1(n3062), .A2(n3796), .B1(n3808), .B2(n3265), .ZN(N640)
         );
  OAI22_X1 U4533 ( .A1(n3191), .A2(n3797), .B1(n3811), .B2(n3058), .ZN(N607)
         );
  OAI22_X1 U4534 ( .A1(n3061), .A2(n3803), .B1(n3819), .B2(n3272), .ZN(N560)
         );
  OAI22_X1 U4535 ( .A1(n3259), .A2(n3803), .B1(n3811), .B2(n3674), .ZN(N606)
         );
  OAI22_X1 U4536 ( .A1(n3016), .A2(n3799), .B1(n3819), .B2(n3279), .ZN(N559)
         );
  OAI22_X1 U4537 ( .A1(n3645), .A2(n3263), .B1(n3013), .B2(n2972), .ZN(N297)
         );
  OAI22_X1 U4538 ( .A1(n3653), .A2(n3294), .B1(n3084), .B2(n3622), .ZN(N296)
         );
  OAI22_X1 U4539 ( .A1(n3639), .A2(n3052), .B1(n3306), .B2(n3622), .ZN(N295)
         );
  OAI22_X1 U4540 ( .A1(n3667), .A2(n3370), .B1(n3416), .B2(n3670), .ZN(N294)
         );
  OAI22_X1 U4541 ( .A1(n3641), .A2(n2181), .B1(n3379), .B2(n3622), .ZN(N293)
         );
  OAI22_X1 U4542 ( .A1(n3660), .A2(n3118), .B1(n3211), .B2(n3469), .ZN(N292)
         );
  OAI22_X1 U4543 ( .A1(n3636), .A2(n2183), .B1(n2327), .B2(n3622), .ZN(N291)
         );
  OAI22_X1 U4544 ( .A1(n3667), .A2(n3296), .B1(n3091), .B2(n3622), .ZN(N290)
         );
  OAI22_X1 U4545 ( .A1(n3669), .A2(n3151), .B1(n2987), .B2(n3247), .ZN(N289)
         );
  OAI22_X1 U4546 ( .A1(n3742), .A2(n3377), .B1(n3374), .B2(n3670), .ZN(N288)
         );
  OAI22_X1 U4547 ( .A1(n3633), .A2(n3388), .B1(n2331), .B2(n3670), .ZN(N287)
         );
  OAI22_X1 U4548 ( .A1(n2979), .A2(n3420), .B1(n3183), .B2(n3670), .ZN(N286)
         );
  NOR3_X1 U4549 ( .A1(n2791), .A2(n2790), .A3(n3418), .ZN(n2788) );
  AOI211_X1 U4550 ( .C1(rC1[7]), .C2(n3183), .A(n3444), .B(n2789), .ZN(n2786)
         );
  AOI22_X1 U4551 ( .A1(rC7[1]), .A2(n3676), .B1(rC7[2]), .B2(n3681), .ZN(n2622) );
  NOR3_X1 U4552 ( .A1(n3431), .A2(rC7[10]), .A3(n3677), .ZN(n3688) );
  NOR3_X1 U4553 ( .A1(n2626), .A2(rC7[10]), .A3(n3677), .ZN(n2621) );
  OAI22_X1 U4554 ( .A1(n3661), .A2(n2337), .B1(n3304), .B2(n3670), .ZN(N409)
         );
  OAI22_X1 U4555 ( .A1(n3668), .A2(n3157), .B1(n3242), .B2(n3622), .ZN(N408)
         );
  OAI22_X1 U4556 ( .A1(n2978), .A2(n3348), .B1(n3139), .B2(n2970), .ZN(N407)
         );
  OAI22_X1 U4557 ( .A1(n3658), .A2(n3338), .B1(n2276), .B2(n2970), .ZN(N342)
         );
  OAI22_X1 U4558 ( .A1(n3657), .A2(n3328), .B1(n3080), .B2(n3670), .ZN(N341)
         );
  OAI22_X1 U4559 ( .A1(n3643), .A2(n3206), .B1(n3141), .B2(n3469), .ZN(N340)
         );
  OAI22_X1 U4560 ( .A1(n2979), .A2(n3262), .B1(n3011), .B2(n2972), .ZN(N339)
         );
  OAI22_X1 U4561 ( .A1(n3644), .A2(n3293), .B1(n3083), .B2(n3670), .ZN(N338)
         );
  OAI22_X1 U4562 ( .A1(n3653), .A2(n3051), .B1(n3305), .B2(n3470), .ZN(N337)
         );
  OAI22_X1 U4563 ( .A1(n3745), .A2(n3197), .B1(n3137), .B2(n3622), .ZN(N336)
         );
  OAI22_X1 U4564 ( .A1(n3302), .A2(n3640), .B1(n3044), .B2(n3670), .ZN(N335)
         );
  OAI22_X1 U4565 ( .A1(n3646), .A2(n3240), .B1(n3155), .B2(n3469), .ZN(N334)
         );
  OAI21_X1 U4566 ( .B1(n2768), .B2(n2769), .A(n2764), .ZN(n2762) );
  AND2_X1 U4567 ( .A1(n2644), .A2(n2645), .ZN(n3689) );
  AND2_X1 U4568 ( .A1(n2646), .A2(n2647), .ZN(n3690) );
  NAND2_X1 U4569 ( .A1(rC2[63]), .A2(n3077), .ZN(n2644) );
  OAI21_X1 U4570 ( .B1(rC2[62]), .B2(n3081), .A(n2731), .ZN(n2645) );
  AOI221_X1 U4571 ( .B1(n3045), .B2(rC2[56]), .C1(n3138), .C2(rC2[57]), .A(
        n2642), .ZN(n2646) );
  OAI22_X1 U4572 ( .A1(rC2[56]), .A2(n3045), .B1(rC2[55]), .B2(n3156), .ZN(
        n2647) );
  AOI21_X1 U4573 ( .B1(rC2[43]), .B2(n3070), .A(n2659), .ZN(n2654) );
  INV_X1 U4574 ( .A(n2659), .ZN(n2213) );
  OAI22_X1 U4575 ( .A1(rC2[44]), .A2(n3222), .B1(rC2[43]), .B2(n3070), .ZN(
        n2656) );
  OAI22_X1 U4576 ( .A1(n3684), .A2(n3797), .B1(n3826), .B2(n3402), .ZN(N613)
         );
  OAI22_X1 U4577 ( .A1(n3402), .A2(n3797), .B1(n3817), .B2(n3684), .ZN(N549)
         );
  AOI22_X1 U4578 ( .A1(n3685), .A2(n3675), .B1(n3000), .B2(n3687), .ZN(n2624)
         );
  NOR2_X1 U4579 ( .A1(n3402), .A2(rC7[12]), .ZN(n2620) );
  OAI22_X1 U4580 ( .A1(n3117), .A2(n3797), .B1(n3819), .B2(n3194), .ZN(N558)
         );
  AOI211_X1 U4581 ( .C1(rC3[9]), .C2(n3419), .A(n2793), .B(n2792), .ZN(n2791)
         );
  OAI22_X1 U4582 ( .A1(rC1[10]), .A2(n3247), .B1(n2794), .B2(n2795), .ZN(n2792) );
  OAI22_X1 U4583 ( .A1(rC3[9]), .A2(n3419), .B1(rC3[8]), .B2(n3606), .ZN(n2795) );
  OAI221_X1 U4584 ( .B1(n2759), .B2(n2760), .C1(n2762), .C2(n2761), .A(n2763), 
        .ZN(n2756) );
  INV_X1 U4585 ( .A(n2639), .ZN(n3793) );
  INV_X1 U4586 ( .A(n3751), .ZN(n3791) );
  OAI221_X1 U4587 ( .B1(n2576), .B2(n2577), .C1(n2579), .C2(n2578), .A(n2580), 
        .ZN(n2571) );
  OAI22_X1 U4588 ( .A1(n3683), .A2(n3619), .B1(n3808), .B2(n3347), .ZN(N537)
         );
  BUF_X2 U4589 ( .A(n3834), .Z(n3819) );
  BUF_X2 U4590 ( .A(n3835), .Z(n3822) );
  OAI22_X1 U4591 ( .A1(n3664), .A2(n3168), .B1(n3469), .B2(n3235), .ZN(N433)
         );
  OAI22_X1 U4592 ( .A1(n2978), .A2(n3321), .B1(n3079), .B2(n3671), .ZN(N432)
         );
  OAI22_X1 U4593 ( .A1(n3644), .A2(n3076), .B1(n3473), .B2(n3189), .ZN(N431)
         );
  OAI22_X1 U4594 ( .A1(n3627), .A2(n3210), .B1(n3150), .B2(n3470), .ZN(N430)
         );
  OAI22_X1 U4595 ( .A1(n3646), .A2(n3329), .B1(n3014), .B2(n3670), .ZN(N429)
         );
  OAI22_X1 U4596 ( .A1(n3645), .A2(n3202), .B1(n3130), .B2(n2983), .ZN(N428)
         );
  OAI22_X1 U4597 ( .A1(n3652), .A2(n3093), .B1(n3340), .B2(n3670), .ZN(N427)
         );
  OAI22_X1 U4598 ( .A1(n3657), .A2(n3256), .B1(n3469), .B2(n3171), .ZN(N426)
         );
  OAI22_X1 U4599 ( .A1(n3662), .A2(n3013), .B1(n3263), .B2(n2983), .ZN(N425)
         );
  OAI22_X1 U4600 ( .A1(n3660), .A2(n3084), .B1(n3294), .B2(n2970), .ZN(N424)
         );
  OAI22_X1 U4601 ( .A1(n3739), .A2(n3306), .B1(n3052), .B2(n3670), .ZN(N423)
         );
  OAI22_X1 U4602 ( .A1(n3659), .A2(n3416), .B1(n3370), .B2(n3472), .ZN(N422)
         );
  AOI211_X1 U4603 ( .C1(n2796), .C2(n2797), .A(n2798), .B(n2790), .ZN(n2787)
         );
  OAI22_X1 U4604 ( .A1(n3285), .A2(n3803), .B1(n3817), .B2(n3092), .ZN(N557)
         );
  OAI211_X1 U4605 ( .C1(rC7[63]), .C2(n3192), .A(n2545), .B(n2546), .ZN(n2544)
         );
  AOI211_X1 U4606 ( .C1(n2650), .C2(n2649), .A(n2651), .B(n2198), .ZN(n2648)
         );
  AOI211_X1 U4607 ( .C1(n2135), .C2(n2750), .A(n2751), .B(n2752), .ZN(n2746)
         );
  OAI211_X1 U4608 ( .C1(rC3[19]), .C2(n3171), .A(n2778), .B(n2779), .ZN(n2777)
         );
  OAI22_X1 U4609 ( .A1(n3655), .A2(n2336), .B1(n3252), .B2(n3481), .ZN(N410)
         );
  OAI22_X1 U4610 ( .A1(n3737), .A2(n3107), .B1(n3470), .B2(n3185), .ZN(N411)
         );
  OAI22_X1 U4611 ( .A1(n3645), .A2(n3033), .B1(n3334), .B2(n3622), .ZN(N412)
         );
  OAI22_X1 U4612 ( .A1(n3656), .A2(n3248), .B1(n3167), .B2(n3459), .ZN(N413)
         );
  OAI22_X1 U4613 ( .A1(n3665), .A2(n3183), .B1(n3420), .B2(n3622), .ZN(N414)
         );
  OAI22_X1 U4614 ( .A1(n3665), .A2(n2331), .B1(n3388), .B2(n3622), .ZN(N415)
         );
  OAI22_X1 U4615 ( .A1(n3772), .A2(n3067), .B1(n3315), .B2(n3755), .ZN(N521)
         );
  OAI22_X1 U4616 ( .A1(n3782), .A2(n3020), .B1(n3307), .B2(n2990), .ZN(N520)
         );
  OAI22_X1 U4617 ( .A1(n3427), .A2(n3103), .B1(n3188), .B2(n3753), .ZN(N519)
         );
  OAI22_X1 U4618 ( .A1(n3763), .A2(n3316), .B1(n3022), .B2(n2990), .ZN(N518)
         );
  OAI22_X1 U4619 ( .A1(n3762), .A2(n3233), .B1(n3114), .B2(n2989), .ZN(N517)
         );
  OAI22_X1 U4620 ( .A1(n3772), .A2(n3166), .B1(n3753), .B2(n3227), .ZN(N516)
         );
  OAI22_X1 U4621 ( .A1(n3783), .A2(n3222), .B1(n3163), .B2(n2990), .ZN(N515)
         );
  OAI22_X1 U4622 ( .A1(n3767), .A2(n3070), .B1(n3297), .B2(n3753), .ZN(N514)
         );
  OAI22_X1 U4623 ( .A1(n3773), .A2(n3105), .B1(n3181), .B2(n2990), .ZN(N513)
         );
  OAI22_X1 U4624 ( .A1(n3779), .A2(n3308), .B1(n3041), .B2(n2990), .ZN(N512)
         );
  OAI22_X1 U4625 ( .A1(n3764), .A2(n3243), .B1(n3158), .B2(n3753), .ZN(N511)
         );
  OAI22_X1 U4626 ( .A1(n3765), .A2(n3121), .B1(n3224), .B2(n3754), .ZN(N510)
         );
  OAI22_X1 U4627 ( .A1(n3764), .A2(n3122), .B1(n3176), .B2(n3752), .ZN(N498)
         );
  OAI22_X1 U4628 ( .A1(n3772), .A2(n3244), .B1(n3159), .B2(n3373), .ZN(N499)
         );
  OAI22_X1 U4629 ( .A1(n3768), .A2(n3309), .B1(n3042), .B2(n3754), .ZN(N500)
         );
  OAI22_X1 U4630 ( .A1(n3773), .A2(n3220), .B1(n3110), .B2(n3754), .ZN(N501)
         );
  OAI22_X1 U4631 ( .A1(n3429), .A2(n3104), .B1(n3180), .B2(n3372), .ZN(N502)
         );
  OAI22_X1 U4632 ( .A1(n3764), .A2(n3335), .B1(n3086), .B2(n3752), .ZN(N503)
         );
  OAI22_X1 U4633 ( .A1(n3772), .A2(n3066), .B1(n2989), .B2(n3317), .ZN(N497)
         );
  OAI22_X1 U4634 ( .A1(n3767), .A2(n3184), .B1(n3170), .B2(n3753), .ZN(N496)
         );
  OAI22_X1 U4635 ( .A1(n3768), .A2(n3059), .B1(n3303), .B2(n3753), .ZN(N495)
         );
  OAI22_X1 U4636 ( .A1(n3422), .A2(n3318), .B1(n3023), .B2(n3373), .ZN(N494)
         );
  OAI22_X1 U4637 ( .A1(n2985), .A2(n3234), .B1(n3115), .B2(n2989), .ZN(N493)
         );
  OAI22_X1 U4638 ( .A1(n3428), .A2(n3034), .B1(n3336), .B2(n2989), .ZN(N492)
         );
  OAI22_X1 U4639 ( .A1(n3767), .A2(n3111), .B1(n3253), .B2(n2989), .ZN(N491)
         );
  OAI22_X1 U4640 ( .A1(n3771), .A2(n3341), .B1(n3094), .B2(n3755), .ZN(N490)
         );
  OAI22_X1 U4641 ( .A1(n3771), .A2(n3012), .B1(n3260), .B2(n3755), .ZN(N489)
         );
  OAI22_X1 U4642 ( .A1(n3771), .A2(n3085), .B1(n3295), .B2(n3755), .ZN(N488)
         );
  OAI22_X1 U4643 ( .A1(n3770), .A2(n3223), .B1(n3112), .B2(n3755), .ZN(N487)
         );
  OAI22_X1 U4644 ( .A1(n2994), .A2(n3464), .B1(n3497), .B2(n2989), .ZN(N486)
         );
  AOI21_X1 U4645 ( .B1(n2674), .B2(n2240), .A(n2671), .ZN(n2665) );
  OAI22_X1 U4646 ( .A1(n3037), .A2(n3799), .B1(n3808), .B2(n3271), .ZN(N639)
         );
  OAI22_X1 U4647 ( .A1(n3134), .A2(n3797), .B1(n3821), .B2(n3219), .ZN(N638)
         );
  OAI22_X1 U4648 ( .A1(n3055), .A2(n3803), .B1(n3817), .B2(n3267), .ZN(N637)
         );
  OAI22_X1 U4649 ( .A1(n3273), .A2(n3803), .B1(n3817), .B2(n3060), .ZN(N636)
         );
  OAI22_X1 U4650 ( .A1(n3283), .A2(n3803), .B1(n3817), .B2(n3015), .ZN(N635)
         );
  OAI22_X1 U4651 ( .A1(n3089), .A2(n3803), .B1(n3818), .B2(n3179), .ZN(N634)
         );
  OAI22_X1 U4652 ( .A1(n3009), .A2(n3799), .B1(n3812), .B2(n3257), .ZN(N633)
         );
  OAI22_X1 U4653 ( .A1(n3126), .A2(n3796), .B1(n3609), .B2(n3214), .ZN(N632)
         );
  OAI22_X1 U4654 ( .A1(n3276), .A2(n3619), .B1(n3820), .B2(n3063), .ZN(N631)
         );
  OAI22_X1 U4655 ( .A1(n3119), .A2(n3797), .B1(n3818), .B2(n3208), .ZN(N630)
         );
  OAI22_X1 U4656 ( .A1(n3018), .A2(n3799), .B1(n3809), .B2(n3278), .ZN(N629)
         );
  OAI22_X1 U4657 ( .A1(n3796), .A2(n3249), .B1(n3828), .B2(n3148), .ZN(N628)
         );
  OAI211_X1 U4658 ( .C1(rC6[58]), .C2(n3237), .A(n2552), .B(n2405), .ZN(n2545)
         );
  AOI22_X1 U4659 ( .A1(n2605), .A2(n3495), .B1(n2606), .B2(n2607), .ZN(n2603)
         );
  INV_X1 U4660 ( .A(n2624), .ZN(n2474) );
  OAI221_X1 U4661 ( .B1(rC7[0]), .B2(n3683), .C1(rC7[1]), .C2(n3676), .A(n3496), .ZN(n2623) );
  OAI22_X1 U4662 ( .A1(n3344), .A2(n3798), .B1(n3468), .B2(n3025), .ZN(N627)
         );
  OAI22_X1 U4663 ( .A1(n3274), .A2(n3798), .B1(n3468), .B2(n3071), .ZN(N626)
         );
  OAI22_X1 U4664 ( .A1(n3054), .A2(n3798), .B1(n3828), .B2(n3266), .ZN(N625)
         );
  OAI22_X1 U4665 ( .A1(n3272), .A2(n3798), .B1(n3828), .B2(n3061), .ZN(N624)
         );
  OAI22_X1 U4666 ( .A1(n3279), .A2(n3798), .B1(n3810), .B2(n3016), .ZN(N623)
         );
  OAI22_X1 U4667 ( .A1(n3194), .A2(n3798), .B1(n3808), .B2(n3117), .ZN(N622)
         );
  OAI22_X1 U4668 ( .A1(n3092), .A2(n3798), .B1(n3617), .B2(n3285), .ZN(N621)
         );
  OAI22_X1 U4669 ( .A1(n3255), .A2(n3798), .B1(n3812), .B2(n3132), .ZN(N620)
         );
  OAI22_X1 U4670 ( .A1(n3193), .A2(n3798), .B1(n3609), .B2(n3099), .ZN(N619)
         );
  OAI22_X1 U4671 ( .A1(n3268), .A2(n3799), .B1(n3810), .B2(n3046), .ZN(N618)
         );
  OAI22_X1 U4672 ( .A1(n3217), .A2(n3460), .B1(n3818), .B2(n3127), .ZN(N617)
         );
  OAI22_X1 U4673 ( .A1(n3008), .A2(n3798), .B1(n3609), .B2(n3258), .ZN(N616)
         );
  OAI22_X1 U4674 ( .A1(n3784), .A2(n2260), .B1(n2992), .B2(n3463), .ZN(N485)
         );
  OAI22_X1 U4675 ( .A1(n3770), .A2(n3198), .B1(n3108), .B2(n2991), .ZN(N484)
         );
  OAI22_X1 U4676 ( .A1(n3772), .A2(n3498), .B1(n2992), .B2(n3478), .ZN(N483)
         );
  OAI22_X1 U4677 ( .A1(n3772), .A2(n2263), .B1(n2993), .B2(n3490), .ZN(N482)
         );
  OAI22_X1 U4678 ( .A1(n3772), .A2(n3241), .B1(n2991), .B2(n3142), .ZN(N481)
         );
  OAI22_X1 U4679 ( .A1(n3768), .A2(n3090), .B1(n3322), .B2(n2991), .ZN(N480)
         );
  OAI22_X1 U4680 ( .A1(n3769), .A2(n2266), .B1(n3310), .B2(n2992), .ZN(N479)
         );
  OAI22_X1 U4681 ( .A1(n2986), .A2(n3169), .B1(n3246), .B2(n2992), .ZN(N478)
         );
  OAI22_X1 U4682 ( .A1(n3422), .A2(n3201), .B1(n3109), .B2(n2993), .ZN(N477)
         );
  OAI22_X1 U4683 ( .A1(n2985), .A2(n3311), .B1(n2995), .B2(n3047), .ZN(N476)
         );
  OAI22_X1 U4684 ( .A1(n3784), .A2(n3236), .B1(n2993), .B2(n3152), .ZN(N475)
         );
  OAI22_X1 U4685 ( .A1(n3784), .A2(n3450), .B1(n2991), .B2(n3332), .ZN(N474)
         );
  OAI221_X1 U4686 ( .B1(n2641), .B2(n2642), .C1(rC2[63]), .C2(n3077), .A(n2643), .ZN(n2639) );
  OAI211_X1 U4687 ( .C1(n2615), .C2(n2616), .A(n2617), .B(n2618), .ZN(n2610)
         );
  OAI22_X1 U4688 ( .A1(n3685), .A2(n3619), .B1(n3817), .B2(n3679), .ZN(N604)
         );
  OAI22_X1 U4689 ( .A1(n3254), .A2(n3796), .B1(n3828), .B2(n3131), .ZN(N605)
         );
  OAI22_X1 U4690 ( .A1(n3800), .A2(n3687), .B1(n3817), .B2(n2999), .ZN(N603)
         );
  OAI22_X1 U4691 ( .A1(n3345), .A2(n3799), .B1(n3813), .B2(n3676), .ZN(N602)
         );
  OAI22_X1 U4692 ( .A1(n3192), .A2(n3804), .B1(n3609), .B2(n3116), .ZN(N600)
         );
  OAI22_X1 U4693 ( .A1(n3264), .A2(n3800), .B1(n3826), .B2(n3053), .ZN(N663)
         );
  OAI22_X1 U4694 ( .A1(n3038), .A2(n3800), .B1(n3808), .B2(n3343), .ZN(N598)
         );
  OAI22_X1 U4695 ( .A1(n3053), .A2(n3461), .B1(n3810), .B2(n3264), .ZN(N599)
         );
  OAI22_X1 U4696 ( .A1(n3203), .A2(n3804), .B1(n3815), .B2(n3147), .ZN(N596)
         );
  OAI22_X1 U4697 ( .A1(n3128), .A2(n3800), .B1(n3808), .B2(n3218), .ZN(N597)
         );
  OAI22_X1 U4698 ( .A1(n3024), .A2(n3800), .B1(n3818), .B2(n3275), .ZN(N594)
         );
  OAI22_X1 U4699 ( .A1(n3125), .A2(n3804), .B1(n3815), .B2(n3237), .ZN(N595)
         );
  OAI22_X1 U4700 ( .A1(n3213), .A2(n3800), .B1(n3813), .B2(n3133), .ZN(N592)
         );
  OAI22_X1 U4701 ( .A1(n3123), .A2(n3804), .B1(n3813), .B2(n3215), .ZN(N593)
         );
  OAI211_X1 U4702 ( .C1(n2571), .C2(n2572), .A(n2427), .B(n2573), .ZN(n2570)
         );
  OAI22_X1 U4703 ( .A1(n3280), .A2(n3801), .B1(n3810), .B2(n3026), .ZN(N590)
         );
  OAI22_X1 U4704 ( .A1(n3135), .A2(n3801), .B1(n3813), .B2(n3216), .ZN(N591)
         );
  OAI22_X1 U4705 ( .A1(n3160), .A2(n3801), .B1(n3812), .B2(n3250), .ZN(N588)
         );
  OAI22_X1 U4706 ( .A1(n3175), .A2(n3801), .B1(n3819), .B2(n3098), .ZN(N589)
         );
  OAI22_X1 U4707 ( .A1(n3173), .A2(n3801), .B1(n3819), .B2(n3096), .ZN(N586)
         );
  OAI22_X1 U4708 ( .A1(n3027), .A2(n3801), .B1(n3819), .B2(n3281), .ZN(N587)
         );
  OAI22_X1 U4709 ( .A1(n3035), .A2(n3801), .B1(n3609), .B2(n3269), .ZN(N584)
         );
  OAI22_X1 U4710 ( .A1(n3100), .A2(n3801), .B1(n3811), .B2(n3199), .ZN(N585)
         );
  OAI22_X1 U4711 ( .A1(n3161), .A2(n3801), .B1(n3817), .B2(n3251), .ZN(N582)
         );
  OAI22_X1 U4712 ( .A1(n3124), .A2(n3801), .B1(n3813), .B2(n3212), .ZN(N583)
         );
  OAI22_X1 U4713 ( .A1(n3801), .A2(n3039), .B1(n3826), .B2(n3282), .ZN(N581)
         );
  OAI22_X1 U4714 ( .A1(n3174), .A2(n3801), .B1(n3609), .B2(n3097), .ZN(N580)
         );
  OAI21_X1 U4715 ( .B1(n2585), .B2(n2586), .A(n3395), .ZN(n2579) );
  AOI221_X1 U4716 ( .B1(n3421), .B2(n2785), .C1(n2786), .C2(n2787), .A(n2788), 
        .ZN(n2781) );
  AOI221_X1 U4717 ( .B1(rC1[18]), .B2(n3013), .C1(n2781), .C2(n2780), .A(n2782), .ZN(n2779) );
  OAI222_X1 U4718 ( .A1(n2755), .A2(n2148), .B1(n2756), .B2(n2757), .C1(
        rC3[42]), .C2(n3078), .ZN(n2753) );
  AOI211_X1 U4719 ( .C1(rC1[43]), .C2(n3068), .A(n2754), .B(n2753), .ZN(n2752)
         );
  OAI22_X1 U4720 ( .A1(n2994), .A2(n3323), .B1(n3057), .B2(n3754), .ZN(N522)
         );
  AOI222_X1 U4721 ( .A1(rC2[42]), .A2(n3105), .B1(n2660), .B2(n2225), .C1(
        n2661), .C2(n2662), .ZN(n2655) );
  AOI221_X1 U4722 ( .B1(n2663), .B2(n2664), .C1(n2665), .C2(n2666), .A(n2667), 
        .ZN(n2660) );
  OAI22_X1 U4723 ( .A1(n3036), .A2(n3802), .B1(n3814), .B2(n3270), .ZN(N578)
         );
  OAI22_X1 U4724 ( .A1(n3101), .A2(n3802), .B1(n3811), .B2(n3200), .ZN(N579)
         );
  OAI22_X1 U4725 ( .A1(n3265), .A2(n3802), .B1(n3811), .B2(n3062), .ZN(N576)
         );
  OAI22_X1 U4726 ( .A1(n3129), .A2(n3454), .B1(n3809), .B2(n3205), .ZN(N577)
         );
  OAI22_X1 U4727 ( .A1(n3219), .A2(n3795), .B1(n3828), .B2(n3134), .ZN(N574)
         );
  OAI22_X1 U4728 ( .A1(n3271), .A2(n3802), .B1(n3609), .B2(n3037), .ZN(N575)
         );
  OAI22_X1 U4729 ( .A1(n3802), .A2(n3060), .B1(n3818), .B2(n3273), .ZN(N572)
         );
  OAI22_X1 U4730 ( .A1(n3267), .A2(n3802), .B1(n3814), .B2(n3055), .ZN(N573)
         );
  OAI22_X1 U4731 ( .A1(n3179), .A2(n3802), .B1(n3818), .B2(n3089), .ZN(N570)
         );
  OAI22_X1 U4732 ( .A1(n3015), .A2(n3802), .B1(n3810), .B2(n3283), .ZN(N571)
         );
  OAI22_X1 U4733 ( .A1(n3214), .A2(n3802), .B1(n3609), .B2(n3126), .ZN(N568)
         );
  OAI22_X1 U4734 ( .A1(n3257), .A2(n3802), .B1(n3818), .B2(n3009), .ZN(N569)
         );
  AOI211_X1 U4735 ( .C1(rC7[52]), .C2(n3175), .A(n2559), .B(n2558), .ZN(n2556)
         );
  OAI22_X1 U4736 ( .A1(n3132), .A2(n3803), .B1(n3818), .B2(n3255), .ZN(N556)
         );
  OAI211_X1 U4737 ( .C1(n2563), .C2(n2564), .A(n2420), .B(n2565), .ZN(n2562)
         );
  OAI221_X1 U4738 ( .B1(rC7[19]), .B2(n3132), .C1(n2596), .C2(n2597), .A(n2598), .ZN(n2595) );
  OAI22_X1 U4739 ( .A1(rC6[12]), .A2(n3684), .B1(rC6[11]), .B2(n3686), .ZN(
        n2626) );
  NOR3_X1 U4740 ( .A1(n2621), .A2(n2619), .A3(n2620), .ZN(n2618) );
  OAI21_X1 U4741 ( .B1(n2625), .B2(n3452), .A(n2606), .ZN(n2601) );
  INV_X2 U4742 ( .A(n3823), .ZN(n3797) );
  INV_X2 U4743 ( .A(n3822), .ZN(n3798) );
  INV_X2 U4744 ( .A(n3823), .ZN(n3799) );
  INV_X2 U4745 ( .A(n3832), .ZN(n3801) );
  INV_X2 U4746 ( .A(n3614), .ZN(n3802) );
  INV_X2 U4747 ( .A(n3823), .ZN(n3803) );
  INV_X1 U4748 ( .A(n3723), .ZN(n3691) );
  INV_X1 U4749 ( .A(n3786), .ZN(n3761) );
  INV_X1 U4750 ( .A(n3868), .ZN(n3836) );
endmodule

