
module GPR ( clk, reset, bus_in, inEn, outEn, bus_out );
  input [15:0] bus_in;
  output [15:0] bus_out;
  input clk, reset, inEn, outEn;
  wire   n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125;
  tri   \bus_out[15] ;
  tri   \bus_out[14] ;
  tri   \bus_out[13] ;
  tri   \bus_out[12] ;
  tri   \bus_out[11] ;
  tri   \bus_out[10] ;
  tri   \bus_out[9] ;
  tri   \bus_out[8] ;
  tri   \bus_out[7] ;
  tri   \bus_out[6] ;
  tri   \bus_out[5] ;
  tri   \bus_out[4] ;
  tri   \bus_out[3] ;
  tri   \bus_out[2] ;
  tri   \bus_out[1] ;
  tri   \bus_out[0] ;

  DFFARX2 \data_reg[14]  ( .D(n80), .CLK(clk), .RSTB(n98), .Q(n83) );
  DFFARX2 \data_reg[13]  ( .D(n79), .CLK(clk), .RSTB(n98), .Q(n84) );
  DFFARX2 \data_reg[9]  ( .D(n75), .CLK(clk), .RSTB(n98), .Q(n88) );
  DFFARX2 \data_reg[7]  ( .D(n73), .CLK(clk), .RSTB(n98), .Q(n90) );
  DFFARX2 \data_reg[6]  ( .D(n72), .CLK(clk), .RSTB(n98), .Q(n91) );
  DFFARX2 \data_reg[4]  ( .D(n70), .CLK(clk), .RSTB(n98), .Q(n93) );
  TNBUFFHX8 \bus_out_tri[0]  ( .IN(n125), .ENB(outEn), .Q(bus_out[0]) );
  TNBUFFHX8 \bus_out_tri[1]  ( .IN(n124), .ENB(outEn), .Q(bus_out[1]) );
  TNBUFFHX8 \bus_out_tri[2]  ( .IN(n123), .ENB(outEn), .Q(bus_out[2]) );
  TNBUFFHX8 \bus_out_tri[3]  ( .IN(n122), .ENB(outEn), .Q(bus_out[3]) );
  TNBUFFHX8 \bus_out_tri[4]  ( .IN(n121), .ENB(outEn), .Q(bus_out[4]) );
  TNBUFFHX8 \bus_out_tri[5]  ( .IN(n120), .ENB(outEn), .Q(bus_out[5]) );
  TNBUFFHX8 \bus_out_tri[6]  ( .IN(n119), .ENB(outEn), .Q(bus_out[6]) );
  TNBUFFHX8 \bus_out_tri[7]  ( .IN(n118), .ENB(outEn), .Q(bus_out[7]) );
  TNBUFFHX8 \bus_out_tri[8]  ( .IN(n117), .ENB(outEn), .Q(bus_out[8]) );
  TNBUFFHX8 \bus_out_tri[9]  ( .IN(n116), .ENB(outEn), .Q(bus_out[9]) );
  TNBUFFHX8 \bus_out_tri[10]  ( .IN(n115), .ENB(outEn), .Q(bus_out[10]) );
  TNBUFFHX8 \bus_out_tri[11]  ( .IN(n114), .ENB(outEn), .Q(bus_out[11]) );
  TNBUFFHX8 \bus_out_tri[12]  ( .IN(n113), .ENB(outEn), .Q(bus_out[12]) );
  TNBUFFHX8 \bus_out_tri[13]  ( .IN(n112), .ENB(outEn), .Q(bus_out[13]) );
  TNBUFFHX8 \bus_out_tri[14]  ( .IN(n111), .ENB(outEn), .Q(bus_out[14]) );
  TNBUFFHX8 \bus_out_tri[15]  ( .IN(n110), .ENB(outEn), .Q(bus_out[15]) );
  AO22X2 U38 ( .IN1(n110), .IN2(n99), .IN3(inEn), .IN4(bus_in[15]), .Q(n81) );
  AO22X2 U39 ( .IN1(n111), .IN2(n99), .IN3(bus_in[14]), .IN4(inEn), .Q(n80) );
  AO22X2 U40 ( .IN1(n112), .IN2(n99), .IN3(bus_in[13]), .IN4(inEn), .Q(n79) );
  AO22X2 U41 ( .IN1(n113), .IN2(n99), .IN3(bus_in[12]), .IN4(inEn), .Q(n78) );
  AO22X2 U42 ( .IN1(n114), .IN2(n99), .IN3(bus_in[11]), .IN4(inEn), .Q(n77) );
  AO22X2 U43 ( .IN1(n115), .IN2(n99), .IN3(bus_in[10]), .IN4(inEn), .Q(n76) );
  AO22X2 U44 ( .IN1(n116), .IN2(n99), .IN3(bus_in[9]), .IN4(inEn), .Q(n75) );
  AO22X2 U45 ( .IN1(n117), .IN2(n99), .IN3(bus_in[8]), .IN4(inEn), .Q(n74) );
  AO22X2 U46 ( .IN1(n118), .IN2(n99), .IN3(bus_in[7]), .IN4(inEn), .Q(n73) );
  AO22X2 U47 ( .IN1(n119), .IN2(n99), .IN3(bus_in[6]), .IN4(inEn), .Q(n72) );
  AO22X2 U48 ( .IN1(n120), .IN2(n99), .IN3(bus_in[5]), .IN4(inEn), .Q(n71) );
  AO22X2 U49 ( .IN1(n121), .IN2(n99), .IN3(bus_in[4]), .IN4(inEn), .Q(n70) );
  AO22X2 U50 ( .IN1(n122), .IN2(n99), .IN3(bus_in[3]), .IN4(inEn), .Q(n69) );
  AO22X2 U51 ( .IN1(n123), .IN2(n99), .IN3(bus_in[2]), .IN4(inEn), .Q(n68) );
  AO22X2 U52 ( .IN1(n124), .IN2(n99), .IN3(bus_in[1]), .IN4(inEn), .Q(n67) );
  AO22X2 U53 ( .IN1(n125), .IN2(n99), .IN3(bus_in[0]), .IN4(inEn), .Q(n66) );
  AODFFARX2 \data_reg[15]  ( .D(n81), .CLK(clk), .RSTB(n98), .Q(n82) );
  AODFFARX2 \data_reg[12]  ( .D(n78), .CLK(clk), .RSTB(n98), .Q(n85) );
  AODFFARX2 \data_reg[11]  ( .D(n77), .CLK(clk), .RSTB(n98), .Q(n86) );
  AODFFARX2 \data_reg[10]  ( .D(n76), .CLK(clk), .RSTB(n98), .Q(n87) );
  AODFFARX2 \data_reg[8]  ( .D(n74), .CLK(clk), .RSTB(n98), .Q(n89) );
  AODFFARX2 \data_reg[5]  ( .D(n71), .CLK(clk), .RSTB(n98), .Q(n92) );
  AODFFARX2 \data_reg[3]  ( .D(n69), .CLK(clk), .RSTB(n98), .Q(n94) );
  AODFFARX2 \data_reg[2]  ( .D(n68), .CLK(clk), .RSTB(n98), .Q(n95) );
  AODFFARX2 \data_reg[1]  ( .D(n67), .CLK(clk), .RSTB(n98), .Q(n96) );
  AODFFARX2 \data_reg[0]  ( .D(n66), .CLK(clk), .RSTB(n98), .Q(n97) );
  NBUFFX16 U54 ( .IN(n82), .Q(n110) );
  NBUFFX16 U55 ( .IN(n83), .Q(n111) );
  NBUFFX16 U56 ( .IN(n84), .Q(n112) );
  NBUFFX16 U57 ( .IN(n85), .Q(n113) );
  NBUFFX16 U58 ( .IN(n86), .Q(n114) );
  NBUFFX16 U59 ( .IN(n87), .Q(n115) );
  NBUFFX16 U60 ( .IN(n88), .Q(n116) );
  NBUFFX16 U61 ( .IN(n89), .Q(n117) );
  NBUFFX16 U62 ( .IN(n90), .Q(n118) );
  NBUFFX16 U63 ( .IN(n91), .Q(n119) );
  NBUFFX16 U64 ( .IN(n92), .Q(n120) );
  NBUFFX16 U65 ( .IN(n93), .Q(n121) );
  NBUFFX16 U66 ( .IN(n94), .Q(n122) );
  NBUFFX16 U67 ( .IN(n95), .Q(n123) );
  NBUFFX16 U68 ( .IN(n96), .Q(n124) );
  NBUFFX16 U69 ( .IN(n97), .Q(n125) );
  AOINVX2 U70 ( .IN(inEn), .QN(n99) );
  AOINVX2 U71 ( .IN(reset), .QN(n98) );
endmodule

