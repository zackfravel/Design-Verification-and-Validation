// Zack Fravel
// System Synthesis and Modeling
// Final Project (Step 4)

module moveImm_FSM(clk, reset, start, PCinc, 
		data_out, Ri1In, Ri2In, Ri3In, Ri4In, p1, p2, finish);

// Port Declartaion

input clk; input reset; input start; input[5:0] p1; input[5:0] p2; 

output reg PCinc; output[15:0] data_out; 
output reg Ri1In; output reg Ri2In; output reg Ri3In; output reg Ri4In; 
output reg finish;

reg[3:0] current_state, next_state;
reg dataTri;		

// Set Parameters for State Signals

parameter init = 4'b0000, one = 4'b0001, two = 4'b0010, three = 4'b0011, 
	four = 4'b0100, five = 4'b0101, six = 4'b0110, 	
	seven = 4'b0111, eight = 4'b1000, nine = 4'b1001, ten = 4'b1010;


// Architecture

always @(posedge clk or posedge reset)			// Current State Transition
begin
   if(reset)
	current_state <= init;
   else
	current_state <= next_state;
end


always @(current_state or start)			// Next State Logic
begin

   case(current_state)

   init: begin
	 	if(start)
	   		next_state <= one;
		else
			next_state <= init;
         end

   one:    begin next_state <= two; end
   two:    begin next_state <= three; end
   three:  begin next_state <= init; end
   default:begin next_state <= init; end

   endcase
end


always @(current_state)					// Output Logic
begin

   case (current_state)

   init:  begin 
		PCinc = 0; dataTri = 0; 
		Ri1In = 0; Ri2In = 0; Ri3In = 0; Ri4In = 0; 
		finish = 0;
	  end
   one:   begin  
		PCinc = 1; dataTri = 1;
		case (p1)
			6'b000001: begin Ri1In = 1; Ri2In = 0; Ri3In = 0; Ri4In = 0; end
			6'b000010: begin Ri2In = 1; Ri1In = 0; Ri3In = 0; Ri4In = 0; end
			6'b000011: begin Ri3In = 1; Ri2In = 0; Ri1In = 0; Ri4In = 0; end
			default  : begin Ri4In = 1; Ri2In = 0; Ri3In = 0; Ri1In = 0; end
		endcase 
	  end
   two:   begin 
		PCinc = 0; dataTri = 0; 
		case (p1)
			6'b000001: begin Ri1In = 0; Ri2In = 0; Ri3In = 0; Ri4In = 0; end
			6'b000010: begin Ri2In = 0; Ri1In = 0; Ri3In = 0; Ri4In = 0; end
			6'b000011: begin Ri3In = 0; Ri2In = 0; Ri1In = 0; Ri4In = 0; end
			default  : begin Ri4In = 0; Ri2In = 0; Ri3In = 0; Ri1In = 0; end
		endcase 
		finish = 1;
	  end
   three: begin 
		PCinc = 0; dataTri = 0; 
		Ri1In = 0; Ri2In = 0; Ri3In = 0; Ri4In = 0; 
		finish = 0;
	  end
   endcase

end

	assign data_out = (dataTri) ? p2:16'hzzzz;


endmodule
