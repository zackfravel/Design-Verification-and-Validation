
module myPMul32_4 ( g_inA0, g_inA1, g_inA2, g_inA3, g_inClk, g_outM );
  input [31:0] g_inA0;
  input [31:0] g_inA1;
  input [31:0] g_inA2;
  input [31:0] g_inA3;
  output [127:0] g_outM;
  input g_inClk;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15,
         N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29,
         N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43,
         N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57,
         N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71,
         N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85,
         N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99,
         N100, N101, N102, N103, N104, N105, N106, N107, N108, N109, N110,
         N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121,
         N122, N123, N124, N125, N126, N127, N128, N129, N130, N131, N132,
         N133, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143,
         N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154,
         N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165,
         N166, N167, N168, N169, N170, N171, N172, N173, N174, N175, N176,
         N177, N178, N179, N180, N181, N182, N183, N184, N185, N186, N187,
         N188, N189, N190, N191, N192, N193, N194, N195, N196, N197, N198,
         N199, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209,
         N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220,
         N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231,
         N232, N233, N234, N235, N236, N237, N238, N239, N240, N241, N242,
         N243, N244, N245, N246, N247, N248, N249, N250, N251, N252, N253,
         N254, N255, \mult_20/n63 , \mult_20/n62 , \mult_20/n61 ,
         \mult_20/n60 , \mult_20/n59 , \mult_20/n58 , \mult_20/n57 ,
         \mult_20/n56 , \mult_20/n55 , \mult_20/n54 , \mult_20/n53 ,
         \mult_20/n52 , \mult_20/n51 , \mult_20/n50 , \mult_20/n49 ,
         \mult_20/n48 , \mult_20/n47 , \mult_20/n46 , \mult_20/n45 ,
         \mult_20/n44 , \mult_20/n43 , \mult_20/n42 , \mult_20/n41 ,
         \mult_20/n40 , \mult_20/n39 , \mult_20/n38 , \mult_20/n37 ,
         \mult_20/n36 , \mult_20/n35 , \mult_20/n34 , \mult_20/n33 ,
         \mult_20/n32 , \mult_20/n31 , \mult_20/n30 , \mult_20/n29 ,
         \mult_20/n28 , \mult_20/n27 , \mult_20/n26 , \mult_20/n25 ,
         \mult_20/n24 , \mult_20/n23 , \mult_20/n22 , \mult_20/n21 ,
         \mult_20/n20 , \mult_20/n19 , \mult_20/n18 , \mult_20/n17 ,
         \mult_20/n16 , \mult_20/n15 , \mult_20/n14 , \mult_20/n13 ,
         \mult_20/n12 , \mult_20/n11 , \mult_20/n10 , \mult_20/n9 ,
         \mult_20/n8 , \mult_20/n7 , \mult_20/n6 , \mult_20/n5 , \mult_20/n4 ,
         \mult_20/n3 , \mult_20/SUMB[16][1] , \mult_20/SUMB[16][2] ,
         \mult_20/SUMB[16][3] , \mult_20/SUMB[16][4] , \mult_20/SUMB[16][5] ,
         \mult_20/SUMB[16][6] , \mult_20/SUMB[16][7] , \mult_20/SUMB[16][8] ,
         \mult_20/SUMB[16][9] , \mult_20/SUMB[16][10] , \mult_20/SUMB[16][11] ,
         \mult_20/SUMB[16][12] , \mult_20/SUMB[16][13] ,
         \mult_20/SUMB[16][14] , \mult_20/SUMB[16][15] ,
         \mult_20/SUMB[16][16] , \mult_20/SUMB[16][17] ,
         \mult_20/SUMB[16][18] , \mult_20/SUMB[16][19] ,
         \mult_20/SUMB[16][20] , \mult_20/SUMB[16][21] ,
         \mult_20/SUMB[16][22] , \mult_20/SUMB[16][23] ,
         \mult_20/SUMB[16][24] , \mult_20/SUMB[16][25] ,
         \mult_20/SUMB[16][26] , \mult_20/SUMB[16][27] ,
         \mult_20/SUMB[16][28] , \mult_20/SUMB[16][29] ,
         \mult_20/SUMB[16][30] , \mult_20/SUMB[17][1] , \mult_20/SUMB[17][2] ,
         \mult_20/SUMB[17][3] , \mult_20/SUMB[17][4] , \mult_20/SUMB[17][5] ,
         \mult_20/SUMB[17][6] , \mult_20/SUMB[17][7] , \mult_20/SUMB[17][8] ,
         \mult_20/SUMB[17][9] , \mult_20/SUMB[17][10] , \mult_20/SUMB[17][11] ,
         \mult_20/SUMB[17][12] , \mult_20/SUMB[17][13] ,
         \mult_20/SUMB[17][14] , \mult_20/SUMB[17][15] ,
         \mult_20/SUMB[17][16] , \mult_20/SUMB[17][17] ,
         \mult_20/SUMB[17][18] , \mult_20/SUMB[17][19] ,
         \mult_20/SUMB[17][20] , \mult_20/SUMB[17][21] ,
         \mult_20/SUMB[17][22] , \mult_20/SUMB[17][23] ,
         \mult_20/SUMB[17][24] , \mult_20/SUMB[17][25] ,
         \mult_20/SUMB[17][26] , \mult_20/SUMB[17][27] ,
         \mult_20/SUMB[17][28] , \mult_20/SUMB[17][29] ,
         \mult_20/SUMB[17][30] , \mult_20/SUMB[18][1] , \mult_20/SUMB[18][2] ,
         \mult_20/SUMB[18][3] , \mult_20/SUMB[18][4] , \mult_20/SUMB[18][5] ,
         \mult_20/SUMB[18][6] , \mult_20/SUMB[18][7] , \mult_20/SUMB[18][8] ,
         \mult_20/SUMB[18][9] , \mult_20/SUMB[18][10] , \mult_20/SUMB[18][11] ,
         \mult_20/SUMB[18][12] , \mult_20/SUMB[18][13] ,
         \mult_20/SUMB[18][14] , \mult_20/SUMB[18][15] ,
         \mult_20/SUMB[18][16] , \mult_20/SUMB[18][17] ,
         \mult_20/SUMB[18][18] , \mult_20/SUMB[18][19] ,
         \mult_20/SUMB[18][20] , \mult_20/SUMB[18][21] ,
         \mult_20/SUMB[18][22] , \mult_20/SUMB[18][23] ,
         \mult_20/SUMB[18][24] , \mult_20/SUMB[18][25] ,
         \mult_20/SUMB[18][26] , \mult_20/SUMB[18][27] ,
         \mult_20/SUMB[18][28] , \mult_20/SUMB[18][29] ,
         \mult_20/SUMB[18][30] , \mult_20/SUMB[19][1] , \mult_20/SUMB[19][2] ,
         \mult_20/SUMB[19][3] , \mult_20/SUMB[19][4] , \mult_20/SUMB[19][5] ,
         \mult_20/SUMB[19][6] , \mult_20/SUMB[19][7] , \mult_20/SUMB[19][8] ,
         \mult_20/SUMB[19][9] , \mult_20/SUMB[19][10] , \mult_20/SUMB[19][11] ,
         \mult_20/SUMB[19][12] , \mult_20/SUMB[19][13] ,
         \mult_20/SUMB[19][14] , \mult_20/SUMB[19][15] ,
         \mult_20/SUMB[19][16] , \mult_20/SUMB[19][17] ,
         \mult_20/SUMB[19][18] , \mult_20/SUMB[19][19] ,
         \mult_20/SUMB[19][20] , \mult_20/SUMB[19][21] ,
         \mult_20/SUMB[19][22] , \mult_20/SUMB[19][23] ,
         \mult_20/SUMB[19][24] , \mult_20/SUMB[19][25] ,
         \mult_20/SUMB[19][26] , \mult_20/SUMB[19][27] ,
         \mult_20/SUMB[19][28] , \mult_20/SUMB[19][29] ,
         \mult_20/SUMB[19][30] , \mult_20/SUMB[20][1] , \mult_20/SUMB[20][2] ,
         \mult_20/SUMB[20][3] , \mult_20/SUMB[20][4] , \mult_20/SUMB[20][5] ,
         \mult_20/SUMB[20][6] , \mult_20/SUMB[20][7] , \mult_20/SUMB[20][8] ,
         \mult_20/SUMB[20][9] , \mult_20/SUMB[20][10] , \mult_20/SUMB[20][11] ,
         \mult_20/SUMB[20][12] , \mult_20/SUMB[20][13] ,
         \mult_20/SUMB[20][14] , \mult_20/SUMB[20][15] ,
         \mult_20/SUMB[20][16] , \mult_20/SUMB[20][17] ,
         \mult_20/SUMB[20][18] , \mult_20/SUMB[20][19] ,
         \mult_20/SUMB[20][20] , \mult_20/SUMB[20][21] ,
         \mult_20/SUMB[20][22] , \mult_20/SUMB[20][23] ,
         \mult_20/SUMB[20][24] , \mult_20/SUMB[20][25] ,
         \mult_20/SUMB[20][26] , \mult_20/SUMB[20][27] ,
         \mult_20/SUMB[20][28] , \mult_20/SUMB[20][29] ,
         \mult_20/SUMB[20][30] , \mult_20/SUMB[21][1] , \mult_20/SUMB[21][2] ,
         \mult_20/SUMB[21][3] , \mult_20/SUMB[21][4] , \mult_20/SUMB[21][5] ,
         \mult_20/SUMB[21][6] , \mult_20/SUMB[21][7] , \mult_20/SUMB[21][8] ,
         \mult_20/SUMB[21][9] , \mult_20/SUMB[21][10] , \mult_20/SUMB[21][11] ,
         \mult_20/SUMB[21][12] , \mult_20/SUMB[21][13] ,
         \mult_20/SUMB[21][14] , \mult_20/SUMB[21][15] ,
         \mult_20/SUMB[21][16] , \mult_20/SUMB[21][17] ,
         \mult_20/SUMB[21][18] , \mult_20/SUMB[21][19] ,
         \mult_20/SUMB[21][20] , \mult_20/SUMB[21][21] ,
         \mult_20/SUMB[21][22] , \mult_20/SUMB[21][23] ,
         \mult_20/SUMB[21][24] , \mult_20/SUMB[21][25] ,
         \mult_20/SUMB[21][26] , \mult_20/SUMB[21][27] ,
         \mult_20/SUMB[21][28] , \mult_20/SUMB[21][29] ,
         \mult_20/SUMB[21][30] , \mult_20/SUMB[22][1] , \mult_20/SUMB[22][2] ,
         \mult_20/SUMB[22][3] , \mult_20/SUMB[22][4] , \mult_20/SUMB[22][5] ,
         \mult_20/SUMB[22][6] , \mult_20/SUMB[22][7] , \mult_20/SUMB[22][8] ,
         \mult_20/SUMB[22][9] , \mult_20/SUMB[22][10] , \mult_20/SUMB[22][11] ,
         \mult_20/SUMB[22][12] , \mult_20/SUMB[22][13] ,
         \mult_20/SUMB[22][14] , \mult_20/SUMB[22][15] ,
         \mult_20/SUMB[22][16] , \mult_20/SUMB[22][17] ,
         \mult_20/SUMB[22][18] , \mult_20/SUMB[22][19] ,
         \mult_20/SUMB[22][20] , \mult_20/SUMB[22][21] ,
         \mult_20/SUMB[22][22] , \mult_20/SUMB[22][23] ,
         \mult_20/SUMB[22][24] , \mult_20/SUMB[22][25] ,
         \mult_20/SUMB[22][26] , \mult_20/SUMB[22][27] ,
         \mult_20/SUMB[22][28] , \mult_20/SUMB[22][29] ,
         \mult_20/SUMB[22][30] , \mult_20/SUMB[23][1] , \mult_20/SUMB[23][2] ,
         \mult_20/SUMB[23][3] , \mult_20/SUMB[23][4] , \mult_20/SUMB[23][5] ,
         \mult_20/SUMB[23][6] , \mult_20/SUMB[23][7] , \mult_20/SUMB[23][8] ,
         \mult_20/SUMB[23][9] , \mult_20/SUMB[23][10] , \mult_20/SUMB[23][11] ,
         \mult_20/SUMB[23][12] , \mult_20/SUMB[23][13] ,
         \mult_20/SUMB[23][14] , \mult_20/SUMB[23][15] ,
         \mult_20/SUMB[23][16] , \mult_20/SUMB[23][17] ,
         \mult_20/SUMB[23][18] , \mult_20/SUMB[23][19] ,
         \mult_20/SUMB[23][20] , \mult_20/SUMB[23][21] ,
         \mult_20/SUMB[23][22] , \mult_20/SUMB[23][23] ,
         \mult_20/SUMB[23][24] , \mult_20/SUMB[23][25] ,
         \mult_20/SUMB[23][26] , \mult_20/SUMB[23][27] ,
         \mult_20/SUMB[23][28] , \mult_20/SUMB[23][29] ,
         \mult_20/SUMB[23][30] , \mult_20/SUMB[24][1] , \mult_20/SUMB[24][2] ,
         \mult_20/SUMB[24][3] , \mult_20/SUMB[24][4] , \mult_20/SUMB[24][5] ,
         \mult_20/SUMB[24][6] , \mult_20/SUMB[24][7] , \mult_20/SUMB[24][8] ,
         \mult_20/SUMB[24][9] , \mult_20/SUMB[24][10] , \mult_20/SUMB[24][11] ,
         \mult_20/SUMB[24][12] , \mult_20/SUMB[24][13] ,
         \mult_20/SUMB[24][14] , \mult_20/SUMB[24][15] ,
         \mult_20/SUMB[24][16] , \mult_20/SUMB[24][17] ,
         \mult_20/SUMB[24][18] , \mult_20/SUMB[24][19] ,
         \mult_20/SUMB[24][20] , \mult_20/SUMB[24][21] ,
         \mult_20/SUMB[24][22] , \mult_20/SUMB[24][23] ,
         \mult_20/SUMB[24][24] , \mult_20/SUMB[24][25] ,
         \mult_20/SUMB[24][26] , \mult_20/SUMB[24][27] ,
         \mult_20/SUMB[24][28] , \mult_20/SUMB[24][29] ,
         \mult_20/SUMB[24][30] , \mult_20/SUMB[25][1] , \mult_20/SUMB[25][2] ,
         \mult_20/SUMB[25][3] , \mult_20/SUMB[25][4] , \mult_20/SUMB[25][5] ,
         \mult_20/SUMB[25][6] , \mult_20/SUMB[25][7] , \mult_20/SUMB[25][8] ,
         \mult_20/SUMB[25][9] , \mult_20/SUMB[25][10] , \mult_20/SUMB[25][11] ,
         \mult_20/SUMB[25][12] , \mult_20/SUMB[25][13] ,
         \mult_20/SUMB[25][14] , \mult_20/SUMB[25][15] ,
         \mult_20/SUMB[25][16] , \mult_20/SUMB[25][17] ,
         \mult_20/SUMB[25][18] , \mult_20/SUMB[25][19] ,
         \mult_20/SUMB[25][20] , \mult_20/SUMB[25][21] ,
         \mult_20/SUMB[25][22] , \mult_20/SUMB[25][23] ,
         \mult_20/SUMB[25][24] , \mult_20/SUMB[25][25] ,
         \mult_20/SUMB[25][26] , \mult_20/SUMB[25][27] ,
         \mult_20/SUMB[25][28] , \mult_20/SUMB[25][29] ,
         \mult_20/SUMB[25][30] , \mult_20/SUMB[26][1] , \mult_20/SUMB[26][2] ,
         \mult_20/SUMB[26][3] , \mult_20/SUMB[26][4] , \mult_20/SUMB[26][5] ,
         \mult_20/SUMB[26][6] , \mult_20/SUMB[26][7] , \mult_20/SUMB[26][8] ,
         \mult_20/SUMB[26][9] , \mult_20/SUMB[26][10] , \mult_20/SUMB[26][11] ,
         \mult_20/SUMB[26][12] , \mult_20/SUMB[26][13] ,
         \mult_20/SUMB[26][14] , \mult_20/SUMB[26][15] ,
         \mult_20/SUMB[26][16] , \mult_20/SUMB[26][17] ,
         \mult_20/SUMB[26][18] , \mult_20/SUMB[26][19] ,
         \mult_20/SUMB[26][20] , \mult_20/SUMB[26][21] ,
         \mult_20/SUMB[26][22] , \mult_20/SUMB[26][23] ,
         \mult_20/SUMB[26][24] , \mult_20/SUMB[26][25] ,
         \mult_20/SUMB[26][26] , \mult_20/SUMB[26][27] ,
         \mult_20/SUMB[26][28] , \mult_20/SUMB[26][29] ,
         \mult_20/SUMB[26][30] , \mult_20/SUMB[27][1] , \mult_20/SUMB[27][2] ,
         \mult_20/SUMB[27][3] , \mult_20/SUMB[27][4] , \mult_20/SUMB[27][5] ,
         \mult_20/SUMB[27][6] , \mult_20/SUMB[27][7] , \mult_20/SUMB[27][8] ,
         \mult_20/SUMB[27][9] , \mult_20/SUMB[27][10] , \mult_20/SUMB[27][11] ,
         \mult_20/SUMB[27][12] , \mult_20/SUMB[27][13] ,
         \mult_20/SUMB[27][14] , \mult_20/SUMB[27][15] ,
         \mult_20/SUMB[27][16] , \mult_20/SUMB[27][17] ,
         \mult_20/SUMB[27][18] , \mult_20/SUMB[27][19] ,
         \mult_20/SUMB[27][20] , \mult_20/SUMB[27][21] ,
         \mult_20/SUMB[27][22] , \mult_20/SUMB[27][23] ,
         \mult_20/SUMB[27][24] , \mult_20/SUMB[27][25] ,
         \mult_20/SUMB[27][26] , \mult_20/SUMB[27][27] ,
         \mult_20/SUMB[27][28] , \mult_20/SUMB[27][29] ,
         \mult_20/SUMB[27][30] , \mult_20/SUMB[28][1] , \mult_20/SUMB[28][2] ,
         \mult_20/SUMB[28][3] , \mult_20/SUMB[28][4] , \mult_20/SUMB[28][5] ,
         \mult_20/SUMB[28][6] , \mult_20/SUMB[28][7] , \mult_20/SUMB[28][8] ,
         \mult_20/SUMB[28][9] , \mult_20/SUMB[28][10] , \mult_20/SUMB[28][11] ,
         \mult_20/SUMB[28][12] , \mult_20/SUMB[28][13] ,
         \mult_20/SUMB[28][14] , \mult_20/SUMB[28][15] ,
         \mult_20/SUMB[28][16] , \mult_20/SUMB[28][17] ,
         \mult_20/SUMB[28][18] , \mult_20/SUMB[28][19] ,
         \mult_20/SUMB[28][20] , \mult_20/SUMB[28][21] ,
         \mult_20/SUMB[28][22] , \mult_20/SUMB[28][23] ,
         \mult_20/SUMB[28][24] , \mult_20/SUMB[28][25] ,
         \mult_20/SUMB[28][26] , \mult_20/SUMB[28][27] ,
         \mult_20/SUMB[28][28] , \mult_20/SUMB[28][29] ,
         \mult_20/SUMB[28][30] , \mult_20/SUMB[29][1] , \mult_20/SUMB[29][2] ,
         \mult_20/SUMB[29][3] , \mult_20/SUMB[29][4] , \mult_20/SUMB[29][5] ,
         \mult_20/SUMB[29][6] , \mult_20/SUMB[29][7] , \mult_20/SUMB[29][8] ,
         \mult_20/SUMB[29][9] , \mult_20/SUMB[29][10] , \mult_20/SUMB[29][11] ,
         \mult_20/SUMB[29][12] , \mult_20/SUMB[29][13] ,
         \mult_20/SUMB[29][14] , \mult_20/SUMB[29][15] ,
         \mult_20/SUMB[29][16] , \mult_20/SUMB[29][17] ,
         \mult_20/SUMB[29][18] , \mult_20/SUMB[29][19] ,
         \mult_20/SUMB[29][20] , \mult_20/SUMB[29][21] ,
         \mult_20/SUMB[29][22] , \mult_20/SUMB[29][23] ,
         \mult_20/SUMB[29][24] , \mult_20/SUMB[29][25] ,
         \mult_20/SUMB[29][26] , \mult_20/SUMB[29][27] ,
         \mult_20/SUMB[29][28] , \mult_20/SUMB[29][29] ,
         \mult_20/SUMB[29][30] , \mult_20/SUMB[30][1] , \mult_20/SUMB[30][2] ,
         \mult_20/SUMB[30][3] , \mult_20/SUMB[30][4] , \mult_20/SUMB[30][5] ,
         \mult_20/SUMB[30][6] , \mult_20/SUMB[30][7] , \mult_20/SUMB[30][8] ,
         \mult_20/SUMB[30][9] , \mult_20/SUMB[30][10] , \mult_20/SUMB[30][11] ,
         \mult_20/SUMB[30][12] , \mult_20/SUMB[30][13] ,
         \mult_20/SUMB[30][14] , \mult_20/SUMB[30][15] ,
         \mult_20/SUMB[30][16] , \mult_20/SUMB[30][17] ,
         \mult_20/SUMB[30][18] , \mult_20/SUMB[30][19] ,
         \mult_20/SUMB[30][20] , \mult_20/SUMB[30][21] ,
         \mult_20/SUMB[30][22] , \mult_20/SUMB[30][23] ,
         \mult_20/SUMB[30][24] , \mult_20/SUMB[30][25] ,
         \mult_20/SUMB[30][26] , \mult_20/SUMB[30][27] ,
         \mult_20/SUMB[30][28] , \mult_20/SUMB[30][29] ,
         \mult_20/SUMB[30][30] , \mult_20/SUMB[31][1] , \mult_20/SUMB[31][2] ,
         \mult_20/SUMB[31][3] , \mult_20/SUMB[31][4] , \mult_20/SUMB[31][5] ,
         \mult_20/SUMB[31][6] , \mult_20/SUMB[31][7] , \mult_20/SUMB[31][8] ,
         \mult_20/SUMB[31][9] , \mult_20/SUMB[31][10] , \mult_20/SUMB[31][11] ,
         \mult_20/SUMB[31][12] , \mult_20/SUMB[31][13] ,
         \mult_20/SUMB[31][14] , \mult_20/SUMB[31][15] ,
         \mult_20/SUMB[31][16] , \mult_20/SUMB[31][17] ,
         \mult_20/SUMB[31][18] , \mult_20/SUMB[31][19] ,
         \mult_20/SUMB[31][20] , \mult_20/SUMB[31][21] ,
         \mult_20/SUMB[31][22] , \mult_20/SUMB[31][23] ,
         \mult_20/SUMB[31][24] , \mult_20/SUMB[31][25] ,
         \mult_20/SUMB[31][26] , \mult_20/SUMB[31][27] ,
         \mult_20/SUMB[31][28] , \mult_20/SUMB[31][29] ,
         \mult_20/SUMB[31][30] , \mult_20/CARRYB[16][0] ,
         \mult_20/CARRYB[16][1] , \mult_20/CARRYB[16][2] ,
         \mult_20/CARRYB[16][3] , \mult_20/CARRYB[16][4] ,
         \mult_20/CARRYB[16][5] , \mult_20/CARRYB[16][6] ,
         \mult_20/CARRYB[16][7] , \mult_20/CARRYB[16][8] ,
         \mult_20/CARRYB[16][9] , \mult_20/CARRYB[16][10] ,
         \mult_20/CARRYB[16][11] , \mult_20/CARRYB[16][12] ,
         \mult_20/CARRYB[16][13] , \mult_20/CARRYB[16][14] ,
         \mult_20/CARRYB[16][15] , \mult_20/CARRYB[16][16] ,
         \mult_20/CARRYB[16][17] , \mult_20/CARRYB[16][18] ,
         \mult_20/CARRYB[16][19] , \mult_20/CARRYB[16][20] ,
         \mult_20/CARRYB[16][21] , \mult_20/CARRYB[16][22] ,
         \mult_20/CARRYB[16][23] , \mult_20/CARRYB[16][24] ,
         \mult_20/CARRYB[16][25] , \mult_20/CARRYB[16][26] ,
         \mult_20/CARRYB[16][27] , \mult_20/CARRYB[16][28] ,
         \mult_20/CARRYB[16][29] , \mult_20/CARRYB[16][30] ,
         \mult_20/CARRYB[17][0] , \mult_20/CARRYB[17][1] ,
         \mult_20/CARRYB[17][2] , \mult_20/CARRYB[17][3] ,
         \mult_20/CARRYB[17][4] , \mult_20/CARRYB[17][5] ,
         \mult_20/CARRYB[17][6] , \mult_20/CARRYB[17][7] ,
         \mult_20/CARRYB[17][8] , \mult_20/CARRYB[17][9] ,
         \mult_20/CARRYB[17][10] , \mult_20/CARRYB[17][11] ,
         \mult_20/CARRYB[17][12] , \mult_20/CARRYB[17][13] ,
         \mult_20/CARRYB[17][14] , \mult_20/CARRYB[17][15] ,
         \mult_20/CARRYB[17][16] , \mult_20/CARRYB[17][17] ,
         \mult_20/CARRYB[17][18] , \mult_20/CARRYB[17][19] ,
         \mult_20/CARRYB[17][20] , \mult_20/CARRYB[17][21] ,
         \mult_20/CARRYB[17][22] , \mult_20/CARRYB[17][23] ,
         \mult_20/CARRYB[17][24] , \mult_20/CARRYB[17][25] ,
         \mult_20/CARRYB[17][26] , \mult_20/CARRYB[17][27] ,
         \mult_20/CARRYB[17][28] , \mult_20/CARRYB[17][29] ,
         \mult_20/CARRYB[17][30] , \mult_20/CARRYB[18][0] ,
         \mult_20/CARRYB[18][1] , \mult_20/CARRYB[18][2] ,
         \mult_20/CARRYB[18][3] , \mult_20/CARRYB[18][4] ,
         \mult_20/CARRYB[18][5] , \mult_20/CARRYB[18][6] ,
         \mult_20/CARRYB[18][7] , \mult_20/CARRYB[18][8] ,
         \mult_20/CARRYB[18][9] , \mult_20/CARRYB[18][10] ,
         \mult_20/CARRYB[18][11] , \mult_20/CARRYB[18][12] ,
         \mult_20/CARRYB[18][13] , \mult_20/CARRYB[18][14] ,
         \mult_20/CARRYB[18][15] , \mult_20/CARRYB[18][16] ,
         \mult_20/CARRYB[18][17] , \mult_20/CARRYB[18][18] ,
         \mult_20/CARRYB[18][19] , \mult_20/CARRYB[18][20] ,
         \mult_20/CARRYB[18][21] , \mult_20/CARRYB[18][22] ,
         \mult_20/CARRYB[18][23] , \mult_20/CARRYB[18][24] ,
         \mult_20/CARRYB[18][25] , \mult_20/CARRYB[18][26] ,
         \mult_20/CARRYB[18][27] , \mult_20/CARRYB[18][28] ,
         \mult_20/CARRYB[18][29] , \mult_20/CARRYB[18][30] ,
         \mult_20/CARRYB[19][0] , \mult_20/CARRYB[19][1] ,
         \mult_20/CARRYB[19][2] , \mult_20/CARRYB[19][3] ,
         \mult_20/CARRYB[19][4] , \mult_20/CARRYB[19][5] ,
         \mult_20/CARRYB[19][6] , \mult_20/CARRYB[19][7] ,
         \mult_20/CARRYB[19][8] , \mult_20/CARRYB[19][9] ,
         \mult_20/CARRYB[19][10] , \mult_20/CARRYB[19][11] ,
         \mult_20/CARRYB[19][12] , \mult_20/CARRYB[19][13] ,
         \mult_20/CARRYB[19][14] , \mult_20/CARRYB[19][15] ,
         \mult_20/CARRYB[19][16] , \mult_20/CARRYB[19][17] ,
         \mult_20/CARRYB[19][18] , \mult_20/CARRYB[19][19] ,
         \mult_20/CARRYB[19][20] , \mult_20/CARRYB[19][21] ,
         \mult_20/CARRYB[19][22] , \mult_20/CARRYB[19][23] ,
         \mult_20/CARRYB[19][24] , \mult_20/CARRYB[19][25] ,
         \mult_20/CARRYB[19][26] , \mult_20/CARRYB[19][27] ,
         \mult_20/CARRYB[19][28] , \mult_20/CARRYB[19][29] ,
         \mult_20/CARRYB[19][30] , \mult_20/CARRYB[20][0] ,
         \mult_20/CARRYB[20][1] , \mult_20/CARRYB[20][2] ,
         \mult_20/CARRYB[20][3] , \mult_20/CARRYB[20][4] ,
         \mult_20/CARRYB[20][5] , \mult_20/CARRYB[20][6] ,
         \mult_20/CARRYB[20][7] , \mult_20/CARRYB[20][8] ,
         \mult_20/CARRYB[20][9] , \mult_20/CARRYB[20][10] ,
         \mult_20/CARRYB[20][11] , \mult_20/CARRYB[20][12] ,
         \mult_20/CARRYB[20][13] , \mult_20/CARRYB[20][14] ,
         \mult_20/CARRYB[20][15] , \mult_20/CARRYB[20][16] ,
         \mult_20/CARRYB[20][17] , \mult_20/CARRYB[20][18] ,
         \mult_20/CARRYB[20][19] , \mult_20/CARRYB[20][20] ,
         \mult_20/CARRYB[20][21] , \mult_20/CARRYB[20][22] ,
         \mult_20/CARRYB[20][23] , \mult_20/CARRYB[20][24] ,
         \mult_20/CARRYB[20][25] , \mult_20/CARRYB[20][26] ,
         \mult_20/CARRYB[20][27] , \mult_20/CARRYB[20][28] ,
         \mult_20/CARRYB[20][29] , \mult_20/CARRYB[20][30] ,
         \mult_20/CARRYB[21][0] , \mult_20/CARRYB[21][1] ,
         \mult_20/CARRYB[21][2] , \mult_20/CARRYB[21][3] ,
         \mult_20/CARRYB[21][4] , \mult_20/CARRYB[21][5] ,
         \mult_20/CARRYB[21][6] , \mult_20/CARRYB[21][7] ,
         \mult_20/CARRYB[21][8] , \mult_20/CARRYB[21][9] ,
         \mult_20/CARRYB[21][10] , \mult_20/CARRYB[21][11] ,
         \mult_20/CARRYB[21][12] , \mult_20/CARRYB[21][13] ,
         \mult_20/CARRYB[21][14] , \mult_20/CARRYB[21][15] ,
         \mult_20/CARRYB[21][16] , \mult_20/CARRYB[21][17] ,
         \mult_20/CARRYB[21][18] , \mult_20/CARRYB[21][19] ,
         \mult_20/CARRYB[21][20] , \mult_20/CARRYB[21][21] ,
         \mult_20/CARRYB[21][22] , \mult_20/CARRYB[21][23] ,
         \mult_20/CARRYB[21][24] , \mult_20/CARRYB[21][25] ,
         \mult_20/CARRYB[21][26] , \mult_20/CARRYB[21][27] ,
         \mult_20/CARRYB[21][28] , \mult_20/CARRYB[21][29] ,
         \mult_20/CARRYB[21][30] , \mult_20/CARRYB[22][0] ,
         \mult_20/CARRYB[22][1] , \mult_20/CARRYB[22][2] ,
         \mult_20/CARRYB[22][3] , \mult_20/CARRYB[22][4] ,
         \mult_20/CARRYB[22][5] , \mult_20/CARRYB[22][6] ,
         \mult_20/CARRYB[22][7] , \mult_20/CARRYB[22][8] ,
         \mult_20/CARRYB[22][9] , \mult_20/CARRYB[22][10] ,
         \mult_20/CARRYB[22][11] , \mult_20/CARRYB[22][12] ,
         \mult_20/CARRYB[22][13] , \mult_20/CARRYB[22][14] ,
         \mult_20/CARRYB[22][15] , \mult_20/CARRYB[22][16] ,
         \mult_20/CARRYB[22][17] , \mult_20/CARRYB[22][18] ,
         \mult_20/CARRYB[22][19] , \mult_20/CARRYB[22][20] ,
         \mult_20/CARRYB[22][21] , \mult_20/CARRYB[22][22] ,
         \mult_20/CARRYB[22][23] , \mult_20/CARRYB[22][24] ,
         \mult_20/CARRYB[22][25] , \mult_20/CARRYB[22][26] ,
         \mult_20/CARRYB[22][27] , \mult_20/CARRYB[22][28] ,
         \mult_20/CARRYB[22][29] , \mult_20/CARRYB[22][30] ,
         \mult_20/CARRYB[23][0] , \mult_20/CARRYB[23][1] ,
         \mult_20/CARRYB[23][2] , \mult_20/CARRYB[23][3] ,
         \mult_20/CARRYB[23][4] , \mult_20/CARRYB[23][5] ,
         \mult_20/CARRYB[23][6] , \mult_20/CARRYB[23][7] ,
         \mult_20/CARRYB[23][8] , \mult_20/CARRYB[23][9] ,
         \mult_20/CARRYB[23][10] , \mult_20/CARRYB[23][11] ,
         \mult_20/CARRYB[23][12] , \mult_20/CARRYB[23][13] ,
         \mult_20/CARRYB[23][14] , \mult_20/CARRYB[23][15] ,
         \mult_20/CARRYB[23][16] , \mult_20/CARRYB[23][17] ,
         \mult_20/CARRYB[23][18] , \mult_20/CARRYB[23][19] ,
         \mult_20/CARRYB[23][20] , \mult_20/CARRYB[23][21] ,
         \mult_20/CARRYB[23][22] , \mult_20/CARRYB[23][23] ,
         \mult_20/CARRYB[23][24] , \mult_20/CARRYB[23][25] ,
         \mult_20/CARRYB[23][26] , \mult_20/CARRYB[23][27] ,
         \mult_20/CARRYB[23][28] , \mult_20/CARRYB[23][29] ,
         \mult_20/CARRYB[23][30] , \mult_20/CARRYB[24][0] ,
         \mult_20/CARRYB[24][1] , \mult_20/CARRYB[24][2] ,
         \mult_20/CARRYB[24][3] , \mult_20/CARRYB[24][4] ,
         \mult_20/CARRYB[24][5] , \mult_20/CARRYB[24][6] ,
         \mult_20/CARRYB[24][7] , \mult_20/CARRYB[24][8] ,
         \mult_20/CARRYB[24][9] , \mult_20/CARRYB[24][10] ,
         \mult_20/CARRYB[24][11] , \mult_20/CARRYB[24][12] ,
         \mult_20/CARRYB[24][13] , \mult_20/CARRYB[24][14] ,
         \mult_20/CARRYB[24][15] , \mult_20/CARRYB[24][16] ,
         \mult_20/CARRYB[24][17] , \mult_20/CARRYB[24][18] ,
         \mult_20/CARRYB[24][19] , \mult_20/CARRYB[24][20] ,
         \mult_20/CARRYB[24][21] , \mult_20/CARRYB[24][22] ,
         \mult_20/CARRYB[24][23] , \mult_20/CARRYB[24][24] ,
         \mult_20/CARRYB[24][25] , \mult_20/CARRYB[24][26] ,
         \mult_20/CARRYB[24][27] , \mult_20/CARRYB[24][28] ,
         \mult_20/CARRYB[24][29] , \mult_20/CARRYB[24][30] ,
         \mult_20/CARRYB[25][0] , \mult_20/CARRYB[25][1] ,
         \mult_20/CARRYB[25][2] , \mult_20/CARRYB[25][3] ,
         \mult_20/CARRYB[25][4] , \mult_20/CARRYB[25][5] ,
         \mult_20/CARRYB[25][6] , \mult_20/CARRYB[25][7] ,
         \mult_20/CARRYB[25][8] , \mult_20/CARRYB[25][9] ,
         \mult_20/CARRYB[25][10] , \mult_20/CARRYB[25][11] ,
         \mult_20/CARRYB[25][12] , \mult_20/CARRYB[25][13] ,
         \mult_20/CARRYB[25][14] , \mult_20/CARRYB[25][15] ,
         \mult_20/CARRYB[25][16] , \mult_20/CARRYB[25][17] ,
         \mult_20/CARRYB[25][18] , \mult_20/CARRYB[25][19] ,
         \mult_20/CARRYB[25][20] , \mult_20/CARRYB[25][21] ,
         \mult_20/CARRYB[25][22] , \mult_20/CARRYB[25][23] ,
         \mult_20/CARRYB[25][24] , \mult_20/CARRYB[25][25] ,
         \mult_20/CARRYB[25][26] , \mult_20/CARRYB[25][27] ,
         \mult_20/CARRYB[25][28] , \mult_20/CARRYB[25][29] ,
         \mult_20/CARRYB[25][30] , \mult_20/CARRYB[26][0] ,
         \mult_20/CARRYB[26][1] , \mult_20/CARRYB[26][2] ,
         \mult_20/CARRYB[26][3] , \mult_20/CARRYB[26][4] ,
         \mult_20/CARRYB[26][5] , \mult_20/CARRYB[26][6] ,
         \mult_20/CARRYB[26][7] , \mult_20/CARRYB[26][8] ,
         \mult_20/CARRYB[26][9] , \mult_20/CARRYB[26][10] ,
         \mult_20/CARRYB[26][11] , \mult_20/CARRYB[26][12] ,
         \mult_20/CARRYB[26][13] , \mult_20/CARRYB[26][14] ,
         \mult_20/CARRYB[26][15] , \mult_20/CARRYB[26][16] ,
         \mult_20/CARRYB[26][17] , \mult_20/CARRYB[26][18] ,
         \mult_20/CARRYB[26][19] , \mult_20/CARRYB[26][20] ,
         \mult_20/CARRYB[26][21] , \mult_20/CARRYB[26][22] ,
         \mult_20/CARRYB[26][23] , \mult_20/CARRYB[26][24] ,
         \mult_20/CARRYB[26][25] , \mult_20/CARRYB[26][26] ,
         \mult_20/CARRYB[26][27] , \mult_20/CARRYB[26][28] ,
         \mult_20/CARRYB[26][29] , \mult_20/CARRYB[26][30] ,
         \mult_20/CARRYB[27][0] , \mult_20/CARRYB[27][1] ,
         \mult_20/CARRYB[27][2] , \mult_20/CARRYB[27][3] ,
         \mult_20/CARRYB[27][4] , \mult_20/CARRYB[27][5] ,
         \mult_20/CARRYB[27][6] , \mult_20/CARRYB[27][7] ,
         \mult_20/CARRYB[27][8] , \mult_20/CARRYB[27][9] ,
         \mult_20/CARRYB[27][10] , \mult_20/CARRYB[27][11] ,
         \mult_20/CARRYB[27][12] , \mult_20/CARRYB[27][13] ,
         \mult_20/CARRYB[27][14] , \mult_20/CARRYB[27][15] ,
         \mult_20/CARRYB[27][16] , \mult_20/CARRYB[27][17] ,
         \mult_20/CARRYB[27][18] , \mult_20/CARRYB[27][19] ,
         \mult_20/CARRYB[27][20] , \mult_20/CARRYB[27][21] ,
         \mult_20/CARRYB[27][22] , \mult_20/CARRYB[27][23] ,
         \mult_20/CARRYB[27][24] , \mult_20/CARRYB[27][25] ,
         \mult_20/CARRYB[27][26] , \mult_20/CARRYB[27][27] ,
         \mult_20/CARRYB[27][28] , \mult_20/CARRYB[27][29] ,
         \mult_20/CARRYB[27][30] , \mult_20/CARRYB[28][0] ,
         \mult_20/CARRYB[28][1] , \mult_20/CARRYB[28][2] ,
         \mult_20/CARRYB[28][3] , \mult_20/CARRYB[28][4] ,
         \mult_20/CARRYB[28][5] , \mult_20/CARRYB[28][6] ,
         \mult_20/CARRYB[28][7] , \mult_20/CARRYB[28][8] ,
         \mult_20/CARRYB[28][9] , \mult_20/CARRYB[28][10] ,
         \mult_20/CARRYB[28][11] , \mult_20/CARRYB[28][12] ,
         \mult_20/CARRYB[28][13] , \mult_20/CARRYB[28][14] ,
         \mult_20/CARRYB[28][15] , \mult_20/CARRYB[28][16] ,
         \mult_20/CARRYB[28][17] , \mult_20/CARRYB[28][18] ,
         \mult_20/CARRYB[28][19] , \mult_20/CARRYB[28][20] ,
         \mult_20/CARRYB[28][21] , \mult_20/CARRYB[28][22] ,
         \mult_20/CARRYB[28][23] , \mult_20/CARRYB[28][24] ,
         \mult_20/CARRYB[28][25] , \mult_20/CARRYB[28][26] ,
         \mult_20/CARRYB[28][27] , \mult_20/CARRYB[28][28] ,
         \mult_20/CARRYB[28][29] , \mult_20/CARRYB[28][30] ,
         \mult_20/CARRYB[29][0] , \mult_20/CARRYB[29][1] ,
         \mult_20/CARRYB[29][2] , \mult_20/CARRYB[29][3] ,
         \mult_20/CARRYB[29][4] , \mult_20/CARRYB[29][5] ,
         \mult_20/CARRYB[29][6] , \mult_20/CARRYB[29][7] ,
         \mult_20/CARRYB[29][8] , \mult_20/CARRYB[29][9] ,
         \mult_20/CARRYB[29][10] , \mult_20/CARRYB[29][11] ,
         \mult_20/CARRYB[29][12] , \mult_20/CARRYB[29][13] ,
         \mult_20/CARRYB[29][14] , \mult_20/CARRYB[29][15] ,
         \mult_20/CARRYB[29][16] , \mult_20/CARRYB[29][17] ,
         \mult_20/CARRYB[29][18] , \mult_20/CARRYB[29][19] ,
         \mult_20/CARRYB[29][20] , \mult_20/CARRYB[29][21] ,
         \mult_20/CARRYB[29][22] , \mult_20/CARRYB[29][23] ,
         \mult_20/CARRYB[29][24] , \mult_20/CARRYB[29][25] ,
         \mult_20/CARRYB[29][26] , \mult_20/CARRYB[29][27] ,
         \mult_20/CARRYB[29][28] , \mult_20/CARRYB[29][29] ,
         \mult_20/CARRYB[29][30] , \mult_20/CARRYB[30][0] ,
         \mult_20/CARRYB[30][1] , \mult_20/CARRYB[30][2] ,
         \mult_20/CARRYB[30][3] , \mult_20/CARRYB[30][4] ,
         \mult_20/CARRYB[30][5] , \mult_20/CARRYB[30][6] ,
         \mult_20/CARRYB[30][7] , \mult_20/CARRYB[30][8] ,
         \mult_20/CARRYB[30][9] , \mult_20/CARRYB[30][10] ,
         \mult_20/CARRYB[30][11] , \mult_20/CARRYB[30][12] ,
         \mult_20/CARRYB[30][13] , \mult_20/CARRYB[30][14] ,
         \mult_20/CARRYB[30][15] , \mult_20/CARRYB[30][16] ,
         \mult_20/CARRYB[30][17] , \mult_20/CARRYB[30][18] ,
         \mult_20/CARRYB[30][19] , \mult_20/CARRYB[30][20] ,
         \mult_20/CARRYB[30][21] , \mult_20/CARRYB[30][22] ,
         \mult_20/CARRYB[30][23] , \mult_20/CARRYB[30][24] ,
         \mult_20/CARRYB[30][25] , \mult_20/CARRYB[30][26] ,
         \mult_20/CARRYB[30][27] , \mult_20/CARRYB[30][28] ,
         \mult_20/CARRYB[30][29] , \mult_20/CARRYB[30][30] ,
         \mult_20/CARRYB[31][0] , \mult_20/CARRYB[31][1] ,
         \mult_20/CARRYB[31][2] , \mult_20/CARRYB[31][3] ,
         \mult_20/CARRYB[31][4] , \mult_20/CARRYB[31][5] ,
         \mult_20/CARRYB[31][6] , \mult_20/CARRYB[31][7] ,
         \mult_20/CARRYB[31][8] , \mult_20/CARRYB[31][9] ,
         \mult_20/CARRYB[31][10] , \mult_20/CARRYB[31][11] ,
         \mult_20/CARRYB[31][12] , \mult_20/CARRYB[31][13] ,
         \mult_20/CARRYB[31][14] , \mult_20/CARRYB[31][15] ,
         \mult_20/CARRYB[31][16] , \mult_20/CARRYB[31][17] ,
         \mult_20/CARRYB[31][18] , \mult_20/CARRYB[31][19] ,
         \mult_20/CARRYB[31][20] , \mult_20/CARRYB[31][21] ,
         \mult_20/CARRYB[31][22] , \mult_20/CARRYB[31][23] ,
         \mult_20/CARRYB[31][24] , \mult_20/CARRYB[31][25] ,
         \mult_20/CARRYB[31][26] , \mult_20/CARRYB[31][27] ,
         \mult_20/CARRYB[31][28] , \mult_20/CARRYB[31][29] ,
         \mult_20/CARRYB[31][30] , \mult_20/SUMB[2][1] , \mult_20/SUMB[2][2] ,
         \mult_20/SUMB[2][3] , \mult_20/SUMB[2][4] , \mult_20/SUMB[2][5] ,
         \mult_20/SUMB[2][6] , \mult_20/SUMB[2][7] , \mult_20/SUMB[2][8] ,
         \mult_20/SUMB[2][9] , \mult_20/SUMB[2][10] , \mult_20/SUMB[2][11] ,
         \mult_20/SUMB[2][12] , \mult_20/SUMB[2][13] , \mult_20/SUMB[2][14] ,
         \mult_20/SUMB[2][15] , \mult_20/SUMB[2][16] , \mult_20/SUMB[2][17] ,
         \mult_20/SUMB[2][18] , \mult_20/SUMB[2][19] , \mult_20/SUMB[2][20] ,
         \mult_20/SUMB[2][21] , \mult_20/SUMB[2][22] , \mult_20/SUMB[2][23] ,
         \mult_20/SUMB[2][24] , \mult_20/SUMB[2][25] , \mult_20/SUMB[2][26] ,
         \mult_20/SUMB[2][27] , \mult_20/SUMB[2][28] , \mult_20/SUMB[2][29] ,
         \mult_20/SUMB[2][30] , \mult_20/SUMB[3][1] , \mult_20/SUMB[3][2] ,
         \mult_20/SUMB[3][3] , \mult_20/SUMB[3][4] , \mult_20/SUMB[3][5] ,
         \mult_20/SUMB[3][6] , \mult_20/SUMB[3][7] , \mult_20/SUMB[3][8] ,
         \mult_20/SUMB[3][9] , \mult_20/SUMB[3][10] , \mult_20/SUMB[3][11] ,
         \mult_20/SUMB[3][12] , \mult_20/SUMB[3][13] , \mult_20/SUMB[3][14] ,
         \mult_20/SUMB[3][15] , \mult_20/SUMB[3][16] , \mult_20/SUMB[3][17] ,
         \mult_20/SUMB[3][18] , \mult_20/SUMB[3][19] , \mult_20/SUMB[3][20] ,
         \mult_20/SUMB[3][21] , \mult_20/SUMB[3][22] , \mult_20/SUMB[3][23] ,
         \mult_20/SUMB[3][24] , \mult_20/SUMB[3][25] , \mult_20/SUMB[3][26] ,
         \mult_20/SUMB[3][27] , \mult_20/SUMB[3][28] , \mult_20/SUMB[3][29] ,
         \mult_20/SUMB[3][30] , \mult_20/SUMB[4][1] , \mult_20/SUMB[4][2] ,
         \mult_20/SUMB[4][3] , \mult_20/SUMB[4][4] , \mult_20/SUMB[4][5] ,
         \mult_20/SUMB[4][6] , \mult_20/SUMB[4][7] , \mult_20/SUMB[4][8] ,
         \mult_20/SUMB[4][9] , \mult_20/SUMB[4][10] , \mult_20/SUMB[4][11] ,
         \mult_20/SUMB[4][12] , \mult_20/SUMB[4][13] , \mult_20/SUMB[4][14] ,
         \mult_20/SUMB[4][15] , \mult_20/SUMB[4][16] , \mult_20/SUMB[4][17] ,
         \mult_20/SUMB[4][18] , \mult_20/SUMB[4][19] , \mult_20/SUMB[4][20] ,
         \mult_20/SUMB[4][21] , \mult_20/SUMB[4][22] , \mult_20/SUMB[4][23] ,
         \mult_20/SUMB[4][24] , \mult_20/SUMB[4][25] , \mult_20/SUMB[4][26] ,
         \mult_20/SUMB[4][27] , \mult_20/SUMB[4][28] , \mult_20/SUMB[4][29] ,
         \mult_20/SUMB[4][30] , \mult_20/SUMB[5][1] , \mult_20/SUMB[5][2] ,
         \mult_20/SUMB[5][3] , \mult_20/SUMB[5][4] , \mult_20/SUMB[5][5] ,
         \mult_20/SUMB[5][6] , \mult_20/SUMB[5][7] , \mult_20/SUMB[5][8] ,
         \mult_20/SUMB[5][9] , \mult_20/SUMB[5][10] , \mult_20/SUMB[5][11] ,
         \mult_20/SUMB[5][12] , \mult_20/SUMB[5][13] , \mult_20/SUMB[5][14] ,
         \mult_20/SUMB[5][15] , \mult_20/SUMB[5][16] , \mult_20/SUMB[5][17] ,
         \mult_20/SUMB[5][18] , \mult_20/SUMB[5][19] , \mult_20/SUMB[5][20] ,
         \mult_20/SUMB[5][21] , \mult_20/SUMB[5][22] , \mult_20/SUMB[5][23] ,
         \mult_20/SUMB[5][24] , \mult_20/SUMB[5][25] , \mult_20/SUMB[5][26] ,
         \mult_20/SUMB[5][27] , \mult_20/SUMB[5][28] , \mult_20/SUMB[5][29] ,
         \mult_20/SUMB[5][30] , \mult_20/SUMB[6][1] , \mult_20/SUMB[6][2] ,
         \mult_20/SUMB[6][3] , \mult_20/SUMB[6][4] , \mult_20/SUMB[6][5] ,
         \mult_20/SUMB[6][6] , \mult_20/SUMB[6][7] , \mult_20/SUMB[6][8] ,
         \mult_20/SUMB[6][9] , \mult_20/SUMB[6][10] , \mult_20/SUMB[6][11] ,
         \mult_20/SUMB[6][12] , \mult_20/SUMB[6][13] , \mult_20/SUMB[6][14] ,
         \mult_20/SUMB[6][15] , \mult_20/SUMB[6][16] , \mult_20/SUMB[6][17] ,
         \mult_20/SUMB[6][18] , \mult_20/SUMB[6][19] , \mult_20/SUMB[6][20] ,
         \mult_20/SUMB[6][21] , \mult_20/SUMB[6][22] , \mult_20/SUMB[6][23] ,
         \mult_20/SUMB[6][24] , \mult_20/SUMB[6][25] , \mult_20/SUMB[6][26] ,
         \mult_20/SUMB[6][27] , \mult_20/SUMB[6][28] , \mult_20/SUMB[6][29] ,
         \mult_20/SUMB[6][30] , \mult_20/SUMB[7][1] , \mult_20/SUMB[7][2] ,
         \mult_20/SUMB[7][3] , \mult_20/SUMB[7][4] , \mult_20/SUMB[7][5] ,
         \mult_20/SUMB[7][6] , \mult_20/SUMB[7][7] , \mult_20/SUMB[7][8] ,
         \mult_20/SUMB[7][9] , \mult_20/SUMB[7][10] , \mult_20/SUMB[7][11] ,
         \mult_20/SUMB[7][12] , \mult_20/SUMB[7][13] , \mult_20/SUMB[7][14] ,
         \mult_20/SUMB[7][15] , \mult_20/SUMB[7][16] , \mult_20/SUMB[7][17] ,
         \mult_20/SUMB[7][18] , \mult_20/SUMB[7][19] , \mult_20/SUMB[7][20] ,
         \mult_20/SUMB[7][21] , \mult_20/SUMB[7][22] , \mult_20/SUMB[7][23] ,
         \mult_20/SUMB[7][24] , \mult_20/SUMB[7][25] , \mult_20/SUMB[7][26] ,
         \mult_20/SUMB[7][27] , \mult_20/SUMB[7][28] , \mult_20/SUMB[7][29] ,
         \mult_20/SUMB[7][30] , \mult_20/SUMB[8][1] , \mult_20/SUMB[8][2] ,
         \mult_20/SUMB[8][3] , \mult_20/SUMB[8][4] , \mult_20/SUMB[8][5] ,
         \mult_20/SUMB[8][6] , \mult_20/SUMB[8][7] , \mult_20/SUMB[8][8] ,
         \mult_20/SUMB[8][9] , \mult_20/SUMB[8][10] , \mult_20/SUMB[8][11] ,
         \mult_20/SUMB[8][12] , \mult_20/SUMB[8][13] , \mult_20/SUMB[8][14] ,
         \mult_20/SUMB[8][15] , \mult_20/SUMB[8][16] , \mult_20/SUMB[8][17] ,
         \mult_20/SUMB[8][18] , \mult_20/SUMB[8][19] , \mult_20/SUMB[8][20] ,
         \mult_20/SUMB[8][21] , \mult_20/SUMB[8][22] , \mult_20/SUMB[8][23] ,
         \mult_20/SUMB[8][24] , \mult_20/SUMB[8][25] , \mult_20/SUMB[8][26] ,
         \mult_20/SUMB[8][27] , \mult_20/SUMB[8][28] , \mult_20/SUMB[8][29] ,
         \mult_20/SUMB[8][30] , \mult_20/SUMB[9][1] , \mult_20/SUMB[9][2] ,
         \mult_20/SUMB[9][3] , \mult_20/SUMB[9][4] , \mult_20/SUMB[9][5] ,
         \mult_20/SUMB[9][6] , \mult_20/SUMB[9][7] , \mult_20/SUMB[9][8] ,
         \mult_20/SUMB[9][9] , \mult_20/SUMB[9][10] , \mult_20/SUMB[9][11] ,
         \mult_20/SUMB[9][12] , \mult_20/SUMB[9][13] , \mult_20/SUMB[9][14] ,
         \mult_20/SUMB[9][15] , \mult_20/SUMB[9][16] , \mult_20/SUMB[9][17] ,
         \mult_20/SUMB[9][18] , \mult_20/SUMB[9][19] , \mult_20/SUMB[9][20] ,
         \mult_20/SUMB[9][21] , \mult_20/SUMB[9][22] , \mult_20/SUMB[9][23] ,
         \mult_20/SUMB[9][24] , \mult_20/SUMB[9][25] , \mult_20/SUMB[9][26] ,
         \mult_20/SUMB[9][27] , \mult_20/SUMB[9][28] , \mult_20/SUMB[9][29] ,
         \mult_20/SUMB[9][30] , \mult_20/SUMB[10][1] , \mult_20/SUMB[10][2] ,
         \mult_20/SUMB[10][3] , \mult_20/SUMB[10][4] , \mult_20/SUMB[10][5] ,
         \mult_20/SUMB[10][6] , \mult_20/SUMB[10][7] , \mult_20/SUMB[10][8] ,
         \mult_20/SUMB[10][9] , \mult_20/SUMB[10][10] , \mult_20/SUMB[10][11] ,
         \mult_20/SUMB[10][12] , \mult_20/SUMB[10][13] ,
         \mult_20/SUMB[10][14] , \mult_20/SUMB[10][15] ,
         \mult_20/SUMB[10][16] , \mult_20/SUMB[10][17] ,
         \mult_20/SUMB[10][18] , \mult_20/SUMB[10][19] ,
         \mult_20/SUMB[10][20] , \mult_20/SUMB[10][21] ,
         \mult_20/SUMB[10][22] , \mult_20/SUMB[10][23] ,
         \mult_20/SUMB[10][24] , \mult_20/SUMB[10][25] ,
         \mult_20/SUMB[10][26] , \mult_20/SUMB[10][27] ,
         \mult_20/SUMB[10][28] , \mult_20/SUMB[10][29] ,
         \mult_20/SUMB[10][30] , \mult_20/SUMB[11][1] , \mult_20/SUMB[11][2] ,
         \mult_20/SUMB[11][3] , \mult_20/SUMB[11][4] , \mult_20/SUMB[11][5] ,
         \mult_20/SUMB[11][6] , \mult_20/SUMB[11][7] , \mult_20/SUMB[11][8] ,
         \mult_20/SUMB[11][9] , \mult_20/SUMB[11][10] , \mult_20/SUMB[11][11] ,
         \mult_20/SUMB[11][12] , \mult_20/SUMB[11][13] ,
         \mult_20/SUMB[11][14] , \mult_20/SUMB[11][15] ,
         \mult_20/SUMB[11][16] , \mult_20/SUMB[11][17] ,
         \mult_20/SUMB[11][18] , \mult_20/SUMB[11][19] ,
         \mult_20/SUMB[11][20] , \mult_20/SUMB[11][21] ,
         \mult_20/SUMB[11][22] , \mult_20/SUMB[11][23] ,
         \mult_20/SUMB[11][24] , \mult_20/SUMB[11][25] ,
         \mult_20/SUMB[11][26] , \mult_20/SUMB[11][27] ,
         \mult_20/SUMB[11][28] , \mult_20/SUMB[11][29] ,
         \mult_20/SUMB[11][30] , \mult_20/SUMB[12][1] , \mult_20/SUMB[12][2] ,
         \mult_20/SUMB[12][3] , \mult_20/SUMB[12][4] , \mult_20/SUMB[12][5] ,
         \mult_20/SUMB[12][6] , \mult_20/SUMB[12][7] , \mult_20/SUMB[12][8] ,
         \mult_20/SUMB[12][9] , \mult_20/SUMB[12][10] , \mult_20/SUMB[12][11] ,
         \mult_20/SUMB[12][12] , \mult_20/SUMB[12][13] ,
         \mult_20/SUMB[12][14] , \mult_20/SUMB[12][15] ,
         \mult_20/SUMB[12][16] , \mult_20/SUMB[12][17] ,
         \mult_20/SUMB[12][18] , \mult_20/SUMB[12][19] ,
         \mult_20/SUMB[12][20] , \mult_20/SUMB[12][21] ,
         \mult_20/SUMB[12][22] , \mult_20/SUMB[12][23] ,
         \mult_20/SUMB[12][24] , \mult_20/SUMB[12][25] ,
         \mult_20/SUMB[12][26] , \mult_20/SUMB[12][27] ,
         \mult_20/SUMB[12][28] , \mult_20/SUMB[12][29] ,
         \mult_20/SUMB[12][30] , \mult_20/SUMB[13][1] , \mult_20/SUMB[13][2] ,
         \mult_20/SUMB[13][3] , \mult_20/SUMB[13][4] , \mult_20/SUMB[13][5] ,
         \mult_20/SUMB[13][6] , \mult_20/SUMB[13][7] , \mult_20/SUMB[13][8] ,
         \mult_20/SUMB[13][9] , \mult_20/SUMB[13][10] , \mult_20/SUMB[13][11] ,
         \mult_20/SUMB[13][12] , \mult_20/SUMB[13][13] ,
         \mult_20/SUMB[13][14] , \mult_20/SUMB[13][15] ,
         \mult_20/SUMB[13][16] , \mult_20/SUMB[13][17] ,
         \mult_20/SUMB[13][18] , \mult_20/SUMB[13][19] ,
         \mult_20/SUMB[13][20] , \mult_20/SUMB[13][21] ,
         \mult_20/SUMB[13][22] , \mult_20/SUMB[13][23] ,
         \mult_20/SUMB[13][24] , \mult_20/SUMB[13][25] ,
         \mult_20/SUMB[13][26] , \mult_20/SUMB[13][27] ,
         \mult_20/SUMB[13][28] , \mult_20/SUMB[13][29] ,
         \mult_20/SUMB[13][30] , \mult_20/SUMB[14][1] , \mult_20/SUMB[14][2] ,
         \mult_20/SUMB[14][3] , \mult_20/SUMB[14][4] , \mult_20/SUMB[14][5] ,
         \mult_20/SUMB[14][6] , \mult_20/SUMB[14][7] , \mult_20/SUMB[14][8] ,
         \mult_20/SUMB[14][9] , \mult_20/SUMB[14][10] , \mult_20/SUMB[14][11] ,
         \mult_20/SUMB[14][12] , \mult_20/SUMB[14][13] ,
         \mult_20/SUMB[14][14] , \mult_20/SUMB[14][15] ,
         \mult_20/SUMB[14][16] , \mult_20/SUMB[14][17] ,
         \mult_20/SUMB[14][18] , \mult_20/SUMB[14][19] ,
         \mult_20/SUMB[14][20] , \mult_20/SUMB[14][21] ,
         \mult_20/SUMB[14][22] , \mult_20/SUMB[14][23] ,
         \mult_20/SUMB[14][24] , \mult_20/SUMB[14][25] ,
         \mult_20/SUMB[14][26] , \mult_20/SUMB[14][27] ,
         \mult_20/SUMB[14][28] , \mult_20/SUMB[14][29] ,
         \mult_20/SUMB[14][30] , \mult_20/SUMB[15][1] , \mult_20/SUMB[15][2] ,
         \mult_20/SUMB[15][3] , \mult_20/SUMB[15][4] , \mult_20/SUMB[15][5] ,
         \mult_20/SUMB[15][6] , \mult_20/SUMB[15][7] , \mult_20/SUMB[15][8] ,
         \mult_20/SUMB[15][9] , \mult_20/SUMB[15][10] , \mult_20/SUMB[15][11] ,
         \mult_20/SUMB[15][12] , \mult_20/SUMB[15][13] ,
         \mult_20/SUMB[15][14] , \mult_20/SUMB[15][15] ,
         \mult_20/SUMB[15][16] , \mult_20/SUMB[15][17] ,
         \mult_20/SUMB[15][18] , \mult_20/SUMB[15][19] ,
         \mult_20/SUMB[15][20] , \mult_20/SUMB[15][21] ,
         \mult_20/SUMB[15][22] , \mult_20/SUMB[15][23] ,
         \mult_20/SUMB[15][24] , \mult_20/SUMB[15][25] ,
         \mult_20/SUMB[15][26] , \mult_20/SUMB[15][27] ,
         \mult_20/SUMB[15][28] , \mult_20/SUMB[15][29] ,
         \mult_20/SUMB[15][30] , \mult_20/CARRYB[2][0] ,
         \mult_20/CARRYB[2][1] , \mult_20/CARRYB[2][2] ,
         \mult_20/CARRYB[2][3] , \mult_20/CARRYB[2][4] ,
         \mult_20/CARRYB[2][5] , \mult_20/CARRYB[2][6] ,
         \mult_20/CARRYB[2][7] , \mult_20/CARRYB[2][8] ,
         \mult_20/CARRYB[2][9] , \mult_20/CARRYB[2][10] ,
         \mult_20/CARRYB[2][11] , \mult_20/CARRYB[2][12] ,
         \mult_20/CARRYB[2][13] , \mult_20/CARRYB[2][14] ,
         \mult_20/CARRYB[2][15] , \mult_20/CARRYB[2][16] ,
         \mult_20/CARRYB[2][17] , \mult_20/CARRYB[2][18] ,
         \mult_20/CARRYB[2][19] , \mult_20/CARRYB[2][20] ,
         \mult_20/CARRYB[2][21] , \mult_20/CARRYB[2][22] ,
         \mult_20/CARRYB[2][23] , \mult_20/CARRYB[2][24] ,
         \mult_20/CARRYB[2][25] , \mult_20/CARRYB[2][26] ,
         \mult_20/CARRYB[2][27] , \mult_20/CARRYB[2][28] ,
         \mult_20/CARRYB[2][29] , \mult_20/CARRYB[2][30] ,
         \mult_20/CARRYB[3][0] , \mult_20/CARRYB[3][1] ,
         \mult_20/CARRYB[3][2] , \mult_20/CARRYB[3][3] ,
         \mult_20/CARRYB[3][4] , \mult_20/CARRYB[3][5] ,
         \mult_20/CARRYB[3][6] , \mult_20/CARRYB[3][7] ,
         \mult_20/CARRYB[3][8] , \mult_20/CARRYB[3][9] ,
         \mult_20/CARRYB[3][10] , \mult_20/CARRYB[3][11] ,
         \mult_20/CARRYB[3][12] , \mult_20/CARRYB[3][13] ,
         \mult_20/CARRYB[3][14] , \mult_20/CARRYB[3][15] ,
         \mult_20/CARRYB[3][16] , \mult_20/CARRYB[3][17] ,
         \mult_20/CARRYB[3][18] , \mult_20/CARRYB[3][19] ,
         \mult_20/CARRYB[3][20] , \mult_20/CARRYB[3][21] ,
         \mult_20/CARRYB[3][22] , \mult_20/CARRYB[3][23] ,
         \mult_20/CARRYB[3][24] , \mult_20/CARRYB[3][25] ,
         \mult_20/CARRYB[3][26] , \mult_20/CARRYB[3][27] ,
         \mult_20/CARRYB[3][28] , \mult_20/CARRYB[3][29] ,
         \mult_20/CARRYB[3][30] , \mult_20/CARRYB[4][0] ,
         \mult_20/CARRYB[4][1] , \mult_20/CARRYB[4][2] ,
         \mult_20/CARRYB[4][3] , \mult_20/CARRYB[4][4] ,
         \mult_20/CARRYB[4][5] , \mult_20/CARRYB[4][6] ,
         \mult_20/CARRYB[4][7] , \mult_20/CARRYB[4][8] ,
         \mult_20/CARRYB[4][9] , \mult_20/CARRYB[4][10] ,
         \mult_20/CARRYB[4][11] , \mult_20/CARRYB[4][12] ,
         \mult_20/CARRYB[4][13] , \mult_20/CARRYB[4][14] ,
         \mult_20/CARRYB[4][15] , \mult_20/CARRYB[4][16] ,
         \mult_20/CARRYB[4][17] , \mult_20/CARRYB[4][18] ,
         \mult_20/CARRYB[4][19] , \mult_20/CARRYB[4][20] ,
         \mult_20/CARRYB[4][21] , \mult_20/CARRYB[4][22] ,
         \mult_20/CARRYB[4][23] , \mult_20/CARRYB[4][24] ,
         \mult_20/CARRYB[4][25] , \mult_20/CARRYB[4][26] ,
         \mult_20/CARRYB[4][27] , \mult_20/CARRYB[4][28] ,
         \mult_20/CARRYB[4][29] , \mult_20/CARRYB[4][30] ,
         \mult_20/CARRYB[5][0] , \mult_20/CARRYB[5][1] ,
         \mult_20/CARRYB[5][2] , \mult_20/CARRYB[5][3] ,
         \mult_20/CARRYB[5][4] , \mult_20/CARRYB[5][5] ,
         \mult_20/CARRYB[5][6] , \mult_20/CARRYB[5][7] ,
         \mult_20/CARRYB[5][8] , \mult_20/CARRYB[5][9] ,
         \mult_20/CARRYB[5][10] , \mult_20/CARRYB[5][11] ,
         \mult_20/CARRYB[5][12] , \mult_20/CARRYB[5][13] ,
         \mult_20/CARRYB[5][14] , \mult_20/CARRYB[5][15] ,
         \mult_20/CARRYB[5][16] , \mult_20/CARRYB[5][17] ,
         \mult_20/CARRYB[5][18] , \mult_20/CARRYB[5][19] ,
         \mult_20/CARRYB[5][20] , \mult_20/CARRYB[5][21] ,
         \mult_20/CARRYB[5][22] , \mult_20/CARRYB[5][23] ,
         \mult_20/CARRYB[5][24] , \mult_20/CARRYB[5][25] ,
         \mult_20/CARRYB[5][26] , \mult_20/CARRYB[5][27] ,
         \mult_20/CARRYB[5][28] , \mult_20/CARRYB[5][29] ,
         \mult_20/CARRYB[5][30] , \mult_20/CARRYB[6][0] ,
         \mult_20/CARRYB[6][1] , \mult_20/CARRYB[6][2] ,
         \mult_20/CARRYB[6][3] , \mult_20/CARRYB[6][4] ,
         \mult_20/CARRYB[6][5] , \mult_20/CARRYB[6][6] ,
         \mult_20/CARRYB[6][7] , \mult_20/CARRYB[6][8] ,
         \mult_20/CARRYB[6][9] , \mult_20/CARRYB[6][10] ,
         \mult_20/CARRYB[6][11] , \mult_20/CARRYB[6][12] ,
         \mult_20/CARRYB[6][13] , \mult_20/CARRYB[6][14] ,
         \mult_20/CARRYB[6][15] , \mult_20/CARRYB[6][16] ,
         \mult_20/CARRYB[6][17] , \mult_20/CARRYB[6][18] ,
         \mult_20/CARRYB[6][19] , \mult_20/CARRYB[6][20] ,
         \mult_20/CARRYB[6][21] , \mult_20/CARRYB[6][22] ,
         \mult_20/CARRYB[6][23] , \mult_20/CARRYB[6][24] ,
         \mult_20/CARRYB[6][25] , \mult_20/CARRYB[6][26] ,
         \mult_20/CARRYB[6][27] , \mult_20/CARRYB[6][28] ,
         \mult_20/CARRYB[6][29] , \mult_20/CARRYB[6][30] ,
         \mult_20/CARRYB[7][0] , \mult_20/CARRYB[7][1] ,
         \mult_20/CARRYB[7][2] , \mult_20/CARRYB[7][3] ,
         \mult_20/CARRYB[7][4] , \mult_20/CARRYB[7][5] ,
         \mult_20/CARRYB[7][6] , \mult_20/CARRYB[7][7] ,
         \mult_20/CARRYB[7][8] , \mult_20/CARRYB[7][9] ,
         \mult_20/CARRYB[7][10] , \mult_20/CARRYB[7][11] ,
         \mult_20/CARRYB[7][12] , \mult_20/CARRYB[7][13] ,
         \mult_20/CARRYB[7][14] , \mult_20/CARRYB[7][15] ,
         \mult_20/CARRYB[7][16] , \mult_20/CARRYB[7][17] ,
         \mult_20/CARRYB[7][18] , \mult_20/CARRYB[7][19] ,
         \mult_20/CARRYB[7][20] , \mult_20/CARRYB[7][21] ,
         \mult_20/CARRYB[7][22] , \mult_20/CARRYB[7][23] ,
         \mult_20/CARRYB[7][24] , \mult_20/CARRYB[7][25] ,
         \mult_20/CARRYB[7][26] , \mult_20/CARRYB[7][27] ,
         \mult_20/CARRYB[7][28] , \mult_20/CARRYB[7][29] ,
         \mult_20/CARRYB[7][30] , \mult_20/CARRYB[8][0] ,
         \mult_20/CARRYB[8][1] , \mult_20/CARRYB[8][2] ,
         \mult_20/CARRYB[8][3] , \mult_20/CARRYB[8][4] ,
         \mult_20/CARRYB[8][5] , \mult_20/CARRYB[8][6] ,
         \mult_20/CARRYB[8][7] , \mult_20/CARRYB[8][8] ,
         \mult_20/CARRYB[8][9] , \mult_20/CARRYB[8][10] ,
         \mult_20/CARRYB[8][11] , \mult_20/CARRYB[8][12] ,
         \mult_20/CARRYB[8][13] , \mult_20/CARRYB[8][14] ,
         \mult_20/CARRYB[8][15] , \mult_20/CARRYB[8][16] ,
         \mult_20/CARRYB[8][17] , \mult_20/CARRYB[8][18] ,
         \mult_20/CARRYB[8][19] , \mult_20/CARRYB[8][20] ,
         \mult_20/CARRYB[8][21] , \mult_20/CARRYB[8][22] ,
         \mult_20/CARRYB[8][23] , \mult_20/CARRYB[8][24] ,
         \mult_20/CARRYB[8][25] , \mult_20/CARRYB[8][26] ,
         \mult_20/CARRYB[8][27] , \mult_20/CARRYB[8][28] ,
         \mult_20/CARRYB[8][29] , \mult_20/CARRYB[8][30] ,
         \mult_20/CARRYB[9][0] , \mult_20/CARRYB[9][1] ,
         \mult_20/CARRYB[9][2] , \mult_20/CARRYB[9][3] ,
         \mult_20/CARRYB[9][4] , \mult_20/CARRYB[9][5] ,
         \mult_20/CARRYB[9][6] , \mult_20/CARRYB[9][7] ,
         \mult_20/CARRYB[9][8] , \mult_20/CARRYB[9][9] ,
         \mult_20/CARRYB[9][10] , \mult_20/CARRYB[9][11] ,
         \mult_20/CARRYB[9][12] , \mult_20/CARRYB[9][13] ,
         \mult_20/CARRYB[9][14] , \mult_20/CARRYB[9][15] ,
         \mult_20/CARRYB[9][16] , \mult_20/CARRYB[9][17] ,
         \mult_20/CARRYB[9][18] , \mult_20/CARRYB[9][19] ,
         \mult_20/CARRYB[9][20] , \mult_20/CARRYB[9][21] ,
         \mult_20/CARRYB[9][22] , \mult_20/CARRYB[9][23] ,
         \mult_20/CARRYB[9][24] , \mult_20/CARRYB[9][25] ,
         \mult_20/CARRYB[9][26] , \mult_20/CARRYB[9][27] ,
         \mult_20/CARRYB[9][28] , \mult_20/CARRYB[9][29] ,
         \mult_20/CARRYB[9][30] , \mult_20/CARRYB[10][0] ,
         \mult_20/CARRYB[10][1] , \mult_20/CARRYB[10][2] ,
         \mult_20/CARRYB[10][3] , \mult_20/CARRYB[10][4] ,
         \mult_20/CARRYB[10][5] , \mult_20/CARRYB[10][6] ,
         \mult_20/CARRYB[10][7] , \mult_20/CARRYB[10][8] ,
         \mult_20/CARRYB[10][9] , \mult_20/CARRYB[10][10] ,
         \mult_20/CARRYB[10][11] , \mult_20/CARRYB[10][12] ,
         \mult_20/CARRYB[10][13] , \mult_20/CARRYB[10][14] ,
         \mult_20/CARRYB[10][15] , \mult_20/CARRYB[10][16] ,
         \mult_20/CARRYB[10][17] , \mult_20/CARRYB[10][18] ,
         \mult_20/CARRYB[10][19] , \mult_20/CARRYB[10][20] ,
         \mult_20/CARRYB[10][21] , \mult_20/CARRYB[10][22] ,
         \mult_20/CARRYB[10][23] , \mult_20/CARRYB[10][24] ,
         \mult_20/CARRYB[10][25] , \mult_20/CARRYB[10][26] ,
         \mult_20/CARRYB[10][27] , \mult_20/CARRYB[10][28] ,
         \mult_20/CARRYB[10][29] , \mult_20/CARRYB[10][30] ,
         \mult_20/CARRYB[11][0] , \mult_20/CARRYB[11][1] ,
         \mult_20/CARRYB[11][2] , \mult_20/CARRYB[11][3] ,
         \mult_20/CARRYB[11][4] , \mult_20/CARRYB[11][5] ,
         \mult_20/CARRYB[11][6] , \mult_20/CARRYB[11][7] ,
         \mult_20/CARRYB[11][8] , \mult_20/CARRYB[11][9] ,
         \mult_20/CARRYB[11][10] , \mult_20/CARRYB[11][11] ,
         \mult_20/CARRYB[11][12] , \mult_20/CARRYB[11][13] ,
         \mult_20/CARRYB[11][14] , \mult_20/CARRYB[11][15] ,
         \mult_20/CARRYB[11][16] , \mult_20/CARRYB[11][17] ,
         \mult_20/CARRYB[11][18] , \mult_20/CARRYB[11][19] ,
         \mult_20/CARRYB[11][20] , \mult_20/CARRYB[11][21] ,
         \mult_20/CARRYB[11][22] , \mult_20/CARRYB[11][23] ,
         \mult_20/CARRYB[11][24] , \mult_20/CARRYB[11][25] ,
         \mult_20/CARRYB[11][26] , \mult_20/CARRYB[11][27] ,
         \mult_20/CARRYB[11][28] , \mult_20/CARRYB[11][29] ,
         \mult_20/CARRYB[11][30] , \mult_20/CARRYB[12][0] ,
         \mult_20/CARRYB[12][1] , \mult_20/CARRYB[12][2] ,
         \mult_20/CARRYB[12][3] , \mult_20/CARRYB[12][4] ,
         \mult_20/CARRYB[12][5] , \mult_20/CARRYB[12][6] ,
         \mult_20/CARRYB[12][7] , \mult_20/CARRYB[12][8] ,
         \mult_20/CARRYB[12][9] , \mult_20/CARRYB[12][10] ,
         \mult_20/CARRYB[12][11] , \mult_20/CARRYB[12][12] ,
         \mult_20/CARRYB[12][13] , \mult_20/CARRYB[12][14] ,
         \mult_20/CARRYB[12][15] , \mult_20/CARRYB[12][16] ,
         \mult_20/CARRYB[12][17] , \mult_20/CARRYB[12][18] ,
         \mult_20/CARRYB[12][19] , \mult_20/CARRYB[12][20] ,
         \mult_20/CARRYB[12][21] , \mult_20/CARRYB[12][22] ,
         \mult_20/CARRYB[12][23] , \mult_20/CARRYB[12][24] ,
         \mult_20/CARRYB[12][25] , \mult_20/CARRYB[12][26] ,
         \mult_20/CARRYB[12][27] , \mult_20/CARRYB[12][28] ,
         \mult_20/CARRYB[12][29] , \mult_20/CARRYB[12][30] ,
         \mult_20/CARRYB[13][0] , \mult_20/CARRYB[13][1] ,
         \mult_20/CARRYB[13][2] , \mult_20/CARRYB[13][3] ,
         \mult_20/CARRYB[13][4] , \mult_20/CARRYB[13][5] ,
         \mult_20/CARRYB[13][6] , \mult_20/CARRYB[13][7] ,
         \mult_20/CARRYB[13][8] , \mult_20/CARRYB[13][9] ,
         \mult_20/CARRYB[13][10] , \mult_20/CARRYB[13][11] ,
         \mult_20/CARRYB[13][12] , \mult_20/CARRYB[13][13] ,
         \mult_20/CARRYB[13][14] , \mult_20/CARRYB[13][15] ,
         \mult_20/CARRYB[13][16] , \mult_20/CARRYB[13][17] ,
         \mult_20/CARRYB[13][18] , \mult_20/CARRYB[13][19] ,
         \mult_20/CARRYB[13][20] , \mult_20/CARRYB[13][21] ,
         \mult_20/CARRYB[13][22] , \mult_20/CARRYB[13][23] ,
         \mult_20/CARRYB[13][24] , \mult_20/CARRYB[13][25] ,
         \mult_20/CARRYB[13][26] , \mult_20/CARRYB[13][27] ,
         \mult_20/CARRYB[13][28] , \mult_20/CARRYB[13][29] ,
         \mult_20/CARRYB[13][30] , \mult_20/CARRYB[14][0] ,
         \mult_20/CARRYB[14][1] , \mult_20/CARRYB[14][2] ,
         \mult_20/CARRYB[14][3] , \mult_20/CARRYB[14][4] ,
         \mult_20/CARRYB[14][5] , \mult_20/CARRYB[14][6] ,
         \mult_20/CARRYB[14][7] , \mult_20/CARRYB[14][8] ,
         \mult_20/CARRYB[14][9] , \mult_20/CARRYB[14][10] ,
         \mult_20/CARRYB[14][11] , \mult_20/CARRYB[14][12] ,
         \mult_20/CARRYB[14][13] , \mult_20/CARRYB[14][14] ,
         \mult_20/CARRYB[14][15] , \mult_20/CARRYB[14][16] ,
         \mult_20/CARRYB[14][17] , \mult_20/CARRYB[14][18] ,
         \mult_20/CARRYB[14][19] , \mult_20/CARRYB[14][20] ,
         \mult_20/CARRYB[14][21] , \mult_20/CARRYB[14][22] ,
         \mult_20/CARRYB[14][23] , \mult_20/CARRYB[14][24] ,
         \mult_20/CARRYB[14][25] , \mult_20/CARRYB[14][26] ,
         \mult_20/CARRYB[14][27] , \mult_20/CARRYB[14][28] ,
         \mult_20/CARRYB[14][29] , \mult_20/CARRYB[14][30] ,
         \mult_20/CARRYB[15][0] , \mult_20/CARRYB[15][1] ,
         \mult_20/CARRYB[15][2] , \mult_20/CARRYB[15][3] ,
         \mult_20/CARRYB[15][4] , \mult_20/CARRYB[15][5] ,
         \mult_20/CARRYB[15][6] , \mult_20/CARRYB[15][7] ,
         \mult_20/CARRYB[15][8] , \mult_20/CARRYB[15][9] ,
         \mult_20/CARRYB[15][10] , \mult_20/CARRYB[15][11] ,
         \mult_20/CARRYB[15][12] , \mult_20/CARRYB[15][13] ,
         \mult_20/CARRYB[15][14] , \mult_20/CARRYB[15][15] ,
         \mult_20/CARRYB[15][16] , \mult_20/CARRYB[15][17] ,
         \mult_20/CARRYB[15][18] , \mult_20/CARRYB[15][19] ,
         \mult_20/CARRYB[15][20] , \mult_20/CARRYB[15][21] ,
         \mult_20/CARRYB[15][22] , \mult_20/CARRYB[15][23] ,
         \mult_20/CARRYB[15][24] , \mult_20/CARRYB[15][25] ,
         \mult_20/CARRYB[15][26] , \mult_20/CARRYB[15][27] ,
         \mult_20/CARRYB[15][28] , \mult_20/CARRYB[15][29] ,
         \mult_20/CARRYB[15][30] , \mult_20/ab[1][31] , \mult_20/ab[2][0] ,
         \mult_20/ab[2][1] , \mult_20/ab[2][2] , \mult_20/ab[2][3] ,
         \mult_20/ab[2][4] , \mult_20/ab[2][5] , \mult_20/ab[2][6] ,
         \mult_20/ab[2][7] , \mult_20/ab[2][8] , \mult_20/ab[2][9] ,
         \mult_20/ab[2][10] , \mult_20/ab[2][11] , \mult_20/ab[2][12] ,
         \mult_20/ab[2][13] , \mult_20/ab[2][14] , \mult_20/ab[2][15] ,
         \mult_20/ab[2][16] , \mult_20/ab[2][17] , \mult_20/ab[2][18] ,
         \mult_20/ab[2][19] , \mult_20/ab[2][20] , \mult_20/ab[2][21] ,
         \mult_20/ab[2][22] , \mult_20/ab[2][23] , \mult_20/ab[2][24] ,
         \mult_20/ab[2][25] , \mult_20/ab[2][26] , \mult_20/ab[2][27] ,
         \mult_20/ab[2][28] , \mult_20/ab[2][29] , \mult_20/ab[2][30] ,
         \mult_20/ab[2][31] , \mult_20/ab[3][0] , \mult_20/ab[3][1] ,
         \mult_20/ab[3][2] , \mult_20/ab[3][3] , \mult_20/ab[3][4] ,
         \mult_20/ab[3][5] , \mult_20/ab[3][6] , \mult_20/ab[3][7] ,
         \mult_20/ab[3][8] , \mult_20/ab[3][9] , \mult_20/ab[3][10] ,
         \mult_20/ab[3][11] , \mult_20/ab[3][12] , \mult_20/ab[3][13] ,
         \mult_20/ab[3][14] , \mult_20/ab[3][15] , \mult_20/ab[3][16] ,
         \mult_20/ab[3][17] , \mult_20/ab[3][18] , \mult_20/ab[3][19] ,
         \mult_20/ab[3][20] , \mult_20/ab[3][21] , \mult_20/ab[3][22] ,
         \mult_20/ab[3][23] , \mult_20/ab[3][24] , \mult_20/ab[3][25] ,
         \mult_20/ab[3][26] , \mult_20/ab[3][27] , \mult_20/ab[3][28] ,
         \mult_20/ab[3][29] , \mult_20/ab[3][30] , \mult_20/ab[3][31] ,
         \mult_20/ab[4][0] , \mult_20/ab[4][1] , \mult_20/ab[4][2] ,
         \mult_20/ab[4][3] , \mult_20/ab[4][4] , \mult_20/ab[4][5] ,
         \mult_20/ab[4][6] , \mult_20/ab[4][7] , \mult_20/ab[4][8] ,
         \mult_20/ab[4][9] , \mult_20/ab[4][10] , \mult_20/ab[4][11] ,
         \mult_20/ab[4][12] , \mult_20/ab[4][13] , \mult_20/ab[4][14] ,
         \mult_20/ab[4][15] , \mult_20/ab[4][16] , \mult_20/ab[4][17] ,
         \mult_20/ab[4][18] , \mult_20/ab[4][19] , \mult_20/ab[4][20] ,
         \mult_20/ab[4][21] , \mult_20/ab[4][22] , \mult_20/ab[4][23] ,
         \mult_20/ab[4][24] , \mult_20/ab[4][25] , \mult_20/ab[4][26] ,
         \mult_20/ab[4][27] , \mult_20/ab[4][28] , \mult_20/ab[4][29] ,
         \mult_20/ab[4][30] , \mult_20/ab[4][31] , \mult_20/ab[5][0] ,
         \mult_20/ab[5][1] , \mult_20/ab[5][2] , \mult_20/ab[5][3] ,
         \mult_20/ab[5][4] , \mult_20/ab[5][5] , \mult_20/ab[5][6] ,
         \mult_20/ab[5][7] , \mult_20/ab[5][8] , \mult_20/ab[5][9] ,
         \mult_20/ab[5][10] , \mult_20/ab[5][11] , \mult_20/ab[5][12] ,
         \mult_20/ab[5][13] , \mult_20/ab[5][14] , \mult_20/ab[5][15] ,
         \mult_20/ab[5][16] , \mult_20/ab[5][17] , \mult_20/ab[5][18] ,
         \mult_20/ab[5][19] , \mult_20/ab[5][20] , \mult_20/ab[5][21] ,
         \mult_20/ab[5][22] , \mult_20/ab[5][23] , \mult_20/ab[5][24] ,
         \mult_20/ab[5][25] , \mult_20/ab[5][26] , \mult_20/ab[5][27] ,
         \mult_20/ab[5][28] , \mult_20/ab[5][29] , \mult_20/ab[5][30] ,
         \mult_20/ab[5][31] , \mult_20/ab[6][0] , \mult_20/ab[6][1] ,
         \mult_20/ab[6][2] , \mult_20/ab[6][3] , \mult_20/ab[6][4] ,
         \mult_20/ab[6][5] , \mult_20/ab[6][6] , \mult_20/ab[6][7] ,
         \mult_20/ab[6][8] , \mult_20/ab[6][9] , \mult_20/ab[6][10] ,
         \mult_20/ab[6][11] , \mult_20/ab[6][12] , \mult_20/ab[6][13] ,
         \mult_20/ab[6][14] , \mult_20/ab[6][15] , \mult_20/ab[6][16] ,
         \mult_20/ab[6][17] , \mult_20/ab[6][18] , \mult_20/ab[6][19] ,
         \mult_20/ab[6][20] , \mult_20/ab[6][21] , \mult_20/ab[6][22] ,
         \mult_20/ab[6][23] , \mult_20/ab[6][24] , \mult_20/ab[6][25] ,
         \mult_20/ab[6][26] , \mult_20/ab[6][27] , \mult_20/ab[6][28] ,
         \mult_20/ab[6][29] , \mult_20/ab[6][30] , \mult_20/ab[6][31] ,
         \mult_20/ab[7][0] , \mult_20/ab[7][1] , \mult_20/ab[7][2] ,
         \mult_20/ab[7][3] , \mult_20/ab[7][4] , \mult_20/ab[7][5] ,
         \mult_20/ab[7][6] , \mult_20/ab[7][7] , \mult_20/ab[7][8] ,
         \mult_20/ab[7][9] , \mult_20/ab[7][10] , \mult_20/ab[7][11] ,
         \mult_20/ab[7][12] , \mult_20/ab[7][13] , \mult_20/ab[7][14] ,
         \mult_20/ab[7][15] , \mult_20/ab[7][16] , \mult_20/ab[7][17] ,
         \mult_20/ab[7][18] , \mult_20/ab[7][19] , \mult_20/ab[7][20] ,
         \mult_20/ab[7][21] , \mult_20/ab[7][22] , \mult_20/ab[7][23] ,
         \mult_20/ab[7][24] , \mult_20/ab[7][25] , \mult_20/ab[7][26] ,
         \mult_20/ab[7][27] , \mult_20/ab[7][28] , \mult_20/ab[7][29] ,
         \mult_20/ab[7][30] , \mult_20/ab[7][31] , \mult_20/ab[8][0] ,
         \mult_20/ab[8][1] , \mult_20/ab[8][2] , \mult_20/ab[8][3] ,
         \mult_20/ab[8][4] , \mult_20/ab[8][5] , \mult_20/ab[8][6] ,
         \mult_20/ab[8][7] , \mult_20/ab[8][8] , \mult_20/ab[8][9] ,
         \mult_20/ab[8][10] , \mult_20/ab[8][11] , \mult_20/ab[8][12] ,
         \mult_20/ab[8][13] , \mult_20/ab[8][14] , \mult_20/ab[8][15] ,
         \mult_20/ab[8][16] , \mult_20/ab[8][17] , \mult_20/ab[8][18] ,
         \mult_20/ab[8][19] , \mult_20/ab[8][20] , \mult_20/ab[8][21] ,
         \mult_20/ab[8][22] , \mult_20/ab[8][23] , \mult_20/ab[8][24] ,
         \mult_20/ab[8][25] , \mult_20/ab[8][26] , \mult_20/ab[8][27] ,
         \mult_20/ab[8][28] , \mult_20/ab[8][29] , \mult_20/ab[8][30] ,
         \mult_20/ab[8][31] , \mult_20/ab[9][0] , \mult_20/ab[9][1] ,
         \mult_20/ab[9][2] , \mult_20/ab[9][3] , \mult_20/ab[9][4] ,
         \mult_20/ab[9][5] , \mult_20/ab[9][6] , \mult_20/ab[9][7] ,
         \mult_20/ab[9][8] , \mult_20/ab[9][9] , \mult_20/ab[9][10] ,
         \mult_20/ab[9][11] , \mult_20/ab[9][12] , \mult_20/ab[9][13] ,
         \mult_20/ab[9][14] , \mult_20/ab[9][15] , \mult_20/ab[9][16] ,
         \mult_20/ab[9][17] , \mult_20/ab[9][18] , \mult_20/ab[9][19] ,
         \mult_20/ab[9][20] , \mult_20/ab[9][21] , \mult_20/ab[9][22] ,
         \mult_20/ab[9][23] , \mult_20/ab[9][24] , \mult_20/ab[9][25] ,
         \mult_20/ab[9][26] , \mult_20/ab[9][27] , \mult_20/ab[9][28] ,
         \mult_20/ab[9][29] , \mult_20/ab[9][30] , \mult_20/ab[9][31] ,
         \mult_20/ab[10][0] , \mult_20/ab[10][1] , \mult_20/ab[10][2] ,
         \mult_20/ab[10][3] , \mult_20/ab[10][4] , \mult_20/ab[10][5] ,
         \mult_20/ab[10][6] , \mult_20/ab[10][7] , \mult_20/ab[10][8] ,
         \mult_20/ab[10][9] , \mult_20/ab[10][10] , \mult_20/ab[10][11] ,
         \mult_20/ab[10][12] , \mult_20/ab[10][13] , \mult_20/ab[10][14] ,
         \mult_20/ab[10][15] , \mult_20/ab[10][16] , \mult_20/ab[10][17] ,
         \mult_20/ab[10][18] , \mult_20/ab[10][19] , \mult_20/ab[10][20] ,
         \mult_20/ab[10][21] , \mult_20/ab[10][22] , \mult_20/ab[10][23] ,
         \mult_20/ab[10][24] , \mult_20/ab[10][25] , \mult_20/ab[10][26] ,
         \mult_20/ab[10][27] , \mult_20/ab[10][28] , \mult_20/ab[10][29] ,
         \mult_20/ab[10][30] , \mult_20/ab[10][31] , \mult_20/ab[11][0] ,
         \mult_20/ab[11][1] , \mult_20/ab[11][2] , \mult_20/ab[11][3] ,
         \mult_20/ab[11][4] , \mult_20/ab[11][5] , \mult_20/ab[11][6] ,
         \mult_20/ab[11][7] , \mult_20/ab[11][8] , \mult_20/ab[11][9] ,
         \mult_20/ab[11][10] , \mult_20/ab[11][11] , \mult_20/ab[11][12] ,
         \mult_20/ab[11][13] , \mult_20/ab[11][14] , \mult_20/ab[11][15] ,
         \mult_20/ab[11][16] , \mult_20/ab[11][17] , \mult_20/ab[11][18] ,
         \mult_20/ab[11][19] , \mult_20/ab[11][20] , \mult_20/ab[11][21] ,
         \mult_20/ab[11][22] , \mult_20/ab[11][23] , \mult_20/ab[11][24] ,
         \mult_20/ab[11][25] , \mult_20/ab[11][26] , \mult_20/ab[11][27] ,
         \mult_20/ab[11][28] , \mult_20/ab[11][29] , \mult_20/ab[11][30] ,
         \mult_20/ab[11][31] , \mult_20/ab[12][0] , \mult_20/ab[12][1] ,
         \mult_20/ab[12][2] , \mult_20/ab[12][3] , \mult_20/ab[12][4] ,
         \mult_20/ab[12][5] , \mult_20/ab[12][6] , \mult_20/ab[12][7] ,
         \mult_20/ab[12][8] , \mult_20/ab[12][9] , \mult_20/ab[12][10] ,
         \mult_20/ab[12][11] , \mult_20/ab[12][12] , \mult_20/ab[12][13] ,
         \mult_20/ab[12][14] , \mult_20/ab[12][15] , \mult_20/ab[12][16] ,
         \mult_20/ab[12][17] , \mult_20/ab[12][18] , \mult_20/ab[12][19] ,
         \mult_20/ab[12][20] , \mult_20/ab[12][21] , \mult_20/ab[12][22] ,
         \mult_20/ab[12][23] , \mult_20/ab[12][24] , \mult_20/ab[12][25] ,
         \mult_20/ab[12][26] , \mult_20/ab[12][27] , \mult_20/ab[12][28] ,
         \mult_20/ab[12][29] , \mult_20/ab[12][30] , \mult_20/ab[12][31] ,
         \mult_20/ab[13][0] , \mult_20/ab[13][1] , \mult_20/ab[13][2] ,
         \mult_20/ab[13][3] , \mult_20/ab[13][4] , \mult_20/ab[13][5] ,
         \mult_20/ab[13][6] , \mult_20/ab[13][7] , \mult_20/ab[13][8] ,
         \mult_20/ab[13][9] , \mult_20/ab[13][10] , \mult_20/ab[13][11] ,
         \mult_20/ab[13][12] , \mult_20/ab[13][13] , \mult_20/ab[13][14] ,
         \mult_20/ab[13][15] , \mult_20/ab[13][16] , \mult_20/ab[13][17] ,
         \mult_20/ab[13][18] , \mult_20/ab[13][19] , \mult_20/ab[13][20] ,
         \mult_20/ab[13][21] , \mult_20/ab[13][22] , \mult_20/ab[13][23] ,
         \mult_20/ab[13][24] , \mult_20/ab[13][25] , \mult_20/ab[13][26] ,
         \mult_20/ab[13][27] , \mult_20/ab[13][28] , \mult_20/ab[13][29] ,
         \mult_20/ab[13][30] , \mult_20/ab[13][31] , \mult_20/ab[14][0] ,
         \mult_20/ab[14][1] , \mult_20/ab[14][2] , \mult_20/ab[14][3] ,
         \mult_20/ab[14][4] , \mult_20/ab[14][5] , \mult_20/ab[14][6] ,
         \mult_20/ab[14][7] , \mult_20/ab[14][8] , \mult_20/ab[14][9] ,
         \mult_20/ab[14][10] , \mult_20/ab[14][11] , \mult_20/ab[14][12] ,
         \mult_20/ab[14][13] , \mult_20/ab[14][14] , \mult_20/ab[14][15] ,
         \mult_20/ab[14][16] , \mult_20/ab[14][17] , \mult_20/ab[14][18] ,
         \mult_20/ab[14][19] , \mult_20/ab[14][20] , \mult_20/ab[14][21] ,
         \mult_20/ab[14][22] , \mult_20/ab[14][23] , \mult_20/ab[14][24] ,
         \mult_20/ab[14][25] , \mult_20/ab[14][26] , \mult_20/ab[14][27] ,
         \mult_20/ab[14][28] , \mult_20/ab[14][29] , \mult_20/ab[14][30] ,
         \mult_20/ab[14][31] , \mult_20/ab[15][0] , \mult_20/ab[15][1] ,
         \mult_20/ab[15][2] , \mult_20/ab[15][3] , \mult_20/ab[15][4] ,
         \mult_20/ab[15][5] , \mult_20/ab[15][6] , \mult_20/ab[15][7] ,
         \mult_20/ab[15][8] , \mult_20/ab[15][9] , \mult_20/ab[15][10] ,
         \mult_20/ab[15][11] , \mult_20/ab[15][12] , \mult_20/ab[15][13] ,
         \mult_20/ab[15][14] , \mult_20/ab[15][15] , \mult_20/ab[15][16] ,
         \mult_20/ab[15][17] , \mult_20/ab[15][18] , \mult_20/ab[15][19] ,
         \mult_20/ab[15][20] , \mult_20/ab[15][21] , \mult_20/ab[15][22] ,
         \mult_20/ab[15][23] , \mult_20/ab[15][24] , \mult_20/ab[15][25] ,
         \mult_20/ab[15][26] , \mult_20/ab[15][27] , \mult_20/ab[15][28] ,
         \mult_20/ab[15][29] , \mult_20/ab[15][30] , \mult_20/ab[15][31] ,
         \mult_20/ab[16][0] , \mult_20/ab[16][1] , \mult_20/ab[16][2] ,
         \mult_20/ab[16][3] , \mult_20/ab[16][4] , \mult_20/ab[16][5] ,
         \mult_20/ab[16][6] , \mult_20/ab[16][7] , \mult_20/ab[16][8] ,
         \mult_20/ab[16][9] , \mult_20/ab[16][10] , \mult_20/ab[16][11] ,
         \mult_20/ab[16][12] , \mult_20/ab[16][13] , \mult_20/ab[16][14] ,
         \mult_20/ab[16][15] , \mult_20/ab[16][16] , \mult_20/ab[16][17] ,
         \mult_20/ab[16][18] , \mult_20/ab[16][19] , \mult_20/ab[16][20] ,
         \mult_20/ab[16][21] , \mult_20/ab[16][22] , \mult_20/ab[16][23] ,
         \mult_20/ab[16][24] , \mult_20/ab[16][25] , \mult_20/ab[16][26] ,
         \mult_20/ab[16][27] , \mult_20/ab[16][28] , \mult_20/ab[16][29] ,
         \mult_20/ab[16][30] , \mult_20/ab[16][31] , \mult_20/ab[17][0] ,
         \mult_20/ab[17][1] , \mult_20/ab[17][2] , \mult_20/ab[17][3] ,
         \mult_20/ab[17][4] , \mult_20/ab[17][5] , \mult_20/ab[17][6] ,
         \mult_20/ab[17][7] , \mult_20/ab[17][8] , \mult_20/ab[17][9] ,
         \mult_20/ab[17][10] , \mult_20/ab[17][11] , \mult_20/ab[17][12] ,
         \mult_20/ab[17][13] , \mult_20/ab[17][14] , \mult_20/ab[17][15] ,
         \mult_20/ab[17][16] , \mult_20/ab[17][17] , \mult_20/ab[17][18] ,
         \mult_20/ab[17][19] , \mult_20/ab[17][20] , \mult_20/ab[17][21] ,
         \mult_20/ab[17][22] , \mult_20/ab[17][23] , \mult_20/ab[17][24] ,
         \mult_20/ab[17][25] , \mult_20/ab[17][26] , \mult_20/ab[17][27] ,
         \mult_20/ab[17][28] , \mult_20/ab[17][29] , \mult_20/ab[17][30] ,
         \mult_20/ab[17][31] , \mult_20/ab[18][0] , \mult_20/ab[18][1] ,
         \mult_20/ab[18][2] , \mult_20/ab[18][3] , \mult_20/ab[18][4] ,
         \mult_20/ab[18][5] , \mult_20/ab[18][6] , \mult_20/ab[18][7] ,
         \mult_20/ab[18][8] , \mult_20/ab[18][9] , \mult_20/ab[18][10] ,
         \mult_20/ab[18][11] , \mult_20/ab[18][12] , \mult_20/ab[18][13] ,
         \mult_20/ab[18][14] , \mult_20/ab[18][15] , \mult_20/ab[18][16] ,
         \mult_20/ab[18][17] , \mult_20/ab[18][18] , \mult_20/ab[18][19] ,
         \mult_20/ab[18][20] , \mult_20/ab[18][21] , \mult_20/ab[18][22] ,
         \mult_20/ab[18][23] , \mult_20/ab[18][24] , \mult_20/ab[18][25] ,
         \mult_20/ab[18][26] , \mult_20/ab[18][27] , \mult_20/ab[18][28] ,
         \mult_20/ab[18][29] , \mult_20/ab[18][30] , \mult_20/ab[18][31] ,
         \mult_20/ab[19][0] , \mult_20/ab[19][1] , \mult_20/ab[19][2] ,
         \mult_20/ab[19][3] , \mult_20/ab[19][4] , \mult_20/ab[19][5] ,
         \mult_20/ab[19][6] , \mult_20/ab[19][7] , \mult_20/ab[19][8] ,
         \mult_20/ab[19][9] , \mult_20/ab[19][10] , \mult_20/ab[19][11] ,
         \mult_20/ab[19][12] , \mult_20/ab[19][13] , \mult_20/ab[19][14] ,
         \mult_20/ab[19][15] , \mult_20/ab[19][16] , \mult_20/ab[19][17] ,
         \mult_20/ab[19][18] , \mult_20/ab[19][19] , \mult_20/ab[19][20] ,
         \mult_20/ab[19][21] , \mult_20/ab[19][22] , \mult_20/ab[19][23] ,
         \mult_20/ab[19][24] , \mult_20/ab[19][25] , \mult_20/ab[19][26] ,
         \mult_20/ab[19][27] , \mult_20/ab[19][28] , \mult_20/ab[19][29] ,
         \mult_20/ab[19][30] , \mult_20/ab[19][31] , \mult_20/ab[20][0] ,
         \mult_20/ab[20][1] , \mult_20/ab[20][2] , \mult_20/ab[20][3] ,
         \mult_20/ab[20][4] , \mult_20/ab[20][5] , \mult_20/ab[20][6] ,
         \mult_20/ab[20][7] , \mult_20/ab[20][8] , \mult_20/ab[20][9] ,
         \mult_20/ab[20][10] , \mult_20/ab[20][11] , \mult_20/ab[20][12] ,
         \mult_20/ab[20][13] , \mult_20/ab[20][14] , \mult_20/ab[20][15] ,
         \mult_20/ab[20][16] , \mult_20/ab[20][17] , \mult_20/ab[20][18] ,
         \mult_20/ab[20][19] , \mult_20/ab[20][20] , \mult_20/ab[20][21] ,
         \mult_20/ab[20][22] , \mult_20/ab[20][23] , \mult_20/ab[20][24] ,
         \mult_20/ab[20][25] , \mult_20/ab[20][26] , \mult_20/ab[20][27] ,
         \mult_20/ab[20][28] , \mult_20/ab[20][29] , \mult_20/ab[20][30] ,
         \mult_20/ab[20][31] , \mult_20/ab[21][0] , \mult_20/ab[21][1] ,
         \mult_20/ab[21][2] , \mult_20/ab[21][3] , \mult_20/ab[21][4] ,
         \mult_20/ab[21][5] , \mult_20/ab[21][6] , \mult_20/ab[21][7] ,
         \mult_20/ab[21][8] , \mult_20/ab[21][9] , \mult_20/ab[21][10] ,
         \mult_20/ab[21][11] , \mult_20/ab[21][12] , \mult_20/ab[21][13] ,
         \mult_20/ab[21][14] , \mult_20/ab[21][15] , \mult_20/ab[21][16] ,
         \mult_20/ab[21][17] , \mult_20/ab[21][18] , \mult_20/ab[21][19] ,
         \mult_20/ab[21][20] , \mult_20/ab[21][21] , \mult_20/ab[21][22] ,
         \mult_20/ab[21][23] , \mult_20/ab[21][24] , \mult_20/ab[21][25] ,
         \mult_20/ab[21][26] , \mult_20/ab[21][27] , \mult_20/ab[21][28] ,
         \mult_20/ab[21][29] , \mult_20/ab[21][30] , \mult_20/ab[21][31] ,
         \mult_20/ab[22][0] , \mult_20/ab[22][1] , \mult_20/ab[22][2] ,
         \mult_20/ab[22][3] , \mult_20/ab[22][4] , \mult_20/ab[22][5] ,
         \mult_20/ab[22][6] , \mult_20/ab[22][7] , \mult_20/ab[22][8] ,
         \mult_20/ab[22][9] , \mult_20/ab[22][10] , \mult_20/ab[22][11] ,
         \mult_20/ab[22][12] , \mult_20/ab[22][13] , \mult_20/ab[22][14] ,
         \mult_20/ab[22][15] , \mult_20/ab[22][16] , \mult_20/ab[22][17] ,
         \mult_20/ab[22][18] , \mult_20/ab[22][19] , \mult_20/ab[22][20] ,
         \mult_20/ab[22][21] , \mult_20/ab[22][22] , \mult_20/ab[22][23] ,
         \mult_20/ab[22][24] , \mult_20/ab[22][25] , \mult_20/ab[22][26] ,
         \mult_20/ab[22][27] , \mult_20/ab[22][28] , \mult_20/ab[22][29] ,
         \mult_20/ab[22][30] , \mult_20/ab[22][31] , \mult_20/ab[23][0] ,
         \mult_20/ab[23][1] , \mult_20/ab[23][2] , \mult_20/ab[23][3] ,
         \mult_20/ab[23][4] , \mult_20/ab[23][5] , \mult_20/ab[23][6] ,
         \mult_20/ab[23][7] , \mult_20/ab[23][8] , \mult_20/ab[23][9] ,
         \mult_20/ab[23][10] , \mult_20/ab[23][11] , \mult_20/ab[23][12] ,
         \mult_20/ab[23][13] , \mult_20/ab[23][14] , \mult_20/ab[23][15] ,
         \mult_20/ab[23][16] , \mult_20/ab[23][17] , \mult_20/ab[23][18] ,
         \mult_20/ab[23][19] , \mult_20/ab[23][20] , \mult_20/ab[23][21] ,
         \mult_20/ab[23][22] , \mult_20/ab[23][23] , \mult_20/ab[23][24] ,
         \mult_20/ab[23][25] , \mult_20/ab[23][26] , \mult_20/ab[23][27] ,
         \mult_20/ab[23][28] , \mult_20/ab[23][29] , \mult_20/ab[23][30] ,
         \mult_20/ab[23][31] , \mult_20/ab[24][0] , \mult_20/ab[24][1] ,
         \mult_20/ab[24][2] , \mult_20/ab[24][3] , \mult_20/ab[24][4] ,
         \mult_20/ab[24][5] , \mult_20/ab[24][6] , \mult_20/ab[24][7] ,
         \mult_20/ab[24][8] , \mult_20/ab[24][9] , \mult_20/ab[24][10] ,
         \mult_20/ab[24][11] , \mult_20/ab[24][12] , \mult_20/ab[24][13] ,
         \mult_20/ab[24][14] , \mult_20/ab[24][15] , \mult_20/ab[24][16] ,
         \mult_20/ab[24][17] , \mult_20/ab[24][18] , \mult_20/ab[24][19] ,
         \mult_20/ab[24][20] , \mult_20/ab[24][21] , \mult_20/ab[24][22] ,
         \mult_20/ab[24][23] , \mult_20/ab[24][24] , \mult_20/ab[24][25] ,
         \mult_20/ab[24][26] , \mult_20/ab[24][27] , \mult_20/ab[24][28] ,
         \mult_20/ab[24][29] , \mult_20/ab[24][30] , \mult_20/ab[24][31] ,
         \mult_20/ab[25][0] , \mult_20/ab[25][1] , \mult_20/ab[25][2] ,
         \mult_20/ab[25][3] , \mult_20/ab[25][4] , \mult_20/ab[25][5] ,
         \mult_20/ab[25][6] , \mult_20/ab[25][7] , \mult_20/ab[25][8] ,
         \mult_20/ab[25][9] , \mult_20/ab[25][10] , \mult_20/ab[25][11] ,
         \mult_20/ab[25][12] , \mult_20/ab[25][13] , \mult_20/ab[25][14] ,
         \mult_20/ab[25][15] , \mult_20/ab[25][16] , \mult_20/ab[25][17] ,
         \mult_20/ab[25][18] , \mult_20/ab[25][19] , \mult_20/ab[25][20] ,
         \mult_20/ab[25][21] , \mult_20/ab[25][22] , \mult_20/ab[25][23] ,
         \mult_20/ab[25][24] , \mult_20/ab[25][25] , \mult_20/ab[25][26] ,
         \mult_20/ab[25][27] , \mult_20/ab[25][28] , \mult_20/ab[25][29] ,
         \mult_20/ab[25][30] , \mult_20/ab[25][31] , \mult_20/ab[26][0] ,
         \mult_20/ab[26][1] , \mult_20/ab[26][2] , \mult_20/ab[26][3] ,
         \mult_20/ab[26][4] , \mult_20/ab[26][5] , \mult_20/ab[26][6] ,
         \mult_20/ab[26][7] , \mult_20/ab[26][8] , \mult_20/ab[26][9] ,
         \mult_20/ab[26][10] , \mult_20/ab[26][11] , \mult_20/ab[26][12] ,
         \mult_20/ab[26][13] , \mult_20/ab[26][14] , \mult_20/ab[26][15] ,
         \mult_20/ab[26][16] , \mult_20/ab[26][17] , \mult_20/ab[26][18] ,
         \mult_20/ab[26][19] , \mult_20/ab[26][20] , \mult_20/ab[26][21] ,
         \mult_20/ab[26][22] , \mult_20/ab[26][23] , \mult_20/ab[26][24] ,
         \mult_20/ab[26][25] , \mult_20/ab[26][26] , \mult_20/ab[26][27] ,
         \mult_20/ab[26][28] , \mult_20/ab[26][29] , \mult_20/ab[26][30] ,
         \mult_20/ab[26][31] , \mult_20/ab[27][0] , \mult_20/ab[27][1] ,
         \mult_20/ab[27][2] , \mult_20/ab[27][3] , \mult_20/ab[27][4] ,
         \mult_20/ab[27][5] , \mult_20/ab[27][6] , \mult_20/ab[27][7] ,
         \mult_20/ab[27][8] , \mult_20/ab[27][9] , \mult_20/ab[27][10] ,
         \mult_20/ab[27][11] , \mult_20/ab[27][12] , \mult_20/ab[27][13] ,
         \mult_20/ab[27][14] , \mult_20/ab[27][15] , \mult_20/ab[27][16] ,
         \mult_20/ab[27][17] , \mult_20/ab[27][18] , \mult_20/ab[27][19] ,
         \mult_20/ab[27][20] , \mult_20/ab[27][21] , \mult_20/ab[27][22] ,
         \mult_20/ab[27][23] , \mult_20/ab[27][24] , \mult_20/ab[27][25] ,
         \mult_20/ab[27][26] , \mult_20/ab[27][27] , \mult_20/ab[27][28] ,
         \mult_20/ab[27][29] , \mult_20/ab[27][30] , \mult_20/ab[27][31] ,
         \mult_20/ab[28][0] , \mult_20/ab[28][1] , \mult_20/ab[28][2] ,
         \mult_20/ab[28][3] , \mult_20/ab[28][4] , \mult_20/ab[28][5] ,
         \mult_20/ab[28][6] , \mult_20/ab[28][7] , \mult_20/ab[28][8] ,
         \mult_20/ab[28][9] , \mult_20/ab[28][10] , \mult_20/ab[28][11] ,
         \mult_20/ab[28][12] , \mult_20/ab[28][13] , \mult_20/ab[28][14] ,
         \mult_20/ab[28][15] , \mult_20/ab[28][16] , \mult_20/ab[28][17] ,
         \mult_20/ab[28][18] , \mult_20/ab[28][19] , \mult_20/ab[28][20] ,
         \mult_20/ab[28][21] , \mult_20/ab[28][22] , \mult_20/ab[28][23] ,
         \mult_20/ab[28][24] , \mult_20/ab[28][25] , \mult_20/ab[28][26] ,
         \mult_20/ab[28][27] , \mult_20/ab[28][28] , \mult_20/ab[28][29] ,
         \mult_20/ab[28][30] , \mult_20/ab[28][31] , \mult_20/ab[29][0] ,
         \mult_20/ab[29][1] , \mult_20/ab[29][2] , \mult_20/ab[29][3] ,
         \mult_20/ab[29][4] , \mult_20/ab[29][5] , \mult_20/ab[29][6] ,
         \mult_20/ab[29][7] , \mult_20/ab[29][8] , \mult_20/ab[29][9] ,
         \mult_20/ab[29][10] , \mult_20/ab[29][11] , \mult_20/ab[29][12] ,
         \mult_20/ab[29][13] , \mult_20/ab[29][14] , \mult_20/ab[29][15] ,
         \mult_20/ab[29][16] , \mult_20/ab[29][17] , \mult_20/ab[29][18] ,
         \mult_20/ab[29][19] , \mult_20/ab[29][20] , \mult_20/ab[29][21] ,
         \mult_20/ab[29][22] , \mult_20/ab[29][23] , \mult_20/ab[29][24] ,
         \mult_20/ab[29][25] , \mult_20/ab[29][26] , \mult_20/ab[29][27] ,
         \mult_20/ab[29][28] , \mult_20/ab[29][29] , \mult_20/ab[29][30] ,
         \mult_20/ab[29][31] , \mult_20/ab[30][0] , \mult_20/ab[30][1] ,
         \mult_20/ab[30][2] , \mult_20/ab[30][3] , \mult_20/ab[30][4] ,
         \mult_20/ab[30][5] , \mult_20/ab[30][6] , \mult_20/ab[30][7] ,
         \mult_20/ab[30][8] , \mult_20/ab[30][9] , \mult_20/ab[30][10] ,
         \mult_20/ab[30][11] , \mult_20/ab[30][12] , \mult_20/ab[30][13] ,
         \mult_20/ab[30][14] , \mult_20/ab[30][15] , \mult_20/ab[30][16] ,
         \mult_20/ab[30][17] , \mult_20/ab[30][18] , \mult_20/ab[30][19] ,
         \mult_20/ab[30][20] , \mult_20/ab[30][21] , \mult_20/ab[30][22] ,
         \mult_20/ab[30][23] , \mult_20/ab[30][24] , \mult_20/ab[30][25] ,
         \mult_20/ab[30][26] , \mult_20/ab[30][27] , \mult_20/ab[30][28] ,
         \mult_20/ab[30][29] , \mult_20/ab[30][30] , \mult_20/ab[30][31] ,
         \mult_20/ab[31][0] , \mult_20/ab[31][1] , \mult_20/ab[31][2] ,
         \mult_20/ab[31][3] , \mult_20/ab[31][4] , \mult_20/ab[31][5] ,
         \mult_20/ab[31][6] , \mult_20/ab[31][7] , \mult_20/ab[31][8] ,
         \mult_20/ab[31][9] , \mult_20/ab[31][10] , \mult_20/ab[31][11] ,
         \mult_20/ab[31][12] , \mult_20/ab[31][13] , \mult_20/ab[31][14] ,
         \mult_20/ab[31][15] , \mult_20/ab[31][16] , \mult_20/ab[31][17] ,
         \mult_20/ab[31][18] , \mult_20/ab[31][19] , \mult_20/ab[31][20] ,
         \mult_20/ab[31][21] , \mult_20/ab[31][22] , \mult_20/ab[31][23] ,
         \mult_20/ab[31][24] , \mult_20/ab[31][25] , \mult_20/ab[31][26] ,
         \mult_20/ab[31][27] , \mult_20/ab[31][28] , \mult_20/ab[31][29] ,
         \mult_20/ab[31][30] , \mult_19/n63 , \mult_19/n62 , \mult_19/n61 ,
         \mult_19/n60 , \mult_19/n59 , \mult_19/n58 , \mult_19/n57 ,
         \mult_19/n56 , \mult_19/n55 , \mult_19/n54 , \mult_19/n53 ,
         \mult_19/n52 , \mult_19/n51 , \mult_19/n50 , \mult_19/n49 ,
         \mult_19/n48 , \mult_19/n47 , \mult_19/n46 , \mult_19/n45 ,
         \mult_19/n44 , \mult_19/n43 , \mult_19/n42 , \mult_19/n41 ,
         \mult_19/n40 , \mult_19/n39 , \mult_19/n38 , \mult_19/n37 ,
         \mult_19/n36 , \mult_19/n35 , \mult_19/n34 , \mult_19/n33 ,
         \mult_19/n32 , \mult_19/n31 , \mult_19/n30 , \mult_19/n29 ,
         \mult_19/n28 , \mult_19/n27 , \mult_19/n26 , \mult_19/n25 ,
         \mult_19/n24 , \mult_19/n23 , \mult_19/n22 , \mult_19/n21 ,
         \mult_19/n20 , \mult_19/n19 , \mult_19/n18 , \mult_19/n17 ,
         \mult_19/n16 , \mult_19/n15 , \mult_19/n14 , \mult_19/n13 ,
         \mult_19/n12 , \mult_19/n11 , \mult_19/n10 , \mult_19/n9 ,
         \mult_19/n8 , \mult_19/n7 , \mult_19/n6 , \mult_19/n5 , \mult_19/n4 ,
         \mult_19/n3 , \mult_19/SUMB[16][1] , \mult_19/SUMB[16][2] ,
         \mult_19/SUMB[16][3] , \mult_19/SUMB[16][4] , \mult_19/SUMB[16][5] ,
         \mult_19/SUMB[16][6] , \mult_19/SUMB[16][7] , \mult_19/SUMB[16][8] ,
         \mult_19/SUMB[16][9] , \mult_19/SUMB[16][10] , \mult_19/SUMB[16][11] ,
         \mult_19/SUMB[16][12] , \mult_19/SUMB[16][13] ,
         \mult_19/SUMB[16][14] , \mult_19/SUMB[16][15] ,
         \mult_19/SUMB[16][16] , \mult_19/SUMB[16][17] ,
         \mult_19/SUMB[16][18] , \mult_19/SUMB[16][19] ,
         \mult_19/SUMB[16][20] , \mult_19/SUMB[16][21] ,
         \mult_19/SUMB[16][22] , \mult_19/SUMB[16][23] ,
         \mult_19/SUMB[16][24] , \mult_19/SUMB[16][25] ,
         \mult_19/SUMB[16][26] , \mult_19/SUMB[16][27] ,
         \mult_19/SUMB[16][28] , \mult_19/SUMB[16][29] ,
         \mult_19/SUMB[16][30] , \mult_19/SUMB[17][1] , \mult_19/SUMB[17][2] ,
         \mult_19/SUMB[17][3] , \mult_19/SUMB[17][4] , \mult_19/SUMB[17][5] ,
         \mult_19/SUMB[17][6] , \mult_19/SUMB[17][7] , \mult_19/SUMB[17][8] ,
         \mult_19/SUMB[17][9] , \mult_19/SUMB[17][10] , \mult_19/SUMB[17][11] ,
         \mult_19/SUMB[17][12] , \mult_19/SUMB[17][13] ,
         \mult_19/SUMB[17][14] , \mult_19/SUMB[17][15] ,
         \mult_19/SUMB[17][16] , \mult_19/SUMB[17][17] ,
         \mult_19/SUMB[17][18] , \mult_19/SUMB[17][19] ,
         \mult_19/SUMB[17][20] , \mult_19/SUMB[17][21] ,
         \mult_19/SUMB[17][22] , \mult_19/SUMB[17][23] ,
         \mult_19/SUMB[17][24] , \mult_19/SUMB[17][25] ,
         \mult_19/SUMB[17][26] , \mult_19/SUMB[17][27] ,
         \mult_19/SUMB[17][28] , \mult_19/SUMB[17][29] ,
         \mult_19/SUMB[17][30] , \mult_19/SUMB[18][1] , \mult_19/SUMB[18][2] ,
         \mult_19/SUMB[18][3] , \mult_19/SUMB[18][4] , \mult_19/SUMB[18][5] ,
         \mult_19/SUMB[18][6] , \mult_19/SUMB[18][7] , \mult_19/SUMB[18][8] ,
         \mult_19/SUMB[18][9] , \mult_19/SUMB[18][10] , \mult_19/SUMB[18][11] ,
         \mult_19/SUMB[18][12] , \mult_19/SUMB[18][13] ,
         \mult_19/SUMB[18][14] , \mult_19/SUMB[18][15] ,
         \mult_19/SUMB[18][16] , \mult_19/SUMB[18][17] ,
         \mult_19/SUMB[18][18] , \mult_19/SUMB[18][19] ,
         \mult_19/SUMB[18][20] , \mult_19/SUMB[18][21] ,
         \mult_19/SUMB[18][22] , \mult_19/SUMB[18][23] ,
         \mult_19/SUMB[18][24] , \mult_19/SUMB[18][25] ,
         \mult_19/SUMB[18][26] , \mult_19/SUMB[18][27] ,
         \mult_19/SUMB[18][28] , \mult_19/SUMB[18][29] ,
         \mult_19/SUMB[18][30] , \mult_19/SUMB[19][1] , \mult_19/SUMB[19][2] ,
         \mult_19/SUMB[19][3] , \mult_19/SUMB[19][4] , \mult_19/SUMB[19][5] ,
         \mult_19/SUMB[19][6] , \mult_19/SUMB[19][7] , \mult_19/SUMB[19][8] ,
         \mult_19/SUMB[19][9] , \mult_19/SUMB[19][10] , \mult_19/SUMB[19][11] ,
         \mult_19/SUMB[19][12] , \mult_19/SUMB[19][13] ,
         \mult_19/SUMB[19][14] , \mult_19/SUMB[19][15] ,
         \mult_19/SUMB[19][16] , \mult_19/SUMB[19][17] ,
         \mult_19/SUMB[19][18] , \mult_19/SUMB[19][19] ,
         \mult_19/SUMB[19][20] , \mult_19/SUMB[19][21] ,
         \mult_19/SUMB[19][22] , \mult_19/SUMB[19][23] ,
         \mult_19/SUMB[19][24] , \mult_19/SUMB[19][25] ,
         \mult_19/SUMB[19][26] , \mult_19/SUMB[19][27] ,
         \mult_19/SUMB[19][28] , \mult_19/SUMB[19][29] ,
         \mult_19/SUMB[19][30] , \mult_19/SUMB[20][1] , \mult_19/SUMB[20][2] ,
         \mult_19/SUMB[20][3] , \mult_19/SUMB[20][4] , \mult_19/SUMB[20][5] ,
         \mult_19/SUMB[20][6] , \mult_19/SUMB[20][7] , \mult_19/SUMB[20][8] ,
         \mult_19/SUMB[20][9] , \mult_19/SUMB[20][10] , \mult_19/SUMB[20][11] ,
         \mult_19/SUMB[20][12] , \mult_19/SUMB[20][13] ,
         \mult_19/SUMB[20][14] , \mult_19/SUMB[20][15] ,
         \mult_19/SUMB[20][16] , \mult_19/SUMB[20][17] ,
         \mult_19/SUMB[20][18] , \mult_19/SUMB[20][19] ,
         \mult_19/SUMB[20][20] , \mult_19/SUMB[20][21] ,
         \mult_19/SUMB[20][22] , \mult_19/SUMB[20][23] ,
         \mult_19/SUMB[20][24] , \mult_19/SUMB[20][25] ,
         \mult_19/SUMB[20][26] , \mult_19/SUMB[20][27] ,
         \mult_19/SUMB[20][28] , \mult_19/SUMB[20][29] ,
         \mult_19/SUMB[20][30] , \mult_19/SUMB[21][1] , \mult_19/SUMB[21][2] ,
         \mult_19/SUMB[21][3] , \mult_19/SUMB[21][4] , \mult_19/SUMB[21][5] ,
         \mult_19/SUMB[21][6] , \mult_19/SUMB[21][7] , \mult_19/SUMB[21][8] ,
         \mult_19/SUMB[21][9] , \mult_19/SUMB[21][10] , \mult_19/SUMB[21][11] ,
         \mult_19/SUMB[21][12] , \mult_19/SUMB[21][13] ,
         \mult_19/SUMB[21][14] , \mult_19/SUMB[21][15] ,
         \mult_19/SUMB[21][16] , \mult_19/SUMB[21][17] ,
         \mult_19/SUMB[21][18] , \mult_19/SUMB[21][19] ,
         \mult_19/SUMB[21][20] , \mult_19/SUMB[21][21] ,
         \mult_19/SUMB[21][22] , \mult_19/SUMB[21][23] ,
         \mult_19/SUMB[21][24] , \mult_19/SUMB[21][25] ,
         \mult_19/SUMB[21][26] , \mult_19/SUMB[21][27] ,
         \mult_19/SUMB[21][28] , \mult_19/SUMB[21][29] ,
         \mult_19/SUMB[21][30] , \mult_19/SUMB[22][1] , \mult_19/SUMB[22][2] ,
         \mult_19/SUMB[22][3] , \mult_19/SUMB[22][4] , \mult_19/SUMB[22][5] ,
         \mult_19/SUMB[22][6] , \mult_19/SUMB[22][7] , \mult_19/SUMB[22][8] ,
         \mult_19/SUMB[22][9] , \mult_19/SUMB[22][10] , \mult_19/SUMB[22][11] ,
         \mult_19/SUMB[22][12] , \mult_19/SUMB[22][13] ,
         \mult_19/SUMB[22][14] , \mult_19/SUMB[22][15] ,
         \mult_19/SUMB[22][16] , \mult_19/SUMB[22][17] ,
         \mult_19/SUMB[22][18] , \mult_19/SUMB[22][19] ,
         \mult_19/SUMB[22][20] , \mult_19/SUMB[22][21] ,
         \mult_19/SUMB[22][22] , \mult_19/SUMB[22][23] ,
         \mult_19/SUMB[22][24] , \mult_19/SUMB[22][25] ,
         \mult_19/SUMB[22][26] , \mult_19/SUMB[22][27] ,
         \mult_19/SUMB[22][28] , \mult_19/SUMB[22][29] ,
         \mult_19/SUMB[22][30] , \mult_19/SUMB[23][1] , \mult_19/SUMB[23][2] ,
         \mult_19/SUMB[23][3] , \mult_19/SUMB[23][4] , \mult_19/SUMB[23][5] ,
         \mult_19/SUMB[23][6] , \mult_19/SUMB[23][7] , \mult_19/SUMB[23][8] ,
         \mult_19/SUMB[23][9] , \mult_19/SUMB[23][10] , \mult_19/SUMB[23][11] ,
         \mult_19/SUMB[23][12] , \mult_19/SUMB[23][13] ,
         \mult_19/SUMB[23][14] , \mult_19/SUMB[23][15] ,
         \mult_19/SUMB[23][16] , \mult_19/SUMB[23][17] ,
         \mult_19/SUMB[23][18] , \mult_19/SUMB[23][19] ,
         \mult_19/SUMB[23][20] , \mult_19/SUMB[23][21] ,
         \mult_19/SUMB[23][22] , \mult_19/SUMB[23][23] ,
         \mult_19/SUMB[23][24] , \mult_19/SUMB[23][25] ,
         \mult_19/SUMB[23][26] , \mult_19/SUMB[23][27] ,
         \mult_19/SUMB[23][28] , \mult_19/SUMB[23][29] ,
         \mult_19/SUMB[23][30] , \mult_19/SUMB[24][1] , \mult_19/SUMB[24][2] ,
         \mult_19/SUMB[24][3] , \mult_19/SUMB[24][4] , \mult_19/SUMB[24][5] ,
         \mult_19/SUMB[24][6] , \mult_19/SUMB[24][7] , \mult_19/SUMB[24][8] ,
         \mult_19/SUMB[24][9] , \mult_19/SUMB[24][10] , \mult_19/SUMB[24][11] ,
         \mult_19/SUMB[24][12] , \mult_19/SUMB[24][13] ,
         \mult_19/SUMB[24][14] , \mult_19/SUMB[24][15] ,
         \mult_19/SUMB[24][16] , \mult_19/SUMB[24][17] ,
         \mult_19/SUMB[24][18] , \mult_19/SUMB[24][19] ,
         \mult_19/SUMB[24][20] , \mult_19/SUMB[24][21] ,
         \mult_19/SUMB[24][22] , \mult_19/SUMB[24][23] ,
         \mult_19/SUMB[24][24] , \mult_19/SUMB[24][25] ,
         \mult_19/SUMB[24][26] , \mult_19/SUMB[24][27] ,
         \mult_19/SUMB[24][28] , \mult_19/SUMB[24][29] ,
         \mult_19/SUMB[24][30] , \mult_19/SUMB[25][1] , \mult_19/SUMB[25][2] ,
         \mult_19/SUMB[25][3] , \mult_19/SUMB[25][4] , \mult_19/SUMB[25][5] ,
         \mult_19/SUMB[25][6] , \mult_19/SUMB[25][7] , \mult_19/SUMB[25][8] ,
         \mult_19/SUMB[25][9] , \mult_19/SUMB[25][10] , \mult_19/SUMB[25][11] ,
         \mult_19/SUMB[25][12] , \mult_19/SUMB[25][13] ,
         \mult_19/SUMB[25][14] , \mult_19/SUMB[25][15] ,
         \mult_19/SUMB[25][16] , \mult_19/SUMB[25][17] ,
         \mult_19/SUMB[25][18] , \mult_19/SUMB[25][19] ,
         \mult_19/SUMB[25][20] , \mult_19/SUMB[25][21] ,
         \mult_19/SUMB[25][22] , \mult_19/SUMB[25][23] ,
         \mult_19/SUMB[25][24] , \mult_19/SUMB[25][25] ,
         \mult_19/SUMB[25][26] , \mult_19/SUMB[25][27] ,
         \mult_19/SUMB[25][28] , \mult_19/SUMB[25][29] ,
         \mult_19/SUMB[25][30] , \mult_19/SUMB[26][1] , \mult_19/SUMB[26][2] ,
         \mult_19/SUMB[26][3] , \mult_19/SUMB[26][4] , \mult_19/SUMB[26][5] ,
         \mult_19/SUMB[26][6] , \mult_19/SUMB[26][7] , \mult_19/SUMB[26][8] ,
         \mult_19/SUMB[26][9] , \mult_19/SUMB[26][10] , \mult_19/SUMB[26][11] ,
         \mult_19/SUMB[26][12] , \mult_19/SUMB[26][13] ,
         \mult_19/SUMB[26][14] , \mult_19/SUMB[26][15] ,
         \mult_19/SUMB[26][16] , \mult_19/SUMB[26][17] ,
         \mult_19/SUMB[26][18] , \mult_19/SUMB[26][19] ,
         \mult_19/SUMB[26][20] , \mult_19/SUMB[26][21] ,
         \mult_19/SUMB[26][22] , \mult_19/SUMB[26][23] ,
         \mult_19/SUMB[26][24] , \mult_19/SUMB[26][25] ,
         \mult_19/SUMB[26][26] , \mult_19/SUMB[26][27] ,
         \mult_19/SUMB[26][28] , \mult_19/SUMB[26][29] ,
         \mult_19/SUMB[26][30] , \mult_19/SUMB[27][1] , \mult_19/SUMB[27][2] ,
         \mult_19/SUMB[27][3] , \mult_19/SUMB[27][4] , \mult_19/SUMB[27][5] ,
         \mult_19/SUMB[27][6] , \mult_19/SUMB[27][7] , \mult_19/SUMB[27][8] ,
         \mult_19/SUMB[27][9] , \mult_19/SUMB[27][10] , \mult_19/SUMB[27][11] ,
         \mult_19/SUMB[27][12] , \mult_19/SUMB[27][13] ,
         \mult_19/SUMB[27][14] , \mult_19/SUMB[27][15] ,
         \mult_19/SUMB[27][16] , \mult_19/SUMB[27][17] ,
         \mult_19/SUMB[27][18] , \mult_19/SUMB[27][19] ,
         \mult_19/SUMB[27][20] , \mult_19/SUMB[27][21] ,
         \mult_19/SUMB[27][22] , \mult_19/SUMB[27][23] ,
         \mult_19/SUMB[27][24] , \mult_19/SUMB[27][25] ,
         \mult_19/SUMB[27][26] , \mult_19/SUMB[27][27] ,
         \mult_19/SUMB[27][28] , \mult_19/SUMB[27][29] ,
         \mult_19/SUMB[27][30] , \mult_19/SUMB[28][1] , \mult_19/SUMB[28][2] ,
         \mult_19/SUMB[28][3] , \mult_19/SUMB[28][4] , \mult_19/SUMB[28][5] ,
         \mult_19/SUMB[28][6] , \mult_19/SUMB[28][7] , \mult_19/SUMB[28][8] ,
         \mult_19/SUMB[28][9] , \mult_19/SUMB[28][10] , \mult_19/SUMB[28][11] ,
         \mult_19/SUMB[28][12] , \mult_19/SUMB[28][13] ,
         \mult_19/SUMB[28][14] , \mult_19/SUMB[28][15] ,
         \mult_19/SUMB[28][16] , \mult_19/SUMB[28][17] ,
         \mult_19/SUMB[28][18] , \mult_19/SUMB[28][19] ,
         \mult_19/SUMB[28][20] , \mult_19/SUMB[28][21] ,
         \mult_19/SUMB[28][22] , \mult_19/SUMB[28][23] ,
         \mult_19/SUMB[28][24] , \mult_19/SUMB[28][25] ,
         \mult_19/SUMB[28][26] , \mult_19/SUMB[28][27] ,
         \mult_19/SUMB[28][28] , \mult_19/SUMB[28][29] ,
         \mult_19/SUMB[28][30] , \mult_19/SUMB[29][1] , \mult_19/SUMB[29][2] ,
         \mult_19/SUMB[29][3] , \mult_19/SUMB[29][4] , \mult_19/SUMB[29][5] ,
         \mult_19/SUMB[29][6] , \mult_19/SUMB[29][7] , \mult_19/SUMB[29][8] ,
         \mult_19/SUMB[29][9] , \mult_19/SUMB[29][10] , \mult_19/SUMB[29][11] ,
         \mult_19/SUMB[29][12] , \mult_19/SUMB[29][13] ,
         \mult_19/SUMB[29][14] , \mult_19/SUMB[29][15] ,
         \mult_19/SUMB[29][16] , \mult_19/SUMB[29][17] ,
         \mult_19/SUMB[29][18] , \mult_19/SUMB[29][19] ,
         \mult_19/SUMB[29][20] , \mult_19/SUMB[29][21] ,
         \mult_19/SUMB[29][22] , \mult_19/SUMB[29][23] ,
         \mult_19/SUMB[29][24] , \mult_19/SUMB[29][25] ,
         \mult_19/SUMB[29][26] , \mult_19/SUMB[29][27] ,
         \mult_19/SUMB[29][28] , \mult_19/SUMB[29][29] ,
         \mult_19/SUMB[29][30] , \mult_19/SUMB[30][1] , \mult_19/SUMB[30][2] ,
         \mult_19/SUMB[30][3] , \mult_19/SUMB[30][4] , \mult_19/SUMB[30][5] ,
         \mult_19/SUMB[30][6] , \mult_19/SUMB[30][7] , \mult_19/SUMB[30][8] ,
         \mult_19/SUMB[30][9] , \mult_19/SUMB[30][10] , \mult_19/SUMB[30][11] ,
         \mult_19/SUMB[30][12] , \mult_19/SUMB[30][13] ,
         \mult_19/SUMB[30][14] , \mult_19/SUMB[30][15] ,
         \mult_19/SUMB[30][16] , \mult_19/SUMB[30][17] ,
         \mult_19/SUMB[30][18] , \mult_19/SUMB[30][19] ,
         \mult_19/SUMB[30][20] , \mult_19/SUMB[30][21] ,
         \mult_19/SUMB[30][22] , \mult_19/SUMB[30][23] ,
         \mult_19/SUMB[30][24] , \mult_19/SUMB[30][25] ,
         \mult_19/SUMB[30][26] , \mult_19/SUMB[30][27] ,
         \mult_19/SUMB[30][28] , \mult_19/SUMB[30][29] ,
         \mult_19/SUMB[30][30] , \mult_19/SUMB[31][1] , \mult_19/SUMB[31][2] ,
         \mult_19/SUMB[31][3] , \mult_19/SUMB[31][4] , \mult_19/SUMB[31][5] ,
         \mult_19/SUMB[31][6] , \mult_19/SUMB[31][7] , \mult_19/SUMB[31][8] ,
         \mult_19/SUMB[31][9] , \mult_19/SUMB[31][10] , \mult_19/SUMB[31][11] ,
         \mult_19/SUMB[31][12] , \mult_19/SUMB[31][13] ,
         \mult_19/SUMB[31][14] , \mult_19/SUMB[31][15] ,
         \mult_19/SUMB[31][16] , \mult_19/SUMB[31][17] ,
         \mult_19/SUMB[31][18] , \mult_19/SUMB[31][19] ,
         \mult_19/SUMB[31][20] , \mult_19/SUMB[31][21] ,
         \mult_19/SUMB[31][22] , \mult_19/SUMB[31][23] ,
         \mult_19/SUMB[31][24] , \mult_19/SUMB[31][25] ,
         \mult_19/SUMB[31][26] , \mult_19/SUMB[31][27] ,
         \mult_19/SUMB[31][28] , \mult_19/SUMB[31][29] ,
         \mult_19/SUMB[31][30] , \mult_19/CARRYB[16][0] ,
         \mult_19/CARRYB[16][1] , \mult_19/CARRYB[16][2] ,
         \mult_19/CARRYB[16][3] , \mult_19/CARRYB[16][4] ,
         \mult_19/CARRYB[16][5] , \mult_19/CARRYB[16][6] ,
         \mult_19/CARRYB[16][7] , \mult_19/CARRYB[16][8] ,
         \mult_19/CARRYB[16][9] , \mult_19/CARRYB[16][10] ,
         \mult_19/CARRYB[16][11] , \mult_19/CARRYB[16][12] ,
         \mult_19/CARRYB[16][13] , \mult_19/CARRYB[16][14] ,
         \mult_19/CARRYB[16][15] , \mult_19/CARRYB[16][16] ,
         \mult_19/CARRYB[16][17] , \mult_19/CARRYB[16][18] ,
         \mult_19/CARRYB[16][19] , \mult_19/CARRYB[16][20] ,
         \mult_19/CARRYB[16][21] , \mult_19/CARRYB[16][22] ,
         \mult_19/CARRYB[16][23] , \mult_19/CARRYB[16][24] ,
         \mult_19/CARRYB[16][25] , \mult_19/CARRYB[16][26] ,
         \mult_19/CARRYB[16][27] , \mult_19/CARRYB[16][28] ,
         \mult_19/CARRYB[16][29] , \mult_19/CARRYB[16][30] ,
         \mult_19/CARRYB[17][0] , \mult_19/CARRYB[17][1] ,
         \mult_19/CARRYB[17][2] , \mult_19/CARRYB[17][3] ,
         \mult_19/CARRYB[17][4] , \mult_19/CARRYB[17][5] ,
         \mult_19/CARRYB[17][6] , \mult_19/CARRYB[17][7] ,
         \mult_19/CARRYB[17][8] , \mult_19/CARRYB[17][9] ,
         \mult_19/CARRYB[17][10] , \mult_19/CARRYB[17][11] ,
         \mult_19/CARRYB[17][12] , \mult_19/CARRYB[17][13] ,
         \mult_19/CARRYB[17][14] , \mult_19/CARRYB[17][15] ,
         \mult_19/CARRYB[17][16] , \mult_19/CARRYB[17][17] ,
         \mult_19/CARRYB[17][18] , \mult_19/CARRYB[17][19] ,
         \mult_19/CARRYB[17][20] , \mult_19/CARRYB[17][21] ,
         \mult_19/CARRYB[17][22] , \mult_19/CARRYB[17][23] ,
         \mult_19/CARRYB[17][24] , \mult_19/CARRYB[17][25] ,
         \mult_19/CARRYB[17][26] , \mult_19/CARRYB[17][27] ,
         \mult_19/CARRYB[17][28] , \mult_19/CARRYB[17][29] ,
         \mult_19/CARRYB[17][30] , \mult_19/CARRYB[18][0] ,
         \mult_19/CARRYB[18][1] , \mult_19/CARRYB[18][2] ,
         \mult_19/CARRYB[18][3] , \mult_19/CARRYB[18][4] ,
         \mult_19/CARRYB[18][5] , \mult_19/CARRYB[18][6] ,
         \mult_19/CARRYB[18][7] , \mult_19/CARRYB[18][8] ,
         \mult_19/CARRYB[18][9] , \mult_19/CARRYB[18][10] ,
         \mult_19/CARRYB[18][11] , \mult_19/CARRYB[18][12] ,
         \mult_19/CARRYB[18][13] , \mult_19/CARRYB[18][14] ,
         \mult_19/CARRYB[18][15] , \mult_19/CARRYB[18][16] ,
         \mult_19/CARRYB[18][17] , \mult_19/CARRYB[18][18] ,
         \mult_19/CARRYB[18][19] , \mult_19/CARRYB[18][20] ,
         \mult_19/CARRYB[18][21] , \mult_19/CARRYB[18][22] ,
         \mult_19/CARRYB[18][23] , \mult_19/CARRYB[18][24] ,
         \mult_19/CARRYB[18][25] , \mult_19/CARRYB[18][26] ,
         \mult_19/CARRYB[18][27] , \mult_19/CARRYB[18][28] ,
         \mult_19/CARRYB[18][29] , \mult_19/CARRYB[18][30] ,
         \mult_19/CARRYB[19][0] , \mult_19/CARRYB[19][1] ,
         \mult_19/CARRYB[19][2] , \mult_19/CARRYB[19][3] ,
         \mult_19/CARRYB[19][4] , \mult_19/CARRYB[19][5] ,
         \mult_19/CARRYB[19][6] , \mult_19/CARRYB[19][7] ,
         \mult_19/CARRYB[19][8] , \mult_19/CARRYB[19][9] ,
         \mult_19/CARRYB[19][10] , \mult_19/CARRYB[19][11] ,
         \mult_19/CARRYB[19][12] , \mult_19/CARRYB[19][13] ,
         \mult_19/CARRYB[19][14] , \mult_19/CARRYB[19][15] ,
         \mult_19/CARRYB[19][16] , \mult_19/CARRYB[19][17] ,
         \mult_19/CARRYB[19][18] , \mult_19/CARRYB[19][19] ,
         \mult_19/CARRYB[19][20] , \mult_19/CARRYB[19][21] ,
         \mult_19/CARRYB[19][22] , \mult_19/CARRYB[19][23] ,
         \mult_19/CARRYB[19][24] , \mult_19/CARRYB[19][25] ,
         \mult_19/CARRYB[19][26] , \mult_19/CARRYB[19][27] ,
         \mult_19/CARRYB[19][28] , \mult_19/CARRYB[19][29] ,
         \mult_19/CARRYB[19][30] , \mult_19/CARRYB[20][0] ,
         \mult_19/CARRYB[20][1] , \mult_19/CARRYB[20][2] ,
         \mult_19/CARRYB[20][3] , \mult_19/CARRYB[20][4] ,
         \mult_19/CARRYB[20][5] , \mult_19/CARRYB[20][6] ,
         \mult_19/CARRYB[20][7] , \mult_19/CARRYB[20][8] ,
         \mult_19/CARRYB[20][9] , \mult_19/CARRYB[20][10] ,
         \mult_19/CARRYB[20][11] , \mult_19/CARRYB[20][12] ,
         \mult_19/CARRYB[20][13] , \mult_19/CARRYB[20][14] ,
         \mult_19/CARRYB[20][15] , \mult_19/CARRYB[20][16] ,
         \mult_19/CARRYB[20][17] , \mult_19/CARRYB[20][18] ,
         \mult_19/CARRYB[20][19] , \mult_19/CARRYB[20][20] ,
         \mult_19/CARRYB[20][21] , \mult_19/CARRYB[20][22] ,
         \mult_19/CARRYB[20][23] , \mult_19/CARRYB[20][24] ,
         \mult_19/CARRYB[20][25] , \mult_19/CARRYB[20][26] ,
         \mult_19/CARRYB[20][27] , \mult_19/CARRYB[20][28] ,
         \mult_19/CARRYB[20][29] , \mult_19/CARRYB[20][30] ,
         \mult_19/CARRYB[21][0] , \mult_19/CARRYB[21][1] ,
         \mult_19/CARRYB[21][2] , \mult_19/CARRYB[21][3] ,
         \mult_19/CARRYB[21][4] , \mult_19/CARRYB[21][5] ,
         \mult_19/CARRYB[21][6] , \mult_19/CARRYB[21][7] ,
         \mult_19/CARRYB[21][8] , \mult_19/CARRYB[21][9] ,
         \mult_19/CARRYB[21][10] , \mult_19/CARRYB[21][11] ,
         \mult_19/CARRYB[21][12] , \mult_19/CARRYB[21][13] ,
         \mult_19/CARRYB[21][14] , \mult_19/CARRYB[21][15] ,
         \mult_19/CARRYB[21][16] , \mult_19/CARRYB[21][17] ,
         \mult_19/CARRYB[21][18] , \mult_19/CARRYB[21][19] ,
         \mult_19/CARRYB[21][20] , \mult_19/CARRYB[21][21] ,
         \mult_19/CARRYB[21][22] , \mult_19/CARRYB[21][23] ,
         \mult_19/CARRYB[21][24] , \mult_19/CARRYB[21][25] ,
         \mult_19/CARRYB[21][26] , \mult_19/CARRYB[21][27] ,
         \mult_19/CARRYB[21][28] , \mult_19/CARRYB[21][29] ,
         \mult_19/CARRYB[21][30] , \mult_19/CARRYB[22][0] ,
         \mult_19/CARRYB[22][1] , \mult_19/CARRYB[22][2] ,
         \mult_19/CARRYB[22][3] , \mult_19/CARRYB[22][4] ,
         \mult_19/CARRYB[22][5] , \mult_19/CARRYB[22][6] ,
         \mult_19/CARRYB[22][7] , \mult_19/CARRYB[22][8] ,
         \mult_19/CARRYB[22][9] , \mult_19/CARRYB[22][10] ,
         \mult_19/CARRYB[22][11] , \mult_19/CARRYB[22][12] ,
         \mult_19/CARRYB[22][13] , \mult_19/CARRYB[22][14] ,
         \mult_19/CARRYB[22][15] , \mult_19/CARRYB[22][16] ,
         \mult_19/CARRYB[22][17] , \mult_19/CARRYB[22][18] ,
         \mult_19/CARRYB[22][19] , \mult_19/CARRYB[22][20] ,
         \mult_19/CARRYB[22][21] , \mult_19/CARRYB[22][22] ,
         \mult_19/CARRYB[22][23] , \mult_19/CARRYB[22][24] ,
         \mult_19/CARRYB[22][25] , \mult_19/CARRYB[22][26] ,
         \mult_19/CARRYB[22][27] , \mult_19/CARRYB[22][28] ,
         \mult_19/CARRYB[22][29] , \mult_19/CARRYB[22][30] ,
         \mult_19/CARRYB[23][0] , \mult_19/CARRYB[23][1] ,
         \mult_19/CARRYB[23][2] , \mult_19/CARRYB[23][3] ,
         \mult_19/CARRYB[23][4] , \mult_19/CARRYB[23][5] ,
         \mult_19/CARRYB[23][6] , \mult_19/CARRYB[23][7] ,
         \mult_19/CARRYB[23][8] , \mult_19/CARRYB[23][9] ,
         \mult_19/CARRYB[23][10] , \mult_19/CARRYB[23][11] ,
         \mult_19/CARRYB[23][12] , \mult_19/CARRYB[23][13] ,
         \mult_19/CARRYB[23][14] , \mult_19/CARRYB[23][15] ,
         \mult_19/CARRYB[23][16] , \mult_19/CARRYB[23][17] ,
         \mult_19/CARRYB[23][18] , \mult_19/CARRYB[23][19] ,
         \mult_19/CARRYB[23][20] , \mult_19/CARRYB[23][21] ,
         \mult_19/CARRYB[23][22] , \mult_19/CARRYB[23][23] ,
         \mult_19/CARRYB[23][24] , \mult_19/CARRYB[23][25] ,
         \mult_19/CARRYB[23][26] , \mult_19/CARRYB[23][27] ,
         \mult_19/CARRYB[23][28] , \mult_19/CARRYB[23][29] ,
         \mult_19/CARRYB[23][30] , \mult_19/CARRYB[24][0] ,
         \mult_19/CARRYB[24][1] , \mult_19/CARRYB[24][2] ,
         \mult_19/CARRYB[24][3] , \mult_19/CARRYB[24][4] ,
         \mult_19/CARRYB[24][5] , \mult_19/CARRYB[24][6] ,
         \mult_19/CARRYB[24][7] , \mult_19/CARRYB[24][8] ,
         \mult_19/CARRYB[24][9] , \mult_19/CARRYB[24][10] ,
         \mult_19/CARRYB[24][11] , \mult_19/CARRYB[24][12] ,
         \mult_19/CARRYB[24][13] , \mult_19/CARRYB[24][14] ,
         \mult_19/CARRYB[24][15] , \mult_19/CARRYB[24][16] ,
         \mult_19/CARRYB[24][17] , \mult_19/CARRYB[24][18] ,
         \mult_19/CARRYB[24][19] , \mult_19/CARRYB[24][20] ,
         \mult_19/CARRYB[24][21] , \mult_19/CARRYB[24][22] ,
         \mult_19/CARRYB[24][23] , \mult_19/CARRYB[24][24] ,
         \mult_19/CARRYB[24][25] , \mult_19/CARRYB[24][26] ,
         \mult_19/CARRYB[24][27] , \mult_19/CARRYB[24][28] ,
         \mult_19/CARRYB[24][29] , \mult_19/CARRYB[24][30] ,
         \mult_19/CARRYB[25][0] , \mult_19/CARRYB[25][1] ,
         \mult_19/CARRYB[25][2] , \mult_19/CARRYB[25][3] ,
         \mult_19/CARRYB[25][4] , \mult_19/CARRYB[25][5] ,
         \mult_19/CARRYB[25][6] , \mult_19/CARRYB[25][7] ,
         \mult_19/CARRYB[25][8] , \mult_19/CARRYB[25][9] ,
         \mult_19/CARRYB[25][10] , \mult_19/CARRYB[25][11] ,
         \mult_19/CARRYB[25][12] , \mult_19/CARRYB[25][13] ,
         \mult_19/CARRYB[25][14] , \mult_19/CARRYB[25][15] ,
         \mult_19/CARRYB[25][16] , \mult_19/CARRYB[25][17] ,
         \mult_19/CARRYB[25][18] , \mult_19/CARRYB[25][19] ,
         \mult_19/CARRYB[25][20] , \mult_19/CARRYB[25][21] ,
         \mult_19/CARRYB[25][22] , \mult_19/CARRYB[25][23] ,
         \mult_19/CARRYB[25][24] , \mult_19/CARRYB[25][25] ,
         \mult_19/CARRYB[25][26] , \mult_19/CARRYB[25][27] ,
         \mult_19/CARRYB[25][28] , \mult_19/CARRYB[25][29] ,
         \mult_19/CARRYB[25][30] , \mult_19/CARRYB[26][0] ,
         \mult_19/CARRYB[26][1] , \mult_19/CARRYB[26][2] ,
         \mult_19/CARRYB[26][3] , \mult_19/CARRYB[26][4] ,
         \mult_19/CARRYB[26][5] , \mult_19/CARRYB[26][6] ,
         \mult_19/CARRYB[26][7] , \mult_19/CARRYB[26][8] ,
         \mult_19/CARRYB[26][9] , \mult_19/CARRYB[26][10] ,
         \mult_19/CARRYB[26][11] , \mult_19/CARRYB[26][12] ,
         \mult_19/CARRYB[26][13] , \mult_19/CARRYB[26][14] ,
         \mult_19/CARRYB[26][15] , \mult_19/CARRYB[26][16] ,
         \mult_19/CARRYB[26][17] , \mult_19/CARRYB[26][18] ,
         \mult_19/CARRYB[26][19] , \mult_19/CARRYB[26][20] ,
         \mult_19/CARRYB[26][21] , \mult_19/CARRYB[26][22] ,
         \mult_19/CARRYB[26][23] , \mult_19/CARRYB[26][24] ,
         \mult_19/CARRYB[26][25] , \mult_19/CARRYB[26][26] ,
         \mult_19/CARRYB[26][27] , \mult_19/CARRYB[26][28] ,
         \mult_19/CARRYB[26][29] , \mult_19/CARRYB[26][30] ,
         \mult_19/CARRYB[27][0] , \mult_19/CARRYB[27][1] ,
         \mult_19/CARRYB[27][2] , \mult_19/CARRYB[27][3] ,
         \mult_19/CARRYB[27][4] , \mult_19/CARRYB[27][5] ,
         \mult_19/CARRYB[27][6] , \mult_19/CARRYB[27][7] ,
         \mult_19/CARRYB[27][8] , \mult_19/CARRYB[27][9] ,
         \mult_19/CARRYB[27][10] , \mult_19/CARRYB[27][11] ,
         \mult_19/CARRYB[27][12] , \mult_19/CARRYB[27][13] ,
         \mult_19/CARRYB[27][14] , \mult_19/CARRYB[27][15] ,
         \mult_19/CARRYB[27][16] , \mult_19/CARRYB[27][17] ,
         \mult_19/CARRYB[27][18] , \mult_19/CARRYB[27][19] ,
         \mult_19/CARRYB[27][20] , \mult_19/CARRYB[27][21] ,
         \mult_19/CARRYB[27][22] , \mult_19/CARRYB[27][23] ,
         \mult_19/CARRYB[27][24] , \mult_19/CARRYB[27][25] ,
         \mult_19/CARRYB[27][26] , \mult_19/CARRYB[27][27] ,
         \mult_19/CARRYB[27][28] , \mult_19/CARRYB[27][29] ,
         \mult_19/CARRYB[27][30] , \mult_19/CARRYB[28][0] ,
         \mult_19/CARRYB[28][1] , \mult_19/CARRYB[28][2] ,
         \mult_19/CARRYB[28][3] , \mult_19/CARRYB[28][4] ,
         \mult_19/CARRYB[28][5] , \mult_19/CARRYB[28][6] ,
         \mult_19/CARRYB[28][7] , \mult_19/CARRYB[28][8] ,
         \mult_19/CARRYB[28][9] , \mult_19/CARRYB[28][10] ,
         \mult_19/CARRYB[28][11] , \mult_19/CARRYB[28][12] ,
         \mult_19/CARRYB[28][13] , \mult_19/CARRYB[28][14] ,
         \mult_19/CARRYB[28][15] , \mult_19/CARRYB[28][16] ,
         \mult_19/CARRYB[28][17] , \mult_19/CARRYB[28][18] ,
         \mult_19/CARRYB[28][19] , \mult_19/CARRYB[28][20] ,
         \mult_19/CARRYB[28][21] , \mult_19/CARRYB[28][22] ,
         \mult_19/CARRYB[28][23] , \mult_19/CARRYB[28][24] ,
         \mult_19/CARRYB[28][25] , \mult_19/CARRYB[28][26] ,
         \mult_19/CARRYB[28][27] , \mult_19/CARRYB[28][28] ,
         \mult_19/CARRYB[28][29] , \mult_19/CARRYB[28][30] ,
         \mult_19/CARRYB[29][0] , \mult_19/CARRYB[29][1] ,
         \mult_19/CARRYB[29][2] , \mult_19/CARRYB[29][3] ,
         \mult_19/CARRYB[29][4] , \mult_19/CARRYB[29][5] ,
         \mult_19/CARRYB[29][6] , \mult_19/CARRYB[29][7] ,
         \mult_19/CARRYB[29][8] , \mult_19/CARRYB[29][9] ,
         \mult_19/CARRYB[29][10] , \mult_19/CARRYB[29][11] ,
         \mult_19/CARRYB[29][12] , \mult_19/CARRYB[29][13] ,
         \mult_19/CARRYB[29][14] , \mult_19/CARRYB[29][15] ,
         \mult_19/CARRYB[29][16] , \mult_19/CARRYB[29][17] ,
         \mult_19/CARRYB[29][18] , \mult_19/CARRYB[29][19] ,
         \mult_19/CARRYB[29][20] , \mult_19/CARRYB[29][21] ,
         \mult_19/CARRYB[29][22] , \mult_19/CARRYB[29][23] ,
         \mult_19/CARRYB[29][24] , \mult_19/CARRYB[29][25] ,
         \mult_19/CARRYB[29][26] , \mult_19/CARRYB[29][27] ,
         \mult_19/CARRYB[29][28] , \mult_19/CARRYB[29][29] ,
         \mult_19/CARRYB[29][30] , \mult_19/CARRYB[30][0] ,
         \mult_19/CARRYB[30][1] , \mult_19/CARRYB[30][2] ,
         \mult_19/CARRYB[30][3] , \mult_19/CARRYB[30][4] ,
         \mult_19/CARRYB[30][5] , \mult_19/CARRYB[30][6] ,
         \mult_19/CARRYB[30][7] , \mult_19/CARRYB[30][8] ,
         \mult_19/CARRYB[30][9] , \mult_19/CARRYB[30][10] ,
         \mult_19/CARRYB[30][11] , \mult_19/CARRYB[30][12] ,
         \mult_19/CARRYB[30][13] , \mult_19/CARRYB[30][14] ,
         \mult_19/CARRYB[30][15] , \mult_19/CARRYB[30][16] ,
         \mult_19/CARRYB[30][17] , \mult_19/CARRYB[30][18] ,
         \mult_19/CARRYB[30][19] , \mult_19/CARRYB[30][20] ,
         \mult_19/CARRYB[30][21] , \mult_19/CARRYB[30][22] ,
         \mult_19/CARRYB[30][23] , \mult_19/CARRYB[30][24] ,
         \mult_19/CARRYB[30][25] , \mult_19/CARRYB[30][26] ,
         \mult_19/CARRYB[30][27] , \mult_19/CARRYB[30][28] ,
         \mult_19/CARRYB[30][29] , \mult_19/CARRYB[30][30] ,
         \mult_19/CARRYB[31][0] , \mult_19/CARRYB[31][1] ,
         \mult_19/CARRYB[31][2] , \mult_19/CARRYB[31][3] ,
         \mult_19/CARRYB[31][4] , \mult_19/CARRYB[31][5] ,
         \mult_19/CARRYB[31][6] , \mult_19/CARRYB[31][7] ,
         \mult_19/CARRYB[31][8] , \mult_19/CARRYB[31][9] ,
         \mult_19/CARRYB[31][10] , \mult_19/CARRYB[31][11] ,
         \mult_19/CARRYB[31][12] , \mult_19/CARRYB[31][13] ,
         \mult_19/CARRYB[31][14] , \mult_19/CARRYB[31][15] ,
         \mult_19/CARRYB[31][16] , \mult_19/CARRYB[31][17] ,
         \mult_19/CARRYB[31][18] , \mult_19/CARRYB[31][19] ,
         \mult_19/CARRYB[31][20] , \mult_19/CARRYB[31][21] ,
         \mult_19/CARRYB[31][22] , \mult_19/CARRYB[31][23] ,
         \mult_19/CARRYB[31][24] , \mult_19/CARRYB[31][25] ,
         \mult_19/CARRYB[31][26] , \mult_19/CARRYB[31][27] ,
         \mult_19/CARRYB[31][28] , \mult_19/CARRYB[31][29] ,
         \mult_19/CARRYB[31][30] , \mult_19/SUMB[2][1] , \mult_19/SUMB[2][2] ,
         \mult_19/SUMB[2][3] , \mult_19/SUMB[2][4] , \mult_19/SUMB[2][5] ,
         \mult_19/SUMB[2][6] , \mult_19/SUMB[2][7] , \mult_19/SUMB[2][8] ,
         \mult_19/SUMB[2][9] , \mult_19/SUMB[2][10] , \mult_19/SUMB[2][11] ,
         \mult_19/SUMB[2][12] , \mult_19/SUMB[2][13] , \mult_19/SUMB[2][14] ,
         \mult_19/SUMB[2][15] , \mult_19/SUMB[2][16] , \mult_19/SUMB[2][17] ,
         \mult_19/SUMB[2][18] , \mult_19/SUMB[2][19] , \mult_19/SUMB[2][20] ,
         \mult_19/SUMB[2][21] , \mult_19/SUMB[2][22] , \mult_19/SUMB[2][23] ,
         \mult_19/SUMB[2][24] , \mult_19/SUMB[2][25] , \mult_19/SUMB[2][26] ,
         \mult_19/SUMB[2][27] , \mult_19/SUMB[2][28] , \mult_19/SUMB[2][29] ,
         \mult_19/SUMB[2][30] , \mult_19/SUMB[3][1] , \mult_19/SUMB[3][2] ,
         \mult_19/SUMB[3][3] , \mult_19/SUMB[3][4] , \mult_19/SUMB[3][5] ,
         \mult_19/SUMB[3][6] , \mult_19/SUMB[3][7] , \mult_19/SUMB[3][8] ,
         \mult_19/SUMB[3][9] , \mult_19/SUMB[3][10] , \mult_19/SUMB[3][11] ,
         \mult_19/SUMB[3][12] , \mult_19/SUMB[3][13] , \mult_19/SUMB[3][14] ,
         \mult_19/SUMB[3][15] , \mult_19/SUMB[3][16] , \mult_19/SUMB[3][17] ,
         \mult_19/SUMB[3][18] , \mult_19/SUMB[3][19] , \mult_19/SUMB[3][20] ,
         \mult_19/SUMB[3][21] , \mult_19/SUMB[3][22] , \mult_19/SUMB[3][23] ,
         \mult_19/SUMB[3][24] , \mult_19/SUMB[3][25] , \mult_19/SUMB[3][26] ,
         \mult_19/SUMB[3][27] , \mult_19/SUMB[3][28] , \mult_19/SUMB[3][29] ,
         \mult_19/SUMB[3][30] , \mult_19/SUMB[4][1] , \mult_19/SUMB[4][2] ,
         \mult_19/SUMB[4][3] , \mult_19/SUMB[4][4] , \mult_19/SUMB[4][5] ,
         \mult_19/SUMB[4][6] , \mult_19/SUMB[4][7] , \mult_19/SUMB[4][8] ,
         \mult_19/SUMB[4][9] , \mult_19/SUMB[4][10] , \mult_19/SUMB[4][11] ,
         \mult_19/SUMB[4][12] , \mult_19/SUMB[4][13] , \mult_19/SUMB[4][14] ,
         \mult_19/SUMB[4][15] , \mult_19/SUMB[4][16] , \mult_19/SUMB[4][17] ,
         \mult_19/SUMB[4][18] , \mult_19/SUMB[4][19] , \mult_19/SUMB[4][20] ,
         \mult_19/SUMB[4][21] , \mult_19/SUMB[4][22] , \mult_19/SUMB[4][23] ,
         \mult_19/SUMB[4][24] , \mult_19/SUMB[4][25] , \mult_19/SUMB[4][26] ,
         \mult_19/SUMB[4][27] , \mult_19/SUMB[4][28] , \mult_19/SUMB[4][29] ,
         \mult_19/SUMB[4][30] , \mult_19/SUMB[5][1] , \mult_19/SUMB[5][2] ,
         \mult_19/SUMB[5][3] , \mult_19/SUMB[5][4] , \mult_19/SUMB[5][5] ,
         \mult_19/SUMB[5][6] , \mult_19/SUMB[5][7] , \mult_19/SUMB[5][8] ,
         \mult_19/SUMB[5][9] , \mult_19/SUMB[5][10] , \mult_19/SUMB[5][11] ,
         \mult_19/SUMB[5][12] , \mult_19/SUMB[5][13] , \mult_19/SUMB[5][14] ,
         \mult_19/SUMB[5][15] , \mult_19/SUMB[5][16] , \mult_19/SUMB[5][17] ,
         \mult_19/SUMB[5][18] , \mult_19/SUMB[5][19] , \mult_19/SUMB[5][20] ,
         \mult_19/SUMB[5][21] , \mult_19/SUMB[5][22] , \mult_19/SUMB[5][23] ,
         \mult_19/SUMB[5][24] , \mult_19/SUMB[5][25] , \mult_19/SUMB[5][26] ,
         \mult_19/SUMB[5][27] , \mult_19/SUMB[5][28] , \mult_19/SUMB[5][29] ,
         \mult_19/SUMB[5][30] , \mult_19/SUMB[6][1] , \mult_19/SUMB[6][2] ,
         \mult_19/SUMB[6][3] , \mult_19/SUMB[6][4] , \mult_19/SUMB[6][5] ,
         \mult_19/SUMB[6][6] , \mult_19/SUMB[6][7] , \mult_19/SUMB[6][8] ,
         \mult_19/SUMB[6][9] , \mult_19/SUMB[6][10] , \mult_19/SUMB[6][11] ,
         \mult_19/SUMB[6][12] , \mult_19/SUMB[6][13] , \mult_19/SUMB[6][14] ,
         \mult_19/SUMB[6][15] , \mult_19/SUMB[6][16] , \mult_19/SUMB[6][17] ,
         \mult_19/SUMB[6][18] , \mult_19/SUMB[6][19] , \mult_19/SUMB[6][20] ,
         \mult_19/SUMB[6][21] , \mult_19/SUMB[6][22] , \mult_19/SUMB[6][23] ,
         \mult_19/SUMB[6][24] , \mult_19/SUMB[6][25] , \mult_19/SUMB[6][26] ,
         \mult_19/SUMB[6][27] , \mult_19/SUMB[6][28] , \mult_19/SUMB[6][29] ,
         \mult_19/SUMB[6][30] , \mult_19/SUMB[7][1] , \mult_19/SUMB[7][2] ,
         \mult_19/SUMB[7][3] , \mult_19/SUMB[7][4] , \mult_19/SUMB[7][5] ,
         \mult_19/SUMB[7][6] , \mult_19/SUMB[7][7] , \mult_19/SUMB[7][8] ,
         \mult_19/SUMB[7][9] , \mult_19/SUMB[7][10] , \mult_19/SUMB[7][11] ,
         \mult_19/SUMB[7][12] , \mult_19/SUMB[7][13] , \mult_19/SUMB[7][14] ,
         \mult_19/SUMB[7][15] , \mult_19/SUMB[7][16] , \mult_19/SUMB[7][17] ,
         \mult_19/SUMB[7][18] , \mult_19/SUMB[7][19] , \mult_19/SUMB[7][20] ,
         \mult_19/SUMB[7][21] , \mult_19/SUMB[7][22] , \mult_19/SUMB[7][23] ,
         \mult_19/SUMB[7][24] , \mult_19/SUMB[7][25] , \mult_19/SUMB[7][26] ,
         \mult_19/SUMB[7][27] , \mult_19/SUMB[7][28] , \mult_19/SUMB[7][29] ,
         \mult_19/SUMB[7][30] , \mult_19/SUMB[8][1] , \mult_19/SUMB[8][2] ,
         \mult_19/SUMB[8][3] , \mult_19/SUMB[8][4] , \mult_19/SUMB[8][5] ,
         \mult_19/SUMB[8][6] , \mult_19/SUMB[8][7] , \mult_19/SUMB[8][8] ,
         \mult_19/SUMB[8][9] , \mult_19/SUMB[8][10] , \mult_19/SUMB[8][11] ,
         \mult_19/SUMB[8][12] , \mult_19/SUMB[8][13] , \mult_19/SUMB[8][14] ,
         \mult_19/SUMB[8][15] , \mult_19/SUMB[8][16] , \mult_19/SUMB[8][17] ,
         \mult_19/SUMB[8][18] , \mult_19/SUMB[8][19] , \mult_19/SUMB[8][20] ,
         \mult_19/SUMB[8][21] , \mult_19/SUMB[8][22] , \mult_19/SUMB[8][23] ,
         \mult_19/SUMB[8][24] , \mult_19/SUMB[8][25] , \mult_19/SUMB[8][26] ,
         \mult_19/SUMB[8][27] , \mult_19/SUMB[8][28] , \mult_19/SUMB[8][29] ,
         \mult_19/SUMB[8][30] , \mult_19/SUMB[9][1] , \mult_19/SUMB[9][2] ,
         \mult_19/SUMB[9][3] , \mult_19/SUMB[9][4] , \mult_19/SUMB[9][5] ,
         \mult_19/SUMB[9][6] , \mult_19/SUMB[9][7] , \mult_19/SUMB[9][8] ,
         \mult_19/SUMB[9][9] , \mult_19/SUMB[9][10] , \mult_19/SUMB[9][11] ,
         \mult_19/SUMB[9][12] , \mult_19/SUMB[9][13] , \mult_19/SUMB[9][14] ,
         \mult_19/SUMB[9][15] , \mult_19/SUMB[9][16] , \mult_19/SUMB[9][17] ,
         \mult_19/SUMB[9][18] , \mult_19/SUMB[9][19] , \mult_19/SUMB[9][20] ,
         \mult_19/SUMB[9][21] , \mult_19/SUMB[9][22] , \mult_19/SUMB[9][23] ,
         \mult_19/SUMB[9][24] , \mult_19/SUMB[9][25] , \mult_19/SUMB[9][26] ,
         \mult_19/SUMB[9][27] , \mult_19/SUMB[9][28] , \mult_19/SUMB[9][29] ,
         \mult_19/SUMB[9][30] , \mult_19/SUMB[10][1] , \mult_19/SUMB[10][2] ,
         \mult_19/SUMB[10][3] , \mult_19/SUMB[10][4] , \mult_19/SUMB[10][5] ,
         \mult_19/SUMB[10][6] , \mult_19/SUMB[10][7] , \mult_19/SUMB[10][8] ,
         \mult_19/SUMB[10][9] , \mult_19/SUMB[10][10] , \mult_19/SUMB[10][11] ,
         \mult_19/SUMB[10][12] , \mult_19/SUMB[10][13] ,
         \mult_19/SUMB[10][14] , \mult_19/SUMB[10][15] ,
         \mult_19/SUMB[10][16] , \mult_19/SUMB[10][17] ,
         \mult_19/SUMB[10][18] , \mult_19/SUMB[10][19] ,
         \mult_19/SUMB[10][20] , \mult_19/SUMB[10][21] ,
         \mult_19/SUMB[10][22] , \mult_19/SUMB[10][23] ,
         \mult_19/SUMB[10][24] , \mult_19/SUMB[10][25] ,
         \mult_19/SUMB[10][26] , \mult_19/SUMB[10][27] ,
         \mult_19/SUMB[10][28] , \mult_19/SUMB[10][29] ,
         \mult_19/SUMB[10][30] , \mult_19/SUMB[11][1] , \mult_19/SUMB[11][2] ,
         \mult_19/SUMB[11][3] , \mult_19/SUMB[11][4] , \mult_19/SUMB[11][5] ,
         \mult_19/SUMB[11][6] , \mult_19/SUMB[11][7] , \mult_19/SUMB[11][8] ,
         \mult_19/SUMB[11][9] , \mult_19/SUMB[11][10] , \mult_19/SUMB[11][11] ,
         \mult_19/SUMB[11][12] , \mult_19/SUMB[11][13] ,
         \mult_19/SUMB[11][14] , \mult_19/SUMB[11][15] ,
         \mult_19/SUMB[11][16] , \mult_19/SUMB[11][17] ,
         \mult_19/SUMB[11][18] , \mult_19/SUMB[11][19] ,
         \mult_19/SUMB[11][20] , \mult_19/SUMB[11][21] ,
         \mult_19/SUMB[11][22] , \mult_19/SUMB[11][23] ,
         \mult_19/SUMB[11][24] , \mult_19/SUMB[11][25] ,
         \mult_19/SUMB[11][26] , \mult_19/SUMB[11][27] ,
         \mult_19/SUMB[11][28] , \mult_19/SUMB[11][29] ,
         \mult_19/SUMB[11][30] , \mult_19/SUMB[12][1] , \mult_19/SUMB[12][2] ,
         \mult_19/SUMB[12][3] , \mult_19/SUMB[12][4] , \mult_19/SUMB[12][5] ,
         \mult_19/SUMB[12][6] , \mult_19/SUMB[12][7] , \mult_19/SUMB[12][8] ,
         \mult_19/SUMB[12][9] , \mult_19/SUMB[12][10] , \mult_19/SUMB[12][11] ,
         \mult_19/SUMB[12][12] , \mult_19/SUMB[12][13] ,
         \mult_19/SUMB[12][14] , \mult_19/SUMB[12][15] ,
         \mult_19/SUMB[12][16] , \mult_19/SUMB[12][17] ,
         \mult_19/SUMB[12][18] , \mult_19/SUMB[12][19] ,
         \mult_19/SUMB[12][20] , \mult_19/SUMB[12][21] ,
         \mult_19/SUMB[12][22] , \mult_19/SUMB[12][23] ,
         \mult_19/SUMB[12][24] , \mult_19/SUMB[12][25] ,
         \mult_19/SUMB[12][26] , \mult_19/SUMB[12][27] ,
         \mult_19/SUMB[12][28] , \mult_19/SUMB[12][29] ,
         \mult_19/SUMB[12][30] , \mult_19/SUMB[13][1] , \mult_19/SUMB[13][2] ,
         \mult_19/SUMB[13][3] , \mult_19/SUMB[13][4] , \mult_19/SUMB[13][5] ,
         \mult_19/SUMB[13][6] , \mult_19/SUMB[13][7] , \mult_19/SUMB[13][8] ,
         \mult_19/SUMB[13][9] , \mult_19/SUMB[13][10] , \mult_19/SUMB[13][11] ,
         \mult_19/SUMB[13][12] , \mult_19/SUMB[13][13] ,
         \mult_19/SUMB[13][14] , \mult_19/SUMB[13][15] ,
         \mult_19/SUMB[13][16] , \mult_19/SUMB[13][17] ,
         \mult_19/SUMB[13][18] , \mult_19/SUMB[13][19] ,
         \mult_19/SUMB[13][20] , \mult_19/SUMB[13][21] ,
         \mult_19/SUMB[13][22] , \mult_19/SUMB[13][23] ,
         \mult_19/SUMB[13][24] , \mult_19/SUMB[13][25] ,
         \mult_19/SUMB[13][26] , \mult_19/SUMB[13][27] ,
         \mult_19/SUMB[13][28] , \mult_19/SUMB[13][29] ,
         \mult_19/SUMB[13][30] , \mult_19/SUMB[14][1] , \mult_19/SUMB[14][2] ,
         \mult_19/SUMB[14][3] , \mult_19/SUMB[14][4] , \mult_19/SUMB[14][5] ,
         \mult_19/SUMB[14][6] , \mult_19/SUMB[14][7] , \mult_19/SUMB[14][8] ,
         \mult_19/SUMB[14][9] , \mult_19/SUMB[14][10] , \mult_19/SUMB[14][11] ,
         \mult_19/SUMB[14][12] , \mult_19/SUMB[14][13] ,
         \mult_19/SUMB[14][14] , \mult_19/SUMB[14][15] ,
         \mult_19/SUMB[14][16] , \mult_19/SUMB[14][17] ,
         \mult_19/SUMB[14][18] , \mult_19/SUMB[14][19] ,
         \mult_19/SUMB[14][20] , \mult_19/SUMB[14][21] ,
         \mult_19/SUMB[14][22] , \mult_19/SUMB[14][23] ,
         \mult_19/SUMB[14][24] , \mult_19/SUMB[14][25] ,
         \mult_19/SUMB[14][26] , \mult_19/SUMB[14][27] ,
         \mult_19/SUMB[14][28] , \mult_19/SUMB[14][29] ,
         \mult_19/SUMB[14][30] , \mult_19/SUMB[15][1] , \mult_19/SUMB[15][2] ,
         \mult_19/SUMB[15][3] , \mult_19/SUMB[15][4] , \mult_19/SUMB[15][5] ,
         \mult_19/SUMB[15][6] , \mult_19/SUMB[15][7] , \mult_19/SUMB[15][8] ,
         \mult_19/SUMB[15][9] , \mult_19/SUMB[15][10] , \mult_19/SUMB[15][11] ,
         \mult_19/SUMB[15][12] , \mult_19/SUMB[15][13] ,
         \mult_19/SUMB[15][14] , \mult_19/SUMB[15][15] ,
         \mult_19/SUMB[15][16] , \mult_19/SUMB[15][17] ,
         \mult_19/SUMB[15][18] , \mult_19/SUMB[15][19] ,
         \mult_19/SUMB[15][20] , \mult_19/SUMB[15][21] ,
         \mult_19/SUMB[15][22] , \mult_19/SUMB[15][23] ,
         \mult_19/SUMB[15][24] , \mult_19/SUMB[15][25] ,
         \mult_19/SUMB[15][26] , \mult_19/SUMB[15][27] ,
         \mult_19/SUMB[15][28] , \mult_19/SUMB[15][29] ,
         \mult_19/SUMB[15][30] , \mult_19/CARRYB[2][0] ,
         \mult_19/CARRYB[2][1] , \mult_19/CARRYB[2][2] ,
         \mult_19/CARRYB[2][3] , \mult_19/CARRYB[2][4] ,
         \mult_19/CARRYB[2][5] , \mult_19/CARRYB[2][6] ,
         \mult_19/CARRYB[2][7] , \mult_19/CARRYB[2][8] ,
         \mult_19/CARRYB[2][9] , \mult_19/CARRYB[2][10] ,
         \mult_19/CARRYB[2][11] , \mult_19/CARRYB[2][12] ,
         \mult_19/CARRYB[2][13] , \mult_19/CARRYB[2][14] ,
         \mult_19/CARRYB[2][15] , \mult_19/CARRYB[2][16] ,
         \mult_19/CARRYB[2][17] , \mult_19/CARRYB[2][18] ,
         \mult_19/CARRYB[2][19] , \mult_19/CARRYB[2][20] ,
         \mult_19/CARRYB[2][21] , \mult_19/CARRYB[2][22] ,
         \mult_19/CARRYB[2][23] , \mult_19/CARRYB[2][24] ,
         \mult_19/CARRYB[2][25] , \mult_19/CARRYB[2][26] ,
         \mult_19/CARRYB[2][27] , \mult_19/CARRYB[2][28] ,
         \mult_19/CARRYB[2][29] , \mult_19/CARRYB[2][30] ,
         \mult_19/CARRYB[3][0] , \mult_19/CARRYB[3][1] ,
         \mult_19/CARRYB[3][2] , \mult_19/CARRYB[3][3] ,
         \mult_19/CARRYB[3][4] , \mult_19/CARRYB[3][5] ,
         \mult_19/CARRYB[3][6] , \mult_19/CARRYB[3][7] ,
         \mult_19/CARRYB[3][8] , \mult_19/CARRYB[3][9] ,
         \mult_19/CARRYB[3][10] , \mult_19/CARRYB[3][11] ,
         \mult_19/CARRYB[3][12] , \mult_19/CARRYB[3][13] ,
         \mult_19/CARRYB[3][14] , \mult_19/CARRYB[3][15] ,
         \mult_19/CARRYB[3][16] , \mult_19/CARRYB[3][17] ,
         \mult_19/CARRYB[3][18] , \mult_19/CARRYB[3][19] ,
         \mult_19/CARRYB[3][20] , \mult_19/CARRYB[3][21] ,
         \mult_19/CARRYB[3][22] , \mult_19/CARRYB[3][23] ,
         \mult_19/CARRYB[3][24] , \mult_19/CARRYB[3][25] ,
         \mult_19/CARRYB[3][26] , \mult_19/CARRYB[3][27] ,
         \mult_19/CARRYB[3][28] , \mult_19/CARRYB[3][29] ,
         \mult_19/CARRYB[3][30] , \mult_19/CARRYB[4][0] ,
         \mult_19/CARRYB[4][1] , \mult_19/CARRYB[4][2] ,
         \mult_19/CARRYB[4][3] , \mult_19/CARRYB[4][4] ,
         \mult_19/CARRYB[4][5] , \mult_19/CARRYB[4][6] ,
         \mult_19/CARRYB[4][7] , \mult_19/CARRYB[4][8] ,
         \mult_19/CARRYB[4][9] , \mult_19/CARRYB[4][10] ,
         \mult_19/CARRYB[4][11] , \mult_19/CARRYB[4][12] ,
         \mult_19/CARRYB[4][13] , \mult_19/CARRYB[4][14] ,
         \mult_19/CARRYB[4][15] , \mult_19/CARRYB[4][16] ,
         \mult_19/CARRYB[4][17] , \mult_19/CARRYB[4][18] ,
         \mult_19/CARRYB[4][19] , \mult_19/CARRYB[4][20] ,
         \mult_19/CARRYB[4][21] , \mult_19/CARRYB[4][22] ,
         \mult_19/CARRYB[4][23] , \mult_19/CARRYB[4][24] ,
         \mult_19/CARRYB[4][25] , \mult_19/CARRYB[4][26] ,
         \mult_19/CARRYB[4][27] , \mult_19/CARRYB[4][28] ,
         \mult_19/CARRYB[4][29] , \mult_19/CARRYB[4][30] ,
         \mult_19/CARRYB[5][0] , \mult_19/CARRYB[5][1] ,
         \mult_19/CARRYB[5][2] , \mult_19/CARRYB[5][3] ,
         \mult_19/CARRYB[5][4] , \mult_19/CARRYB[5][5] ,
         \mult_19/CARRYB[5][6] , \mult_19/CARRYB[5][7] ,
         \mult_19/CARRYB[5][8] , \mult_19/CARRYB[5][9] ,
         \mult_19/CARRYB[5][10] , \mult_19/CARRYB[5][11] ,
         \mult_19/CARRYB[5][12] , \mult_19/CARRYB[5][13] ,
         \mult_19/CARRYB[5][14] , \mult_19/CARRYB[5][15] ,
         \mult_19/CARRYB[5][16] , \mult_19/CARRYB[5][17] ,
         \mult_19/CARRYB[5][18] , \mult_19/CARRYB[5][19] ,
         \mult_19/CARRYB[5][20] , \mult_19/CARRYB[5][21] ,
         \mult_19/CARRYB[5][22] , \mult_19/CARRYB[5][23] ,
         \mult_19/CARRYB[5][24] , \mult_19/CARRYB[5][25] ,
         \mult_19/CARRYB[5][26] , \mult_19/CARRYB[5][27] ,
         \mult_19/CARRYB[5][28] , \mult_19/CARRYB[5][29] ,
         \mult_19/CARRYB[5][30] , \mult_19/CARRYB[6][0] ,
         \mult_19/CARRYB[6][1] , \mult_19/CARRYB[6][2] ,
         \mult_19/CARRYB[6][3] , \mult_19/CARRYB[6][4] ,
         \mult_19/CARRYB[6][5] , \mult_19/CARRYB[6][6] ,
         \mult_19/CARRYB[6][7] , \mult_19/CARRYB[6][8] ,
         \mult_19/CARRYB[6][9] , \mult_19/CARRYB[6][10] ,
         \mult_19/CARRYB[6][11] , \mult_19/CARRYB[6][12] ,
         \mult_19/CARRYB[6][13] , \mult_19/CARRYB[6][14] ,
         \mult_19/CARRYB[6][15] , \mult_19/CARRYB[6][16] ,
         \mult_19/CARRYB[6][17] , \mult_19/CARRYB[6][18] ,
         \mult_19/CARRYB[6][19] , \mult_19/CARRYB[6][20] ,
         \mult_19/CARRYB[6][21] , \mult_19/CARRYB[6][22] ,
         \mult_19/CARRYB[6][23] , \mult_19/CARRYB[6][24] ,
         \mult_19/CARRYB[6][25] , \mult_19/CARRYB[6][26] ,
         \mult_19/CARRYB[6][27] , \mult_19/CARRYB[6][28] ,
         \mult_19/CARRYB[6][29] , \mult_19/CARRYB[6][30] ,
         \mult_19/CARRYB[7][0] , \mult_19/CARRYB[7][1] ,
         \mult_19/CARRYB[7][2] , \mult_19/CARRYB[7][3] ,
         \mult_19/CARRYB[7][4] , \mult_19/CARRYB[7][5] ,
         \mult_19/CARRYB[7][6] , \mult_19/CARRYB[7][7] ,
         \mult_19/CARRYB[7][8] , \mult_19/CARRYB[7][9] ,
         \mult_19/CARRYB[7][10] , \mult_19/CARRYB[7][11] ,
         \mult_19/CARRYB[7][12] , \mult_19/CARRYB[7][13] ,
         \mult_19/CARRYB[7][14] , \mult_19/CARRYB[7][15] ,
         \mult_19/CARRYB[7][16] , \mult_19/CARRYB[7][17] ,
         \mult_19/CARRYB[7][18] , \mult_19/CARRYB[7][19] ,
         \mult_19/CARRYB[7][20] , \mult_19/CARRYB[7][21] ,
         \mult_19/CARRYB[7][22] , \mult_19/CARRYB[7][23] ,
         \mult_19/CARRYB[7][24] , \mult_19/CARRYB[7][25] ,
         \mult_19/CARRYB[7][26] , \mult_19/CARRYB[7][27] ,
         \mult_19/CARRYB[7][28] , \mult_19/CARRYB[7][29] ,
         \mult_19/CARRYB[7][30] , \mult_19/CARRYB[8][0] ,
         \mult_19/CARRYB[8][1] , \mult_19/CARRYB[8][2] ,
         \mult_19/CARRYB[8][3] , \mult_19/CARRYB[8][4] ,
         \mult_19/CARRYB[8][5] , \mult_19/CARRYB[8][6] ,
         \mult_19/CARRYB[8][7] , \mult_19/CARRYB[8][8] ,
         \mult_19/CARRYB[8][9] , \mult_19/CARRYB[8][10] ,
         \mult_19/CARRYB[8][11] , \mult_19/CARRYB[8][12] ,
         \mult_19/CARRYB[8][13] , \mult_19/CARRYB[8][14] ,
         \mult_19/CARRYB[8][15] , \mult_19/CARRYB[8][16] ,
         \mult_19/CARRYB[8][17] , \mult_19/CARRYB[8][18] ,
         \mult_19/CARRYB[8][19] , \mult_19/CARRYB[8][20] ,
         \mult_19/CARRYB[8][21] , \mult_19/CARRYB[8][22] ,
         \mult_19/CARRYB[8][23] , \mult_19/CARRYB[8][24] ,
         \mult_19/CARRYB[8][25] , \mult_19/CARRYB[8][26] ,
         \mult_19/CARRYB[8][27] , \mult_19/CARRYB[8][28] ,
         \mult_19/CARRYB[8][29] , \mult_19/CARRYB[8][30] ,
         \mult_19/CARRYB[9][0] , \mult_19/CARRYB[9][1] ,
         \mult_19/CARRYB[9][2] , \mult_19/CARRYB[9][3] ,
         \mult_19/CARRYB[9][4] , \mult_19/CARRYB[9][5] ,
         \mult_19/CARRYB[9][6] , \mult_19/CARRYB[9][7] ,
         \mult_19/CARRYB[9][8] , \mult_19/CARRYB[9][9] ,
         \mult_19/CARRYB[9][10] , \mult_19/CARRYB[9][11] ,
         \mult_19/CARRYB[9][12] , \mult_19/CARRYB[9][13] ,
         \mult_19/CARRYB[9][14] , \mult_19/CARRYB[9][15] ,
         \mult_19/CARRYB[9][16] , \mult_19/CARRYB[9][17] ,
         \mult_19/CARRYB[9][18] , \mult_19/CARRYB[9][19] ,
         \mult_19/CARRYB[9][20] , \mult_19/CARRYB[9][21] ,
         \mult_19/CARRYB[9][22] , \mult_19/CARRYB[9][23] ,
         \mult_19/CARRYB[9][24] , \mult_19/CARRYB[9][25] ,
         \mult_19/CARRYB[9][26] , \mult_19/CARRYB[9][27] ,
         \mult_19/CARRYB[9][28] , \mult_19/CARRYB[9][29] ,
         \mult_19/CARRYB[9][30] , \mult_19/CARRYB[10][0] ,
         \mult_19/CARRYB[10][1] , \mult_19/CARRYB[10][2] ,
         \mult_19/CARRYB[10][3] , \mult_19/CARRYB[10][4] ,
         \mult_19/CARRYB[10][5] , \mult_19/CARRYB[10][6] ,
         \mult_19/CARRYB[10][7] , \mult_19/CARRYB[10][8] ,
         \mult_19/CARRYB[10][9] , \mult_19/CARRYB[10][10] ,
         \mult_19/CARRYB[10][11] , \mult_19/CARRYB[10][12] ,
         \mult_19/CARRYB[10][13] , \mult_19/CARRYB[10][14] ,
         \mult_19/CARRYB[10][15] , \mult_19/CARRYB[10][16] ,
         \mult_19/CARRYB[10][17] , \mult_19/CARRYB[10][18] ,
         \mult_19/CARRYB[10][19] , \mult_19/CARRYB[10][20] ,
         \mult_19/CARRYB[10][21] , \mult_19/CARRYB[10][22] ,
         \mult_19/CARRYB[10][23] , \mult_19/CARRYB[10][24] ,
         \mult_19/CARRYB[10][25] , \mult_19/CARRYB[10][26] ,
         \mult_19/CARRYB[10][27] , \mult_19/CARRYB[10][28] ,
         \mult_19/CARRYB[10][29] , \mult_19/CARRYB[10][30] ,
         \mult_19/CARRYB[11][0] , \mult_19/CARRYB[11][1] ,
         \mult_19/CARRYB[11][2] , \mult_19/CARRYB[11][3] ,
         \mult_19/CARRYB[11][4] , \mult_19/CARRYB[11][5] ,
         \mult_19/CARRYB[11][6] , \mult_19/CARRYB[11][7] ,
         \mult_19/CARRYB[11][8] , \mult_19/CARRYB[11][9] ,
         \mult_19/CARRYB[11][10] , \mult_19/CARRYB[11][11] ,
         \mult_19/CARRYB[11][12] , \mult_19/CARRYB[11][13] ,
         \mult_19/CARRYB[11][14] , \mult_19/CARRYB[11][15] ,
         \mult_19/CARRYB[11][16] , \mult_19/CARRYB[11][17] ,
         \mult_19/CARRYB[11][18] , \mult_19/CARRYB[11][19] ,
         \mult_19/CARRYB[11][20] , \mult_19/CARRYB[11][21] ,
         \mult_19/CARRYB[11][22] , \mult_19/CARRYB[11][23] ,
         \mult_19/CARRYB[11][24] , \mult_19/CARRYB[11][25] ,
         \mult_19/CARRYB[11][26] , \mult_19/CARRYB[11][27] ,
         \mult_19/CARRYB[11][28] , \mult_19/CARRYB[11][29] ,
         \mult_19/CARRYB[11][30] , \mult_19/CARRYB[12][0] ,
         \mult_19/CARRYB[12][1] , \mult_19/CARRYB[12][2] ,
         \mult_19/CARRYB[12][3] , \mult_19/CARRYB[12][4] ,
         \mult_19/CARRYB[12][5] , \mult_19/CARRYB[12][6] ,
         \mult_19/CARRYB[12][7] , \mult_19/CARRYB[12][8] ,
         \mult_19/CARRYB[12][9] , \mult_19/CARRYB[12][10] ,
         \mult_19/CARRYB[12][11] , \mult_19/CARRYB[12][12] ,
         \mult_19/CARRYB[12][13] , \mult_19/CARRYB[12][14] ,
         \mult_19/CARRYB[12][15] , \mult_19/CARRYB[12][16] ,
         \mult_19/CARRYB[12][17] , \mult_19/CARRYB[12][18] ,
         \mult_19/CARRYB[12][19] , \mult_19/CARRYB[12][20] ,
         \mult_19/CARRYB[12][21] , \mult_19/CARRYB[12][22] ,
         \mult_19/CARRYB[12][23] , \mult_19/CARRYB[12][24] ,
         \mult_19/CARRYB[12][25] , \mult_19/CARRYB[12][26] ,
         \mult_19/CARRYB[12][27] , \mult_19/CARRYB[12][28] ,
         \mult_19/CARRYB[12][29] , \mult_19/CARRYB[12][30] ,
         \mult_19/CARRYB[13][0] , \mult_19/CARRYB[13][1] ,
         \mult_19/CARRYB[13][2] , \mult_19/CARRYB[13][3] ,
         \mult_19/CARRYB[13][4] , \mult_19/CARRYB[13][5] ,
         \mult_19/CARRYB[13][6] , \mult_19/CARRYB[13][7] ,
         \mult_19/CARRYB[13][8] , \mult_19/CARRYB[13][9] ,
         \mult_19/CARRYB[13][10] , \mult_19/CARRYB[13][11] ,
         \mult_19/CARRYB[13][12] , \mult_19/CARRYB[13][13] ,
         \mult_19/CARRYB[13][14] , \mult_19/CARRYB[13][15] ,
         \mult_19/CARRYB[13][16] , \mult_19/CARRYB[13][17] ,
         \mult_19/CARRYB[13][18] , \mult_19/CARRYB[13][19] ,
         \mult_19/CARRYB[13][20] , \mult_19/CARRYB[13][21] ,
         \mult_19/CARRYB[13][22] , \mult_19/CARRYB[13][23] ,
         \mult_19/CARRYB[13][24] , \mult_19/CARRYB[13][25] ,
         \mult_19/CARRYB[13][26] , \mult_19/CARRYB[13][27] ,
         \mult_19/CARRYB[13][28] , \mult_19/CARRYB[13][29] ,
         \mult_19/CARRYB[13][30] , \mult_19/CARRYB[14][0] ,
         \mult_19/CARRYB[14][1] , \mult_19/CARRYB[14][2] ,
         \mult_19/CARRYB[14][3] , \mult_19/CARRYB[14][4] ,
         \mult_19/CARRYB[14][5] , \mult_19/CARRYB[14][6] ,
         \mult_19/CARRYB[14][7] , \mult_19/CARRYB[14][8] ,
         \mult_19/CARRYB[14][9] , \mult_19/CARRYB[14][10] ,
         \mult_19/CARRYB[14][11] , \mult_19/CARRYB[14][12] ,
         \mult_19/CARRYB[14][13] , \mult_19/CARRYB[14][14] ,
         \mult_19/CARRYB[14][15] , \mult_19/CARRYB[14][16] ,
         \mult_19/CARRYB[14][17] , \mult_19/CARRYB[14][18] ,
         \mult_19/CARRYB[14][19] , \mult_19/CARRYB[14][20] ,
         \mult_19/CARRYB[14][21] , \mult_19/CARRYB[14][22] ,
         \mult_19/CARRYB[14][23] , \mult_19/CARRYB[14][24] ,
         \mult_19/CARRYB[14][25] , \mult_19/CARRYB[14][26] ,
         \mult_19/CARRYB[14][27] , \mult_19/CARRYB[14][28] ,
         \mult_19/CARRYB[14][29] , \mult_19/CARRYB[14][30] ,
         \mult_19/CARRYB[15][0] , \mult_19/CARRYB[15][1] ,
         \mult_19/CARRYB[15][2] , \mult_19/CARRYB[15][3] ,
         \mult_19/CARRYB[15][4] , \mult_19/CARRYB[15][5] ,
         \mult_19/CARRYB[15][6] , \mult_19/CARRYB[15][7] ,
         \mult_19/CARRYB[15][8] , \mult_19/CARRYB[15][9] ,
         \mult_19/CARRYB[15][10] , \mult_19/CARRYB[15][11] ,
         \mult_19/CARRYB[15][12] , \mult_19/CARRYB[15][13] ,
         \mult_19/CARRYB[15][14] , \mult_19/CARRYB[15][15] ,
         \mult_19/CARRYB[15][16] , \mult_19/CARRYB[15][17] ,
         \mult_19/CARRYB[15][18] , \mult_19/CARRYB[15][19] ,
         \mult_19/CARRYB[15][20] , \mult_19/CARRYB[15][21] ,
         \mult_19/CARRYB[15][22] , \mult_19/CARRYB[15][23] ,
         \mult_19/CARRYB[15][24] , \mult_19/CARRYB[15][25] ,
         \mult_19/CARRYB[15][26] , \mult_19/CARRYB[15][27] ,
         \mult_19/CARRYB[15][28] , \mult_19/CARRYB[15][29] ,
         \mult_19/CARRYB[15][30] , \mult_19/ab[1][31] , \mult_19/ab[2][0] ,
         \mult_19/ab[2][1] , \mult_19/ab[2][2] , \mult_19/ab[2][3] ,
         \mult_19/ab[2][4] , \mult_19/ab[2][5] , \mult_19/ab[2][6] ,
         \mult_19/ab[2][7] , \mult_19/ab[2][8] , \mult_19/ab[2][9] ,
         \mult_19/ab[2][10] , \mult_19/ab[2][11] , \mult_19/ab[2][12] ,
         \mult_19/ab[2][13] , \mult_19/ab[2][14] , \mult_19/ab[2][15] ,
         \mult_19/ab[2][16] , \mult_19/ab[2][17] , \mult_19/ab[2][18] ,
         \mult_19/ab[2][19] , \mult_19/ab[2][20] , \mult_19/ab[2][21] ,
         \mult_19/ab[2][22] , \mult_19/ab[2][23] , \mult_19/ab[2][24] ,
         \mult_19/ab[2][25] , \mult_19/ab[2][26] , \mult_19/ab[2][27] ,
         \mult_19/ab[2][28] , \mult_19/ab[2][29] , \mult_19/ab[2][30] ,
         \mult_19/ab[2][31] , \mult_19/ab[3][0] , \mult_19/ab[3][1] ,
         \mult_19/ab[3][2] , \mult_19/ab[3][3] , \mult_19/ab[3][4] ,
         \mult_19/ab[3][5] , \mult_19/ab[3][6] , \mult_19/ab[3][7] ,
         \mult_19/ab[3][8] , \mult_19/ab[3][9] , \mult_19/ab[3][10] ,
         \mult_19/ab[3][11] , \mult_19/ab[3][12] , \mult_19/ab[3][13] ,
         \mult_19/ab[3][14] , \mult_19/ab[3][15] , \mult_19/ab[3][16] ,
         \mult_19/ab[3][17] , \mult_19/ab[3][18] , \mult_19/ab[3][19] ,
         \mult_19/ab[3][20] , \mult_19/ab[3][21] , \mult_19/ab[3][22] ,
         \mult_19/ab[3][23] , \mult_19/ab[3][24] , \mult_19/ab[3][25] ,
         \mult_19/ab[3][26] , \mult_19/ab[3][27] , \mult_19/ab[3][28] ,
         \mult_19/ab[3][29] , \mult_19/ab[3][30] , \mult_19/ab[3][31] ,
         \mult_19/ab[4][0] , \mult_19/ab[4][1] , \mult_19/ab[4][2] ,
         \mult_19/ab[4][3] , \mult_19/ab[4][4] , \mult_19/ab[4][5] ,
         \mult_19/ab[4][6] , \mult_19/ab[4][7] , \mult_19/ab[4][8] ,
         \mult_19/ab[4][9] , \mult_19/ab[4][10] , \mult_19/ab[4][11] ,
         \mult_19/ab[4][12] , \mult_19/ab[4][13] , \mult_19/ab[4][14] ,
         \mult_19/ab[4][15] , \mult_19/ab[4][16] , \mult_19/ab[4][17] ,
         \mult_19/ab[4][18] , \mult_19/ab[4][19] , \mult_19/ab[4][20] ,
         \mult_19/ab[4][21] , \mult_19/ab[4][22] , \mult_19/ab[4][23] ,
         \mult_19/ab[4][24] , \mult_19/ab[4][25] , \mult_19/ab[4][26] ,
         \mult_19/ab[4][27] , \mult_19/ab[4][28] , \mult_19/ab[4][29] ,
         \mult_19/ab[4][30] , \mult_19/ab[4][31] , \mult_19/ab[5][0] ,
         \mult_19/ab[5][1] , \mult_19/ab[5][2] , \mult_19/ab[5][3] ,
         \mult_19/ab[5][4] , \mult_19/ab[5][5] , \mult_19/ab[5][6] ,
         \mult_19/ab[5][7] , \mult_19/ab[5][8] , \mult_19/ab[5][9] ,
         \mult_19/ab[5][10] , \mult_19/ab[5][11] , \mult_19/ab[5][12] ,
         \mult_19/ab[5][13] , \mult_19/ab[5][14] , \mult_19/ab[5][15] ,
         \mult_19/ab[5][16] , \mult_19/ab[5][17] , \mult_19/ab[5][18] ,
         \mult_19/ab[5][19] , \mult_19/ab[5][20] , \mult_19/ab[5][21] ,
         \mult_19/ab[5][22] , \mult_19/ab[5][23] , \mult_19/ab[5][24] ,
         \mult_19/ab[5][25] , \mult_19/ab[5][26] , \mult_19/ab[5][27] ,
         \mult_19/ab[5][28] , \mult_19/ab[5][29] , \mult_19/ab[5][30] ,
         \mult_19/ab[5][31] , \mult_19/ab[6][0] , \mult_19/ab[6][1] ,
         \mult_19/ab[6][2] , \mult_19/ab[6][3] , \mult_19/ab[6][4] ,
         \mult_19/ab[6][5] , \mult_19/ab[6][6] , \mult_19/ab[6][7] ,
         \mult_19/ab[6][8] , \mult_19/ab[6][9] , \mult_19/ab[6][10] ,
         \mult_19/ab[6][11] , \mult_19/ab[6][12] , \mult_19/ab[6][13] ,
         \mult_19/ab[6][14] , \mult_19/ab[6][15] , \mult_19/ab[6][16] ,
         \mult_19/ab[6][17] , \mult_19/ab[6][18] , \mult_19/ab[6][19] ,
         \mult_19/ab[6][20] , \mult_19/ab[6][21] , \mult_19/ab[6][22] ,
         \mult_19/ab[6][23] , \mult_19/ab[6][24] , \mult_19/ab[6][25] ,
         \mult_19/ab[6][26] , \mult_19/ab[6][27] , \mult_19/ab[6][28] ,
         \mult_19/ab[6][29] , \mult_19/ab[6][30] , \mult_19/ab[6][31] ,
         \mult_19/ab[7][0] , \mult_19/ab[7][1] , \mult_19/ab[7][2] ,
         \mult_19/ab[7][3] , \mult_19/ab[7][4] , \mult_19/ab[7][5] ,
         \mult_19/ab[7][6] , \mult_19/ab[7][7] , \mult_19/ab[7][8] ,
         \mult_19/ab[7][9] , \mult_19/ab[7][10] , \mult_19/ab[7][11] ,
         \mult_19/ab[7][12] , \mult_19/ab[7][13] , \mult_19/ab[7][14] ,
         \mult_19/ab[7][15] , \mult_19/ab[7][16] , \mult_19/ab[7][17] ,
         \mult_19/ab[7][18] , \mult_19/ab[7][19] , \mult_19/ab[7][20] ,
         \mult_19/ab[7][21] , \mult_19/ab[7][22] , \mult_19/ab[7][23] ,
         \mult_19/ab[7][24] , \mult_19/ab[7][25] , \mult_19/ab[7][26] ,
         \mult_19/ab[7][27] , \mult_19/ab[7][28] , \mult_19/ab[7][29] ,
         \mult_19/ab[7][30] , \mult_19/ab[7][31] , \mult_19/ab[8][0] ,
         \mult_19/ab[8][1] , \mult_19/ab[8][2] , \mult_19/ab[8][3] ,
         \mult_19/ab[8][4] , \mult_19/ab[8][5] , \mult_19/ab[8][6] ,
         \mult_19/ab[8][7] , \mult_19/ab[8][8] , \mult_19/ab[8][9] ,
         \mult_19/ab[8][10] , \mult_19/ab[8][11] , \mult_19/ab[8][12] ,
         \mult_19/ab[8][13] , \mult_19/ab[8][14] , \mult_19/ab[8][15] ,
         \mult_19/ab[8][16] , \mult_19/ab[8][17] , \mult_19/ab[8][18] ,
         \mult_19/ab[8][19] , \mult_19/ab[8][20] , \mult_19/ab[8][21] ,
         \mult_19/ab[8][22] , \mult_19/ab[8][23] , \mult_19/ab[8][24] ,
         \mult_19/ab[8][25] , \mult_19/ab[8][26] , \mult_19/ab[8][27] ,
         \mult_19/ab[8][28] , \mult_19/ab[8][29] , \mult_19/ab[8][30] ,
         \mult_19/ab[8][31] , \mult_19/ab[9][0] , \mult_19/ab[9][1] ,
         \mult_19/ab[9][2] , \mult_19/ab[9][3] , \mult_19/ab[9][4] ,
         \mult_19/ab[9][5] , \mult_19/ab[9][6] , \mult_19/ab[9][7] ,
         \mult_19/ab[9][8] , \mult_19/ab[9][9] , \mult_19/ab[9][10] ,
         \mult_19/ab[9][11] , \mult_19/ab[9][12] , \mult_19/ab[9][13] ,
         \mult_19/ab[9][14] , \mult_19/ab[9][15] , \mult_19/ab[9][16] ,
         \mult_19/ab[9][17] , \mult_19/ab[9][18] , \mult_19/ab[9][19] ,
         \mult_19/ab[9][20] , \mult_19/ab[9][21] , \mult_19/ab[9][22] ,
         \mult_19/ab[9][23] , \mult_19/ab[9][24] , \mult_19/ab[9][25] ,
         \mult_19/ab[9][26] , \mult_19/ab[9][27] , \mult_19/ab[9][28] ,
         \mult_19/ab[9][29] , \mult_19/ab[9][30] , \mult_19/ab[9][31] ,
         \mult_19/ab[10][0] , \mult_19/ab[10][1] , \mult_19/ab[10][2] ,
         \mult_19/ab[10][3] , \mult_19/ab[10][4] , \mult_19/ab[10][5] ,
         \mult_19/ab[10][6] , \mult_19/ab[10][7] , \mult_19/ab[10][8] ,
         \mult_19/ab[10][9] , \mult_19/ab[10][10] , \mult_19/ab[10][11] ,
         \mult_19/ab[10][12] , \mult_19/ab[10][13] , \mult_19/ab[10][14] ,
         \mult_19/ab[10][15] , \mult_19/ab[10][16] , \mult_19/ab[10][17] ,
         \mult_19/ab[10][18] , \mult_19/ab[10][19] , \mult_19/ab[10][20] ,
         \mult_19/ab[10][21] , \mult_19/ab[10][22] , \mult_19/ab[10][23] ,
         \mult_19/ab[10][24] , \mult_19/ab[10][25] , \mult_19/ab[10][26] ,
         \mult_19/ab[10][27] , \mult_19/ab[10][28] , \mult_19/ab[10][29] ,
         \mult_19/ab[10][30] , \mult_19/ab[10][31] , \mult_19/ab[11][0] ,
         \mult_19/ab[11][1] , \mult_19/ab[11][2] , \mult_19/ab[11][3] ,
         \mult_19/ab[11][4] , \mult_19/ab[11][5] , \mult_19/ab[11][6] ,
         \mult_19/ab[11][7] , \mult_19/ab[11][8] , \mult_19/ab[11][9] ,
         \mult_19/ab[11][10] , \mult_19/ab[11][11] , \mult_19/ab[11][12] ,
         \mult_19/ab[11][13] , \mult_19/ab[11][14] , \mult_19/ab[11][15] ,
         \mult_19/ab[11][16] , \mult_19/ab[11][17] , \mult_19/ab[11][18] ,
         \mult_19/ab[11][19] , \mult_19/ab[11][20] , \mult_19/ab[11][21] ,
         \mult_19/ab[11][22] , \mult_19/ab[11][23] , \mult_19/ab[11][24] ,
         \mult_19/ab[11][25] , \mult_19/ab[11][26] , \mult_19/ab[11][27] ,
         \mult_19/ab[11][28] , \mult_19/ab[11][29] , \mult_19/ab[11][30] ,
         \mult_19/ab[11][31] , \mult_19/ab[12][0] , \mult_19/ab[12][1] ,
         \mult_19/ab[12][2] , \mult_19/ab[12][3] , \mult_19/ab[12][4] ,
         \mult_19/ab[12][5] , \mult_19/ab[12][6] , \mult_19/ab[12][7] ,
         \mult_19/ab[12][8] , \mult_19/ab[12][9] , \mult_19/ab[12][10] ,
         \mult_19/ab[12][11] , \mult_19/ab[12][12] , \mult_19/ab[12][13] ,
         \mult_19/ab[12][14] , \mult_19/ab[12][15] , \mult_19/ab[12][16] ,
         \mult_19/ab[12][17] , \mult_19/ab[12][18] , \mult_19/ab[12][19] ,
         \mult_19/ab[12][20] , \mult_19/ab[12][21] , \mult_19/ab[12][22] ,
         \mult_19/ab[12][23] , \mult_19/ab[12][24] , \mult_19/ab[12][25] ,
         \mult_19/ab[12][26] , \mult_19/ab[12][27] , \mult_19/ab[12][28] ,
         \mult_19/ab[12][29] , \mult_19/ab[12][30] , \mult_19/ab[12][31] ,
         \mult_19/ab[13][0] , \mult_19/ab[13][1] , \mult_19/ab[13][2] ,
         \mult_19/ab[13][3] , \mult_19/ab[13][4] , \mult_19/ab[13][5] ,
         \mult_19/ab[13][6] , \mult_19/ab[13][7] , \mult_19/ab[13][8] ,
         \mult_19/ab[13][9] , \mult_19/ab[13][10] , \mult_19/ab[13][11] ,
         \mult_19/ab[13][12] , \mult_19/ab[13][13] , \mult_19/ab[13][14] ,
         \mult_19/ab[13][15] , \mult_19/ab[13][16] , \mult_19/ab[13][17] ,
         \mult_19/ab[13][18] , \mult_19/ab[13][19] , \mult_19/ab[13][20] ,
         \mult_19/ab[13][21] , \mult_19/ab[13][22] , \mult_19/ab[13][23] ,
         \mult_19/ab[13][24] , \mult_19/ab[13][25] , \mult_19/ab[13][26] ,
         \mult_19/ab[13][27] , \mult_19/ab[13][28] , \mult_19/ab[13][29] ,
         \mult_19/ab[13][30] , \mult_19/ab[13][31] , \mult_19/ab[14][0] ,
         \mult_19/ab[14][1] , \mult_19/ab[14][2] , \mult_19/ab[14][3] ,
         \mult_19/ab[14][4] , \mult_19/ab[14][5] , \mult_19/ab[14][6] ,
         \mult_19/ab[14][7] , \mult_19/ab[14][8] , \mult_19/ab[14][9] ,
         \mult_19/ab[14][10] , \mult_19/ab[14][11] , \mult_19/ab[14][12] ,
         \mult_19/ab[14][13] , \mult_19/ab[14][14] , \mult_19/ab[14][15] ,
         \mult_19/ab[14][16] , \mult_19/ab[14][17] , \mult_19/ab[14][18] ,
         \mult_19/ab[14][19] , \mult_19/ab[14][20] , \mult_19/ab[14][21] ,
         \mult_19/ab[14][22] , \mult_19/ab[14][23] , \mult_19/ab[14][24] ,
         \mult_19/ab[14][25] , \mult_19/ab[14][26] , \mult_19/ab[14][27] ,
         \mult_19/ab[14][28] , \mult_19/ab[14][29] , \mult_19/ab[14][30] ,
         \mult_19/ab[14][31] , \mult_19/ab[15][0] , \mult_19/ab[15][1] ,
         \mult_19/ab[15][2] , \mult_19/ab[15][3] , \mult_19/ab[15][4] ,
         \mult_19/ab[15][5] , \mult_19/ab[15][6] , \mult_19/ab[15][7] ,
         \mult_19/ab[15][8] , \mult_19/ab[15][9] , \mult_19/ab[15][10] ,
         \mult_19/ab[15][11] , \mult_19/ab[15][12] , \mult_19/ab[15][13] ,
         \mult_19/ab[15][14] , \mult_19/ab[15][15] , \mult_19/ab[15][16] ,
         \mult_19/ab[15][17] , \mult_19/ab[15][18] , \mult_19/ab[15][19] ,
         \mult_19/ab[15][20] , \mult_19/ab[15][21] , \mult_19/ab[15][22] ,
         \mult_19/ab[15][23] , \mult_19/ab[15][24] , \mult_19/ab[15][25] ,
         \mult_19/ab[15][26] , \mult_19/ab[15][27] , \mult_19/ab[15][28] ,
         \mult_19/ab[15][29] , \mult_19/ab[15][30] , \mult_19/ab[15][31] ,
         \mult_19/ab[16][0] , \mult_19/ab[16][1] , \mult_19/ab[16][2] ,
         \mult_19/ab[16][3] , \mult_19/ab[16][4] , \mult_19/ab[16][5] ,
         \mult_19/ab[16][6] , \mult_19/ab[16][7] , \mult_19/ab[16][8] ,
         \mult_19/ab[16][9] , \mult_19/ab[16][10] , \mult_19/ab[16][11] ,
         \mult_19/ab[16][12] , \mult_19/ab[16][13] , \mult_19/ab[16][14] ,
         \mult_19/ab[16][15] , \mult_19/ab[16][16] , \mult_19/ab[16][17] ,
         \mult_19/ab[16][18] , \mult_19/ab[16][19] , \mult_19/ab[16][20] ,
         \mult_19/ab[16][21] , \mult_19/ab[16][22] , \mult_19/ab[16][23] ,
         \mult_19/ab[16][24] , \mult_19/ab[16][25] , \mult_19/ab[16][26] ,
         \mult_19/ab[16][27] , \mult_19/ab[16][28] , \mult_19/ab[16][29] ,
         \mult_19/ab[16][30] , \mult_19/ab[16][31] , \mult_19/ab[17][0] ,
         \mult_19/ab[17][1] , \mult_19/ab[17][2] , \mult_19/ab[17][3] ,
         \mult_19/ab[17][4] , \mult_19/ab[17][5] , \mult_19/ab[17][6] ,
         \mult_19/ab[17][7] , \mult_19/ab[17][8] , \mult_19/ab[17][9] ,
         \mult_19/ab[17][10] , \mult_19/ab[17][11] , \mult_19/ab[17][12] ,
         \mult_19/ab[17][13] , \mult_19/ab[17][14] , \mult_19/ab[17][15] ,
         \mult_19/ab[17][16] , \mult_19/ab[17][17] , \mult_19/ab[17][18] ,
         \mult_19/ab[17][19] , \mult_19/ab[17][20] , \mult_19/ab[17][21] ,
         \mult_19/ab[17][22] , \mult_19/ab[17][23] , \mult_19/ab[17][24] ,
         \mult_19/ab[17][25] , \mult_19/ab[17][26] , \mult_19/ab[17][27] ,
         \mult_19/ab[17][28] , \mult_19/ab[17][29] , \mult_19/ab[17][30] ,
         \mult_19/ab[17][31] , \mult_19/ab[18][0] , \mult_19/ab[18][1] ,
         \mult_19/ab[18][2] , \mult_19/ab[18][3] , \mult_19/ab[18][4] ,
         \mult_19/ab[18][5] , \mult_19/ab[18][6] , \mult_19/ab[18][7] ,
         \mult_19/ab[18][8] , \mult_19/ab[18][9] , \mult_19/ab[18][10] ,
         \mult_19/ab[18][11] , \mult_19/ab[18][12] , \mult_19/ab[18][13] ,
         \mult_19/ab[18][14] , \mult_19/ab[18][15] , \mult_19/ab[18][16] ,
         \mult_19/ab[18][17] , \mult_19/ab[18][18] , \mult_19/ab[18][19] ,
         \mult_19/ab[18][20] , \mult_19/ab[18][21] , \mult_19/ab[18][22] ,
         \mult_19/ab[18][23] , \mult_19/ab[18][24] , \mult_19/ab[18][25] ,
         \mult_19/ab[18][26] , \mult_19/ab[18][27] , \mult_19/ab[18][28] ,
         \mult_19/ab[18][29] , \mult_19/ab[18][30] , \mult_19/ab[18][31] ,
         \mult_19/ab[19][0] , \mult_19/ab[19][1] , \mult_19/ab[19][2] ,
         \mult_19/ab[19][3] , \mult_19/ab[19][4] , \mult_19/ab[19][5] ,
         \mult_19/ab[19][6] , \mult_19/ab[19][7] , \mult_19/ab[19][8] ,
         \mult_19/ab[19][9] , \mult_19/ab[19][10] , \mult_19/ab[19][11] ,
         \mult_19/ab[19][12] , \mult_19/ab[19][13] , \mult_19/ab[19][14] ,
         \mult_19/ab[19][15] , \mult_19/ab[19][16] , \mult_19/ab[19][17] ,
         \mult_19/ab[19][18] , \mult_19/ab[19][19] , \mult_19/ab[19][20] ,
         \mult_19/ab[19][21] , \mult_19/ab[19][22] , \mult_19/ab[19][23] ,
         \mult_19/ab[19][24] , \mult_19/ab[19][25] , \mult_19/ab[19][26] ,
         \mult_19/ab[19][27] , \mult_19/ab[19][28] , \mult_19/ab[19][29] ,
         \mult_19/ab[19][30] , \mult_19/ab[19][31] , \mult_19/ab[20][0] ,
         \mult_19/ab[20][1] , \mult_19/ab[20][2] , \mult_19/ab[20][3] ,
         \mult_19/ab[20][4] , \mult_19/ab[20][5] , \mult_19/ab[20][6] ,
         \mult_19/ab[20][7] , \mult_19/ab[20][8] , \mult_19/ab[20][9] ,
         \mult_19/ab[20][10] , \mult_19/ab[20][11] , \mult_19/ab[20][12] ,
         \mult_19/ab[20][13] , \mult_19/ab[20][14] , \mult_19/ab[20][15] ,
         \mult_19/ab[20][16] , \mult_19/ab[20][17] , \mult_19/ab[20][18] ,
         \mult_19/ab[20][19] , \mult_19/ab[20][20] , \mult_19/ab[20][21] ,
         \mult_19/ab[20][22] , \mult_19/ab[20][23] , \mult_19/ab[20][24] ,
         \mult_19/ab[20][25] , \mult_19/ab[20][26] , \mult_19/ab[20][27] ,
         \mult_19/ab[20][28] , \mult_19/ab[20][29] , \mult_19/ab[20][30] ,
         \mult_19/ab[20][31] , \mult_19/ab[21][0] , \mult_19/ab[21][1] ,
         \mult_19/ab[21][2] , \mult_19/ab[21][3] , \mult_19/ab[21][4] ,
         \mult_19/ab[21][5] , \mult_19/ab[21][6] , \mult_19/ab[21][7] ,
         \mult_19/ab[21][8] , \mult_19/ab[21][9] , \mult_19/ab[21][10] ,
         \mult_19/ab[21][11] , \mult_19/ab[21][12] , \mult_19/ab[21][13] ,
         \mult_19/ab[21][14] , \mult_19/ab[21][15] , \mult_19/ab[21][16] ,
         \mult_19/ab[21][17] , \mult_19/ab[21][18] , \mult_19/ab[21][19] ,
         \mult_19/ab[21][20] , \mult_19/ab[21][21] , \mult_19/ab[21][22] ,
         \mult_19/ab[21][23] , \mult_19/ab[21][24] , \mult_19/ab[21][25] ,
         \mult_19/ab[21][26] , \mult_19/ab[21][27] , \mult_19/ab[21][28] ,
         \mult_19/ab[21][29] , \mult_19/ab[21][30] , \mult_19/ab[21][31] ,
         \mult_19/ab[22][0] , \mult_19/ab[22][1] , \mult_19/ab[22][2] ,
         \mult_19/ab[22][3] , \mult_19/ab[22][4] , \mult_19/ab[22][5] ,
         \mult_19/ab[22][6] , \mult_19/ab[22][7] , \mult_19/ab[22][8] ,
         \mult_19/ab[22][9] , \mult_19/ab[22][10] , \mult_19/ab[22][11] ,
         \mult_19/ab[22][12] , \mult_19/ab[22][13] , \mult_19/ab[22][14] ,
         \mult_19/ab[22][15] , \mult_19/ab[22][16] , \mult_19/ab[22][17] ,
         \mult_19/ab[22][18] , \mult_19/ab[22][19] , \mult_19/ab[22][20] ,
         \mult_19/ab[22][21] , \mult_19/ab[22][22] , \mult_19/ab[22][23] ,
         \mult_19/ab[22][24] , \mult_19/ab[22][25] , \mult_19/ab[22][26] ,
         \mult_19/ab[22][27] , \mult_19/ab[22][28] , \mult_19/ab[22][29] ,
         \mult_19/ab[22][30] , \mult_19/ab[22][31] , \mult_19/ab[23][0] ,
         \mult_19/ab[23][1] , \mult_19/ab[23][2] , \mult_19/ab[23][3] ,
         \mult_19/ab[23][4] , \mult_19/ab[23][5] , \mult_19/ab[23][6] ,
         \mult_19/ab[23][7] , \mult_19/ab[23][8] , \mult_19/ab[23][9] ,
         \mult_19/ab[23][10] , \mult_19/ab[23][11] , \mult_19/ab[23][12] ,
         \mult_19/ab[23][13] , \mult_19/ab[23][14] , \mult_19/ab[23][15] ,
         \mult_19/ab[23][16] , \mult_19/ab[23][17] , \mult_19/ab[23][18] ,
         \mult_19/ab[23][19] , \mult_19/ab[23][20] , \mult_19/ab[23][21] ,
         \mult_19/ab[23][22] , \mult_19/ab[23][23] , \mult_19/ab[23][24] ,
         \mult_19/ab[23][25] , \mult_19/ab[23][26] , \mult_19/ab[23][27] ,
         \mult_19/ab[23][28] , \mult_19/ab[23][29] , \mult_19/ab[23][30] ,
         \mult_19/ab[23][31] , \mult_19/ab[24][0] , \mult_19/ab[24][1] ,
         \mult_19/ab[24][2] , \mult_19/ab[24][3] , \mult_19/ab[24][4] ,
         \mult_19/ab[24][5] , \mult_19/ab[24][6] , \mult_19/ab[24][7] ,
         \mult_19/ab[24][8] , \mult_19/ab[24][9] , \mult_19/ab[24][10] ,
         \mult_19/ab[24][11] , \mult_19/ab[24][12] , \mult_19/ab[24][13] ,
         \mult_19/ab[24][14] , \mult_19/ab[24][15] , \mult_19/ab[24][16] ,
         \mult_19/ab[24][17] , \mult_19/ab[24][18] , \mult_19/ab[24][19] ,
         \mult_19/ab[24][20] , \mult_19/ab[24][21] , \mult_19/ab[24][22] ,
         \mult_19/ab[24][23] , \mult_19/ab[24][24] , \mult_19/ab[24][25] ,
         \mult_19/ab[24][26] , \mult_19/ab[24][27] , \mult_19/ab[24][28] ,
         \mult_19/ab[24][29] , \mult_19/ab[24][30] , \mult_19/ab[24][31] ,
         \mult_19/ab[25][0] , \mult_19/ab[25][1] , \mult_19/ab[25][2] ,
         \mult_19/ab[25][3] , \mult_19/ab[25][4] , \mult_19/ab[25][5] ,
         \mult_19/ab[25][6] , \mult_19/ab[25][7] , \mult_19/ab[25][8] ,
         \mult_19/ab[25][9] , \mult_19/ab[25][10] , \mult_19/ab[25][11] ,
         \mult_19/ab[25][12] , \mult_19/ab[25][13] , \mult_19/ab[25][14] ,
         \mult_19/ab[25][15] , \mult_19/ab[25][16] , \mult_19/ab[25][17] ,
         \mult_19/ab[25][18] , \mult_19/ab[25][19] , \mult_19/ab[25][20] ,
         \mult_19/ab[25][21] , \mult_19/ab[25][22] , \mult_19/ab[25][23] ,
         \mult_19/ab[25][24] , \mult_19/ab[25][25] , \mult_19/ab[25][26] ,
         \mult_19/ab[25][27] , \mult_19/ab[25][28] , \mult_19/ab[25][29] ,
         \mult_19/ab[25][30] , \mult_19/ab[25][31] , \mult_19/ab[26][0] ,
         \mult_19/ab[26][1] , \mult_19/ab[26][2] , \mult_19/ab[26][3] ,
         \mult_19/ab[26][4] , \mult_19/ab[26][5] , \mult_19/ab[26][6] ,
         \mult_19/ab[26][7] , \mult_19/ab[26][8] , \mult_19/ab[26][9] ,
         \mult_19/ab[26][10] , \mult_19/ab[26][11] , \mult_19/ab[26][12] ,
         \mult_19/ab[26][13] , \mult_19/ab[26][14] , \mult_19/ab[26][15] ,
         \mult_19/ab[26][16] , \mult_19/ab[26][17] , \mult_19/ab[26][18] ,
         \mult_19/ab[26][19] , \mult_19/ab[26][20] , \mult_19/ab[26][21] ,
         \mult_19/ab[26][22] , \mult_19/ab[26][23] , \mult_19/ab[26][24] ,
         \mult_19/ab[26][25] , \mult_19/ab[26][26] , \mult_19/ab[26][27] ,
         \mult_19/ab[26][28] , \mult_19/ab[26][29] , \mult_19/ab[26][30] ,
         \mult_19/ab[26][31] , \mult_19/ab[27][0] , \mult_19/ab[27][1] ,
         \mult_19/ab[27][2] , \mult_19/ab[27][3] , \mult_19/ab[27][4] ,
         \mult_19/ab[27][5] , \mult_19/ab[27][6] , \mult_19/ab[27][7] ,
         \mult_19/ab[27][8] , \mult_19/ab[27][9] , \mult_19/ab[27][10] ,
         \mult_19/ab[27][11] , \mult_19/ab[27][12] , \mult_19/ab[27][13] ,
         \mult_19/ab[27][14] , \mult_19/ab[27][15] , \mult_19/ab[27][16] ,
         \mult_19/ab[27][17] , \mult_19/ab[27][18] , \mult_19/ab[27][19] ,
         \mult_19/ab[27][20] , \mult_19/ab[27][21] , \mult_19/ab[27][22] ,
         \mult_19/ab[27][23] , \mult_19/ab[27][24] , \mult_19/ab[27][25] ,
         \mult_19/ab[27][26] , \mult_19/ab[27][27] , \mult_19/ab[27][28] ,
         \mult_19/ab[27][29] , \mult_19/ab[27][30] , \mult_19/ab[27][31] ,
         \mult_19/ab[28][0] , \mult_19/ab[28][1] , \mult_19/ab[28][2] ,
         \mult_19/ab[28][3] , \mult_19/ab[28][4] , \mult_19/ab[28][5] ,
         \mult_19/ab[28][6] , \mult_19/ab[28][7] , \mult_19/ab[28][8] ,
         \mult_19/ab[28][9] , \mult_19/ab[28][10] , \mult_19/ab[28][11] ,
         \mult_19/ab[28][12] , \mult_19/ab[28][13] , \mult_19/ab[28][14] ,
         \mult_19/ab[28][15] , \mult_19/ab[28][16] , \mult_19/ab[28][17] ,
         \mult_19/ab[28][18] , \mult_19/ab[28][19] , \mult_19/ab[28][20] ,
         \mult_19/ab[28][21] , \mult_19/ab[28][22] , \mult_19/ab[28][23] ,
         \mult_19/ab[28][24] , \mult_19/ab[28][25] , \mult_19/ab[28][26] ,
         \mult_19/ab[28][27] , \mult_19/ab[28][28] , \mult_19/ab[28][29] ,
         \mult_19/ab[28][30] , \mult_19/ab[28][31] , \mult_19/ab[29][0] ,
         \mult_19/ab[29][1] , \mult_19/ab[29][2] , \mult_19/ab[29][3] ,
         \mult_19/ab[29][4] , \mult_19/ab[29][5] , \mult_19/ab[29][6] ,
         \mult_19/ab[29][7] , \mult_19/ab[29][8] , \mult_19/ab[29][9] ,
         \mult_19/ab[29][10] , \mult_19/ab[29][11] , \mult_19/ab[29][12] ,
         \mult_19/ab[29][13] , \mult_19/ab[29][14] , \mult_19/ab[29][15] ,
         \mult_19/ab[29][16] , \mult_19/ab[29][17] , \mult_19/ab[29][18] ,
         \mult_19/ab[29][19] , \mult_19/ab[29][20] , \mult_19/ab[29][21] ,
         \mult_19/ab[29][22] , \mult_19/ab[29][23] , \mult_19/ab[29][24] ,
         \mult_19/ab[29][25] , \mult_19/ab[29][26] , \mult_19/ab[29][27] ,
         \mult_19/ab[29][28] , \mult_19/ab[29][29] , \mult_19/ab[29][30] ,
         \mult_19/ab[29][31] , \mult_19/ab[30][0] , \mult_19/ab[30][1] ,
         \mult_19/ab[30][2] , \mult_19/ab[30][3] , \mult_19/ab[30][4] ,
         \mult_19/ab[30][5] , \mult_19/ab[30][6] , \mult_19/ab[30][7] ,
         \mult_19/ab[30][8] , \mult_19/ab[30][9] , \mult_19/ab[30][10] ,
         \mult_19/ab[30][11] , \mult_19/ab[30][12] , \mult_19/ab[30][13] ,
         \mult_19/ab[30][14] , \mult_19/ab[30][15] , \mult_19/ab[30][16] ,
         \mult_19/ab[30][17] , \mult_19/ab[30][18] , \mult_19/ab[30][19] ,
         \mult_19/ab[30][20] , \mult_19/ab[30][21] , \mult_19/ab[30][22] ,
         \mult_19/ab[30][23] , \mult_19/ab[30][24] , \mult_19/ab[30][25] ,
         \mult_19/ab[30][26] , \mult_19/ab[30][27] , \mult_19/ab[30][28] ,
         \mult_19/ab[30][29] , \mult_19/ab[30][30] , \mult_19/ab[30][31] ,
         \mult_19/ab[31][0] , \mult_19/ab[31][1] , \mult_19/ab[31][2] ,
         \mult_19/ab[31][3] , \mult_19/ab[31][4] , \mult_19/ab[31][5] ,
         \mult_19/ab[31][6] , \mult_19/ab[31][7] , \mult_19/ab[31][8] ,
         \mult_19/ab[31][9] , \mult_19/ab[31][10] , \mult_19/ab[31][11] ,
         \mult_19/ab[31][12] , \mult_19/ab[31][13] , \mult_19/ab[31][14] ,
         \mult_19/ab[31][15] , \mult_19/ab[31][16] , \mult_19/ab[31][17] ,
         \mult_19/ab[31][18] , \mult_19/ab[31][19] , \mult_19/ab[31][20] ,
         \mult_19/ab[31][21] , \mult_19/ab[31][22] , \mult_19/ab[31][23] ,
         \mult_19/ab[31][24] , \mult_19/ab[31][25] , \mult_19/ab[31][26] ,
         \mult_19/ab[31][27] , \mult_19/ab[31][28] , \mult_19/ab[31][29] ,
         \mult_19/ab[31][30] , \mult_22/n325 , \mult_22/n324 , \mult_22/n323 ,
         \mult_22/n322 , \mult_22/n196 , \mult_22/n195 , \mult_22/n194 ,
         \mult_22/n181 , \mult_22/n163 , \mult_22/n159 , \mult_22/n114 ,
         \mult_22/n113 , \mult_22/n112 , \mult_22/n111 , \mult_22/n110 ,
         \mult_22/n109 , \mult_22/n108 , \mult_22/n107 , \mult_22/n106 ,
         \mult_22/n105 , \mult_22/n104 , \mult_22/n103 , \mult_22/n102 ,
         \mult_22/n101 , \mult_22/n100 , \mult_22/n99 , \mult_22/n98 ,
         \mult_22/n97 , \mult_22/n96 , \mult_22/n95 , \mult_22/n94 ,
         \mult_22/n93 , \mult_22/n92 , \mult_22/n91 , \mult_22/n90 ,
         \mult_22/n89 , \mult_22/n88 , \mult_22/n87 , \mult_22/n86 ,
         \mult_22/n85 , \mult_22/n84 , \mult_22/n83 , \mult_22/n82 ,
         \mult_22/n81 , \mult_22/n80 , \mult_22/n79 , \mult_22/n78 ,
         \mult_22/n77 , \mult_22/n76 , \mult_22/n75 , \mult_22/n74 ,
         \mult_22/n73 , \mult_22/n72 , \mult_22/n71 , \mult_22/n70 ,
         \mult_22/n69 , \mult_22/n68 , \mult_22/n67 , \mult_22/n66 ,
         \mult_22/n65 , \mult_22/n64 , \mult_22/n63 , \mult_22/n62 ,
         \mult_22/n61 , \mult_22/n60 , \mult_22/n59 , \mult_22/n58 ,
         \mult_22/n57 , \mult_22/n56 , \mult_22/n55 , \mult_22/n54 ,
         \mult_22/n53 , \mult_22/n52 , \mult_22/n51 , \mult_22/n50 ,
         \mult_22/n49 , \mult_22/n48 , \mult_22/n47 , \mult_22/n46 ,
         \mult_22/n45 , \mult_22/n44 , \mult_22/n43 , \mult_22/n42 ,
         \mult_22/n41 , \mult_22/n40 , \mult_22/n39 , \mult_22/n38 ,
         \mult_22/n37 , \mult_22/n36 , \mult_22/n35 , \mult_22/n34 ,
         \mult_22/n33 , \mult_22/n32 , \mult_22/n31 , \mult_22/n30 ,
         \mult_22/n29 , \mult_22/n28 , \mult_22/n27 , \mult_22/n26 ,
         \mult_22/n25 , \mult_22/n24 , \mult_22/n23 , \mult_22/n22 ,
         \mult_22/n21 , \mult_22/n20 , \mult_22/n19 , \mult_22/n18 ,
         \mult_22/n17 , \mult_22/n16 , \mult_22/n15 , \mult_22/n14 ,
         \mult_22/n13 , \mult_22/n12 , \mult_22/n11 , \mult_22/n10 ,
         \mult_22/n9 , \mult_22/n8 , \mult_22/n7 , \mult_22/n6 , \mult_22/n5 ,
         \mult_22/SUMB[56][1] , \mult_22/SUMB[56][2] , \mult_22/SUMB[56][3] ,
         \mult_22/SUMB[56][4] , \mult_22/SUMB[56][5] , \mult_22/SUMB[56][6] ,
         \mult_22/SUMB[56][7] , \mult_22/SUMB[56][8] , \mult_22/SUMB[56][9] ,
         \mult_22/SUMB[56][10] , \mult_22/SUMB[56][11] ,
         \mult_22/SUMB[56][12] , \mult_22/SUMB[56][13] ,
         \mult_22/SUMB[56][14] , \mult_22/SUMB[56][15] ,
         \mult_22/SUMB[56][16] , \mult_22/SUMB[56][17] ,
         \mult_22/SUMB[56][18] , \mult_22/SUMB[56][19] ,
         \mult_22/SUMB[56][20] , \mult_22/SUMB[56][21] ,
         \mult_22/SUMB[56][22] , \mult_22/SUMB[56][23] ,
         \mult_22/SUMB[56][24] , \mult_22/SUMB[56][25] ,
         \mult_22/SUMB[56][26] , \mult_22/SUMB[56][27] ,
         \mult_22/SUMB[56][28] , \mult_22/SUMB[56][29] ,
         \mult_22/SUMB[56][30] , \mult_22/SUMB[56][31] ,
         \mult_22/SUMB[56][32] , \mult_22/SUMB[56][33] ,
         \mult_22/SUMB[56][34] , \mult_22/SUMB[56][35] ,
         \mult_22/SUMB[56][36] , \mult_22/SUMB[56][37] ,
         \mult_22/SUMB[56][38] , \mult_22/SUMB[56][39] ,
         \mult_22/SUMB[56][40] , \mult_22/SUMB[56][41] ,
         \mult_22/SUMB[56][42] , \mult_22/SUMB[56][43] ,
         \mult_22/SUMB[56][44] , \mult_22/SUMB[56][45] ,
         \mult_22/SUMB[56][46] , \mult_22/SUMB[56][47] ,
         \mult_22/SUMB[56][48] , \mult_22/SUMB[56][49] ,
         \mult_22/SUMB[56][50] , \mult_22/SUMB[56][51] ,
         \mult_22/SUMB[56][52] , \mult_22/SUMB[56][53] ,
         \mult_22/SUMB[56][54] , \mult_22/SUMB[56][55] ,
         \mult_22/SUMB[56][56] , \mult_22/SUMB[56][57] ,
         \mult_22/SUMB[56][58] , \mult_22/SUMB[56][59] ,
         \mult_22/SUMB[56][60] , \mult_22/SUMB[56][61] ,
         \mult_22/SUMB[56][62] , \mult_22/SUMB[57][1] , \mult_22/SUMB[57][2] ,
         \mult_22/SUMB[57][3] , \mult_22/SUMB[57][4] , \mult_22/SUMB[57][5] ,
         \mult_22/SUMB[57][6] , \mult_22/SUMB[57][7] , \mult_22/SUMB[57][8] ,
         \mult_22/SUMB[57][9] , \mult_22/SUMB[57][10] , \mult_22/SUMB[57][11] ,
         \mult_22/SUMB[57][12] , \mult_22/SUMB[57][13] ,
         \mult_22/SUMB[57][14] , \mult_22/SUMB[57][15] ,
         \mult_22/SUMB[57][16] , \mult_22/SUMB[57][17] ,
         \mult_22/SUMB[57][18] , \mult_22/SUMB[57][19] ,
         \mult_22/SUMB[57][20] , \mult_22/SUMB[57][21] ,
         \mult_22/SUMB[57][22] , \mult_22/SUMB[57][23] ,
         \mult_22/SUMB[57][24] , \mult_22/SUMB[57][25] ,
         \mult_22/SUMB[57][26] , \mult_22/SUMB[57][27] ,
         \mult_22/SUMB[57][28] , \mult_22/SUMB[57][29] ,
         \mult_22/SUMB[57][30] , \mult_22/SUMB[57][31] ,
         \mult_22/SUMB[57][32] , \mult_22/SUMB[57][33] ,
         \mult_22/SUMB[57][34] , \mult_22/SUMB[57][35] ,
         \mult_22/SUMB[57][36] , \mult_22/SUMB[57][37] ,
         \mult_22/SUMB[57][38] , \mult_22/SUMB[57][39] ,
         \mult_22/SUMB[57][40] , \mult_22/SUMB[57][41] ,
         \mult_22/SUMB[57][42] , \mult_22/SUMB[57][43] ,
         \mult_22/SUMB[57][44] , \mult_22/SUMB[57][45] ,
         \mult_22/SUMB[57][46] , \mult_22/SUMB[57][47] ,
         \mult_22/SUMB[57][48] , \mult_22/SUMB[57][49] ,
         \mult_22/SUMB[57][50] , \mult_22/SUMB[57][51] ,
         \mult_22/SUMB[57][52] , \mult_22/SUMB[57][53] ,
         \mult_22/SUMB[57][54] , \mult_22/SUMB[57][55] ,
         \mult_22/SUMB[57][56] , \mult_22/SUMB[57][57] ,
         \mult_22/SUMB[57][58] , \mult_22/SUMB[57][59] ,
         \mult_22/SUMB[57][60] , \mult_22/SUMB[57][61] ,
         \mult_22/SUMB[57][62] , \mult_22/SUMB[58][1] , \mult_22/SUMB[58][2] ,
         \mult_22/SUMB[58][3] , \mult_22/SUMB[58][4] , \mult_22/SUMB[58][5] ,
         \mult_22/SUMB[58][6] , \mult_22/SUMB[58][7] , \mult_22/SUMB[58][8] ,
         \mult_22/SUMB[58][9] , \mult_22/SUMB[58][10] , \mult_22/SUMB[58][11] ,
         \mult_22/SUMB[58][12] , \mult_22/SUMB[58][13] ,
         \mult_22/SUMB[58][14] , \mult_22/SUMB[58][15] ,
         \mult_22/SUMB[58][16] , \mult_22/SUMB[58][17] ,
         \mult_22/SUMB[58][18] , \mult_22/SUMB[58][19] ,
         \mult_22/SUMB[58][20] , \mult_22/SUMB[58][21] ,
         \mult_22/SUMB[58][22] , \mult_22/SUMB[58][23] ,
         \mult_22/SUMB[58][24] , \mult_22/SUMB[58][25] ,
         \mult_22/SUMB[58][26] , \mult_22/SUMB[58][27] ,
         \mult_22/SUMB[58][28] , \mult_22/SUMB[58][29] ,
         \mult_22/SUMB[58][30] , \mult_22/SUMB[58][31] ,
         \mult_22/SUMB[58][32] , \mult_22/SUMB[58][33] ,
         \mult_22/SUMB[58][34] , \mult_22/SUMB[58][35] ,
         \mult_22/SUMB[58][36] , \mult_22/SUMB[58][37] ,
         \mult_22/SUMB[58][38] , \mult_22/SUMB[58][39] ,
         \mult_22/SUMB[58][40] , \mult_22/SUMB[58][41] ,
         \mult_22/SUMB[58][42] , \mult_22/SUMB[58][43] ,
         \mult_22/SUMB[58][44] , \mult_22/SUMB[58][45] ,
         \mult_22/SUMB[58][46] , \mult_22/SUMB[58][47] ,
         \mult_22/SUMB[58][48] , \mult_22/SUMB[58][49] ,
         \mult_22/SUMB[58][50] , \mult_22/SUMB[58][51] ,
         \mult_22/SUMB[58][52] , \mult_22/SUMB[58][53] ,
         \mult_22/SUMB[58][54] , \mult_22/SUMB[58][55] ,
         \mult_22/SUMB[58][56] , \mult_22/SUMB[58][57] ,
         \mult_22/SUMB[58][58] , \mult_22/SUMB[58][59] ,
         \mult_22/SUMB[58][60] , \mult_22/SUMB[58][61] ,
         \mult_22/SUMB[58][62] , \mult_22/SUMB[59][1] , \mult_22/SUMB[59][2] ,
         \mult_22/SUMB[59][3] , \mult_22/SUMB[59][4] , \mult_22/SUMB[59][5] ,
         \mult_22/SUMB[59][6] , \mult_22/SUMB[59][7] , \mult_22/SUMB[59][8] ,
         \mult_22/SUMB[59][9] , \mult_22/SUMB[59][10] , \mult_22/SUMB[59][11] ,
         \mult_22/SUMB[59][12] , \mult_22/SUMB[59][13] ,
         \mult_22/SUMB[59][14] , \mult_22/SUMB[59][15] ,
         \mult_22/SUMB[59][16] , \mult_22/SUMB[59][17] ,
         \mult_22/SUMB[59][18] , \mult_22/SUMB[59][19] ,
         \mult_22/SUMB[59][20] , \mult_22/SUMB[59][21] ,
         \mult_22/SUMB[59][22] , \mult_22/SUMB[59][23] ,
         \mult_22/SUMB[59][24] , \mult_22/SUMB[59][25] ,
         \mult_22/SUMB[59][26] , \mult_22/SUMB[59][27] ,
         \mult_22/SUMB[59][28] , \mult_22/SUMB[59][29] ,
         \mult_22/SUMB[59][30] , \mult_22/SUMB[59][31] ,
         \mult_22/SUMB[59][32] , \mult_22/SUMB[59][33] ,
         \mult_22/SUMB[59][34] , \mult_22/SUMB[59][35] ,
         \mult_22/SUMB[59][36] , \mult_22/SUMB[59][37] ,
         \mult_22/SUMB[59][38] , \mult_22/SUMB[59][39] ,
         \mult_22/SUMB[59][40] , \mult_22/SUMB[59][41] ,
         \mult_22/SUMB[59][42] , \mult_22/SUMB[59][43] ,
         \mult_22/SUMB[59][44] , \mult_22/SUMB[59][45] ,
         \mult_22/SUMB[59][46] , \mult_22/SUMB[59][47] ,
         \mult_22/SUMB[59][48] , \mult_22/SUMB[59][49] ,
         \mult_22/SUMB[59][50] , \mult_22/SUMB[59][51] ,
         \mult_22/SUMB[59][52] , \mult_22/SUMB[59][53] ,
         \mult_22/SUMB[59][54] , \mult_22/SUMB[59][55] ,
         \mult_22/SUMB[59][56] , \mult_22/SUMB[59][57] ,
         \mult_22/SUMB[59][58] , \mult_22/SUMB[59][59] ,
         \mult_22/SUMB[59][60] , \mult_22/SUMB[59][61] ,
         \mult_22/SUMB[59][62] , \mult_22/SUMB[60][1] , \mult_22/SUMB[60][2] ,
         \mult_22/SUMB[60][3] , \mult_22/SUMB[60][4] , \mult_22/SUMB[60][5] ,
         \mult_22/SUMB[60][6] , \mult_22/SUMB[60][7] , \mult_22/SUMB[60][8] ,
         \mult_22/SUMB[60][9] , \mult_22/SUMB[60][10] , \mult_22/SUMB[60][11] ,
         \mult_22/SUMB[60][12] , \mult_22/SUMB[60][13] ,
         \mult_22/SUMB[60][14] , \mult_22/SUMB[60][15] ,
         \mult_22/SUMB[60][16] , \mult_22/SUMB[60][17] ,
         \mult_22/SUMB[60][18] , \mult_22/SUMB[60][19] ,
         \mult_22/SUMB[60][20] , \mult_22/SUMB[60][21] ,
         \mult_22/SUMB[60][22] , \mult_22/SUMB[60][23] ,
         \mult_22/SUMB[60][24] , \mult_22/SUMB[60][25] ,
         \mult_22/SUMB[60][26] , \mult_22/SUMB[60][27] ,
         \mult_22/SUMB[60][28] , \mult_22/SUMB[60][29] ,
         \mult_22/SUMB[60][30] , \mult_22/SUMB[60][31] ,
         \mult_22/SUMB[60][32] , \mult_22/SUMB[60][33] ,
         \mult_22/SUMB[60][34] , \mult_22/SUMB[60][35] ,
         \mult_22/SUMB[60][36] , \mult_22/SUMB[60][37] ,
         \mult_22/SUMB[60][38] , \mult_22/SUMB[60][39] ,
         \mult_22/SUMB[60][40] , \mult_22/SUMB[60][41] ,
         \mult_22/SUMB[60][42] , \mult_22/SUMB[60][43] ,
         \mult_22/SUMB[60][44] , \mult_22/SUMB[60][45] ,
         \mult_22/SUMB[60][46] , \mult_22/SUMB[60][47] ,
         \mult_22/SUMB[60][48] , \mult_22/SUMB[60][49] ,
         \mult_22/SUMB[60][50] , \mult_22/SUMB[60][51] ,
         \mult_22/SUMB[60][52] , \mult_22/SUMB[60][53] ,
         \mult_22/SUMB[60][54] , \mult_22/SUMB[60][55] ,
         \mult_22/SUMB[60][56] , \mult_22/SUMB[60][57] ,
         \mult_22/SUMB[60][58] , \mult_22/SUMB[60][59] ,
         \mult_22/SUMB[60][60] , \mult_22/SUMB[60][61] ,
         \mult_22/SUMB[60][62] , \mult_22/SUMB[61][1] , \mult_22/SUMB[61][2] ,
         \mult_22/SUMB[61][3] , \mult_22/SUMB[61][4] , \mult_22/SUMB[61][5] ,
         \mult_22/SUMB[61][6] , \mult_22/SUMB[61][7] , \mult_22/SUMB[61][8] ,
         \mult_22/SUMB[61][9] , \mult_22/SUMB[61][10] , \mult_22/SUMB[61][11] ,
         \mult_22/SUMB[61][12] , \mult_22/SUMB[61][13] ,
         \mult_22/SUMB[61][14] , \mult_22/SUMB[61][15] ,
         \mult_22/SUMB[61][16] , \mult_22/SUMB[61][17] ,
         \mult_22/SUMB[61][18] , \mult_22/SUMB[61][19] ,
         \mult_22/SUMB[61][20] , \mult_22/SUMB[61][21] ,
         \mult_22/SUMB[61][22] , \mult_22/SUMB[61][23] ,
         \mult_22/SUMB[61][24] , \mult_22/SUMB[61][25] ,
         \mult_22/SUMB[61][26] , \mult_22/SUMB[61][27] ,
         \mult_22/SUMB[61][28] , \mult_22/SUMB[61][29] ,
         \mult_22/SUMB[61][30] , \mult_22/SUMB[61][31] ,
         \mult_22/SUMB[61][32] , \mult_22/SUMB[61][33] ,
         \mult_22/SUMB[61][34] , \mult_22/SUMB[61][35] ,
         \mult_22/SUMB[61][36] , \mult_22/SUMB[61][37] ,
         \mult_22/SUMB[61][38] , \mult_22/SUMB[61][39] ,
         \mult_22/SUMB[61][40] , \mult_22/SUMB[61][41] ,
         \mult_22/SUMB[61][42] , \mult_22/SUMB[61][43] ,
         \mult_22/SUMB[61][44] , \mult_22/SUMB[61][45] ,
         \mult_22/SUMB[61][46] , \mult_22/SUMB[61][47] ,
         \mult_22/SUMB[61][48] , \mult_22/SUMB[61][49] ,
         \mult_22/SUMB[61][50] , \mult_22/SUMB[61][51] ,
         \mult_22/SUMB[61][52] , \mult_22/SUMB[61][53] ,
         \mult_22/SUMB[61][54] , \mult_22/SUMB[61][55] ,
         \mult_22/SUMB[61][56] , \mult_22/SUMB[61][57] ,
         \mult_22/SUMB[61][58] , \mult_22/SUMB[61][59] ,
         \mult_22/SUMB[61][60] , \mult_22/SUMB[61][61] ,
         \mult_22/SUMB[61][62] , \mult_22/SUMB[62][1] , \mult_22/SUMB[62][2] ,
         \mult_22/SUMB[62][3] , \mult_22/SUMB[62][4] , \mult_22/SUMB[62][5] ,
         \mult_22/SUMB[62][6] , \mult_22/SUMB[62][7] , \mult_22/SUMB[62][8] ,
         \mult_22/SUMB[62][9] , \mult_22/SUMB[62][10] , \mult_22/SUMB[62][11] ,
         \mult_22/SUMB[62][12] , \mult_22/SUMB[62][13] ,
         \mult_22/SUMB[62][14] , \mult_22/SUMB[62][15] ,
         \mult_22/SUMB[62][16] , \mult_22/SUMB[62][17] ,
         \mult_22/SUMB[62][18] , \mult_22/SUMB[62][19] ,
         \mult_22/SUMB[62][20] , \mult_22/SUMB[62][21] ,
         \mult_22/SUMB[62][22] , \mult_22/SUMB[62][23] ,
         \mult_22/SUMB[62][24] , \mult_22/SUMB[62][25] ,
         \mult_22/SUMB[62][26] , \mult_22/SUMB[62][27] ,
         \mult_22/SUMB[62][28] , \mult_22/SUMB[62][29] ,
         \mult_22/SUMB[62][30] , \mult_22/SUMB[62][31] ,
         \mult_22/SUMB[62][32] , \mult_22/SUMB[62][33] ,
         \mult_22/SUMB[62][34] , \mult_22/SUMB[62][35] ,
         \mult_22/SUMB[62][36] , \mult_22/SUMB[62][37] ,
         \mult_22/SUMB[62][38] , \mult_22/SUMB[62][39] ,
         \mult_22/SUMB[62][40] , \mult_22/SUMB[62][41] ,
         \mult_22/SUMB[62][42] , \mult_22/SUMB[62][43] ,
         \mult_22/SUMB[62][44] , \mult_22/SUMB[62][45] ,
         \mult_22/SUMB[62][46] , \mult_22/SUMB[62][47] ,
         \mult_22/SUMB[62][48] , \mult_22/SUMB[62][49] ,
         \mult_22/SUMB[62][50] , \mult_22/SUMB[62][51] ,
         \mult_22/SUMB[62][52] , \mult_22/SUMB[62][53] ,
         \mult_22/SUMB[62][54] , \mult_22/SUMB[62][55] ,
         \mult_22/SUMB[62][56] , \mult_22/SUMB[62][57] ,
         \mult_22/SUMB[62][58] , \mult_22/SUMB[62][59] ,
         \mult_22/SUMB[62][60] , \mult_22/SUMB[62][61] ,
         \mult_22/SUMB[62][62] , \mult_22/SUMB[63][1] , \mult_22/SUMB[63][2] ,
         \mult_22/SUMB[63][3] , \mult_22/SUMB[63][4] , \mult_22/SUMB[63][5] ,
         \mult_22/SUMB[63][6] , \mult_22/SUMB[63][7] , \mult_22/SUMB[63][8] ,
         \mult_22/SUMB[63][9] , \mult_22/SUMB[63][10] , \mult_22/SUMB[63][11] ,
         \mult_22/SUMB[63][12] , \mult_22/SUMB[63][13] ,
         \mult_22/SUMB[63][14] , \mult_22/SUMB[63][15] ,
         \mult_22/SUMB[63][16] , \mult_22/SUMB[63][17] ,
         \mult_22/SUMB[63][18] , \mult_22/SUMB[63][19] ,
         \mult_22/SUMB[63][20] , \mult_22/SUMB[63][21] ,
         \mult_22/SUMB[63][22] , \mult_22/SUMB[63][23] ,
         \mult_22/SUMB[63][24] , \mult_22/SUMB[63][25] ,
         \mult_22/SUMB[63][26] , \mult_22/SUMB[63][27] ,
         \mult_22/SUMB[63][28] , \mult_22/SUMB[63][29] ,
         \mult_22/SUMB[63][30] , \mult_22/SUMB[63][31] ,
         \mult_22/SUMB[63][32] , \mult_22/SUMB[63][33] ,
         \mult_22/SUMB[63][34] , \mult_22/SUMB[63][35] ,
         \mult_22/SUMB[63][36] , \mult_22/SUMB[63][37] ,
         \mult_22/SUMB[63][38] , \mult_22/SUMB[63][39] ,
         \mult_22/SUMB[63][40] , \mult_22/SUMB[63][41] ,
         \mult_22/SUMB[63][42] , \mult_22/SUMB[63][43] ,
         \mult_22/SUMB[63][44] , \mult_22/SUMB[63][45] ,
         \mult_22/SUMB[63][46] , \mult_22/SUMB[63][47] ,
         \mult_22/SUMB[63][48] , \mult_22/SUMB[63][49] ,
         \mult_22/SUMB[63][50] , \mult_22/SUMB[63][51] ,
         \mult_22/SUMB[63][52] , \mult_22/SUMB[63][53] ,
         \mult_22/SUMB[63][54] , \mult_22/SUMB[63][55] ,
         \mult_22/SUMB[63][56] , \mult_22/SUMB[63][57] ,
         \mult_22/SUMB[63][58] , \mult_22/SUMB[63][59] ,
         \mult_22/SUMB[63][60] , \mult_22/SUMB[63][61] ,
         \mult_22/SUMB[63][62] , \mult_22/CARRYB[56][0] ,
         \mult_22/CARRYB[56][1] , \mult_22/CARRYB[56][2] ,
         \mult_22/CARRYB[56][3] , \mult_22/CARRYB[56][4] ,
         \mult_22/CARRYB[56][5] , \mult_22/CARRYB[56][6] ,
         \mult_22/CARRYB[56][7] , \mult_22/CARRYB[56][8] ,
         \mult_22/CARRYB[56][9] , \mult_22/CARRYB[56][10] ,
         \mult_22/CARRYB[56][11] , \mult_22/CARRYB[56][12] ,
         \mult_22/CARRYB[56][13] , \mult_22/CARRYB[56][14] ,
         \mult_22/CARRYB[56][15] , \mult_22/CARRYB[56][16] ,
         \mult_22/CARRYB[56][17] , \mult_22/CARRYB[56][18] ,
         \mult_22/CARRYB[56][19] , \mult_22/CARRYB[56][20] ,
         \mult_22/CARRYB[56][21] , \mult_22/CARRYB[56][22] ,
         \mult_22/CARRYB[56][23] , \mult_22/CARRYB[56][24] ,
         \mult_22/CARRYB[56][25] , \mult_22/CARRYB[56][26] ,
         \mult_22/CARRYB[56][27] , \mult_22/CARRYB[56][28] ,
         \mult_22/CARRYB[56][29] , \mult_22/CARRYB[56][30] ,
         \mult_22/CARRYB[56][31] , \mult_22/CARRYB[56][32] ,
         \mult_22/CARRYB[56][33] , \mult_22/CARRYB[56][34] ,
         \mult_22/CARRYB[56][35] , \mult_22/CARRYB[56][36] ,
         \mult_22/CARRYB[56][37] , \mult_22/CARRYB[56][38] ,
         \mult_22/CARRYB[56][39] , \mult_22/CARRYB[56][40] ,
         \mult_22/CARRYB[56][41] , \mult_22/CARRYB[56][42] ,
         \mult_22/CARRYB[56][43] , \mult_22/CARRYB[56][44] ,
         \mult_22/CARRYB[56][45] , \mult_22/CARRYB[56][46] ,
         \mult_22/CARRYB[56][47] , \mult_22/CARRYB[56][48] ,
         \mult_22/CARRYB[56][49] , \mult_22/CARRYB[56][50] ,
         \mult_22/CARRYB[56][51] , \mult_22/CARRYB[56][52] ,
         \mult_22/CARRYB[56][53] , \mult_22/CARRYB[56][54] ,
         \mult_22/CARRYB[56][55] , \mult_22/CARRYB[56][56] ,
         \mult_22/CARRYB[56][57] , \mult_22/CARRYB[56][58] ,
         \mult_22/CARRYB[56][59] , \mult_22/CARRYB[56][60] ,
         \mult_22/CARRYB[56][61] , \mult_22/CARRYB[56][62] ,
         \mult_22/CARRYB[57][0] , \mult_22/CARRYB[57][1] ,
         \mult_22/CARRYB[57][2] , \mult_22/CARRYB[57][3] ,
         \mult_22/CARRYB[57][4] , \mult_22/CARRYB[57][5] ,
         \mult_22/CARRYB[57][6] , \mult_22/CARRYB[57][7] ,
         \mult_22/CARRYB[57][8] , \mult_22/CARRYB[57][9] ,
         \mult_22/CARRYB[57][10] , \mult_22/CARRYB[57][11] ,
         \mult_22/CARRYB[57][12] , \mult_22/CARRYB[57][13] ,
         \mult_22/CARRYB[57][14] , \mult_22/CARRYB[57][15] ,
         \mult_22/CARRYB[57][16] , \mult_22/CARRYB[57][17] ,
         \mult_22/CARRYB[57][18] , \mult_22/CARRYB[57][19] ,
         \mult_22/CARRYB[57][20] , \mult_22/CARRYB[57][21] ,
         \mult_22/CARRYB[57][22] , \mult_22/CARRYB[57][23] ,
         \mult_22/CARRYB[57][24] , \mult_22/CARRYB[57][25] ,
         \mult_22/CARRYB[57][26] , \mult_22/CARRYB[57][27] ,
         \mult_22/CARRYB[57][28] , \mult_22/CARRYB[57][29] ,
         \mult_22/CARRYB[57][30] , \mult_22/CARRYB[57][31] ,
         \mult_22/CARRYB[57][32] , \mult_22/CARRYB[57][33] ,
         \mult_22/CARRYB[57][34] , \mult_22/CARRYB[57][35] ,
         \mult_22/CARRYB[57][36] , \mult_22/CARRYB[57][37] ,
         \mult_22/CARRYB[57][38] , \mult_22/CARRYB[57][39] ,
         \mult_22/CARRYB[57][40] , \mult_22/CARRYB[57][41] ,
         \mult_22/CARRYB[57][42] , \mult_22/CARRYB[57][43] ,
         \mult_22/CARRYB[57][44] , \mult_22/CARRYB[57][45] ,
         \mult_22/CARRYB[57][46] , \mult_22/CARRYB[57][47] ,
         \mult_22/CARRYB[57][48] , \mult_22/CARRYB[57][49] ,
         \mult_22/CARRYB[57][50] , \mult_22/CARRYB[57][51] ,
         \mult_22/CARRYB[57][52] , \mult_22/CARRYB[57][53] ,
         \mult_22/CARRYB[57][54] , \mult_22/CARRYB[57][55] ,
         \mult_22/CARRYB[57][56] , \mult_22/CARRYB[57][57] ,
         \mult_22/CARRYB[57][58] , \mult_22/CARRYB[57][59] ,
         \mult_22/CARRYB[57][60] , \mult_22/CARRYB[57][61] ,
         \mult_22/CARRYB[57][62] , \mult_22/CARRYB[58][0] ,
         \mult_22/CARRYB[58][1] , \mult_22/CARRYB[58][2] ,
         \mult_22/CARRYB[58][3] , \mult_22/CARRYB[58][4] ,
         \mult_22/CARRYB[58][5] , \mult_22/CARRYB[58][6] ,
         \mult_22/CARRYB[58][7] , \mult_22/CARRYB[58][8] ,
         \mult_22/CARRYB[58][9] , \mult_22/CARRYB[58][10] ,
         \mult_22/CARRYB[58][11] , \mult_22/CARRYB[58][12] ,
         \mult_22/CARRYB[58][13] , \mult_22/CARRYB[58][14] ,
         \mult_22/CARRYB[58][15] , \mult_22/CARRYB[58][16] ,
         \mult_22/CARRYB[58][17] , \mult_22/CARRYB[58][18] ,
         \mult_22/CARRYB[58][19] , \mult_22/CARRYB[58][20] ,
         \mult_22/CARRYB[58][21] , \mult_22/CARRYB[58][22] ,
         \mult_22/CARRYB[58][23] , \mult_22/CARRYB[58][24] ,
         \mult_22/CARRYB[58][25] , \mult_22/CARRYB[58][26] ,
         \mult_22/CARRYB[58][27] , \mult_22/CARRYB[58][28] ,
         \mult_22/CARRYB[58][29] , \mult_22/CARRYB[58][30] ,
         \mult_22/CARRYB[58][31] , \mult_22/CARRYB[58][32] ,
         \mult_22/CARRYB[58][33] , \mult_22/CARRYB[58][34] ,
         \mult_22/CARRYB[58][35] , \mult_22/CARRYB[58][36] ,
         \mult_22/CARRYB[58][37] , \mult_22/CARRYB[58][38] ,
         \mult_22/CARRYB[58][39] , \mult_22/CARRYB[58][40] ,
         \mult_22/CARRYB[58][41] , \mult_22/CARRYB[58][42] ,
         \mult_22/CARRYB[58][43] , \mult_22/CARRYB[58][44] ,
         \mult_22/CARRYB[58][45] , \mult_22/CARRYB[58][46] ,
         \mult_22/CARRYB[58][47] , \mult_22/CARRYB[58][48] ,
         \mult_22/CARRYB[58][49] , \mult_22/CARRYB[58][50] ,
         \mult_22/CARRYB[58][51] , \mult_22/CARRYB[58][52] ,
         \mult_22/CARRYB[58][53] , \mult_22/CARRYB[58][54] ,
         \mult_22/CARRYB[58][55] , \mult_22/CARRYB[58][56] ,
         \mult_22/CARRYB[58][57] , \mult_22/CARRYB[58][58] ,
         \mult_22/CARRYB[58][59] , \mult_22/CARRYB[58][60] ,
         \mult_22/CARRYB[58][61] , \mult_22/CARRYB[58][62] ,
         \mult_22/CARRYB[59][0] , \mult_22/CARRYB[59][1] ,
         \mult_22/CARRYB[59][2] , \mult_22/CARRYB[59][3] ,
         \mult_22/CARRYB[59][4] , \mult_22/CARRYB[59][5] ,
         \mult_22/CARRYB[59][6] , \mult_22/CARRYB[59][7] ,
         \mult_22/CARRYB[59][8] , \mult_22/CARRYB[59][9] ,
         \mult_22/CARRYB[59][10] , \mult_22/CARRYB[59][11] ,
         \mult_22/CARRYB[59][12] , \mult_22/CARRYB[59][13] ,
         \mult_22/CARRYB[59][14] , \mult_22/CARRYB[59][15] ,
         \mult_22/CARRYB[59][16] , \mult_22/CARRYB[59][17] ,
         \mult_22/CARRYB[59][18] , \mult_22/CARRYB[59][19] ,
         \mult_22/CARRYB[59][20] , \mult_22/CARRYB[59][21] ,
         \mult_22/CARRYB[59][22] , \mult_22/CARRYB[59][23] ,
         \mult_22/CARRYB[59][24] , \mult_22/CARRYB[59][25] ,
         \mult_22/CARRYB[59][26] , \mult_22/CARRYB[59][27] ,
         \mult_22/CARRYB[59][28] , \mult_22/CARRYB[59][29] ,
         \mult_22/CARRYB[59][30] , \mult_22/CARRYB[59][31] ,
         \mult_22/CARRYB[59][32] , \mult_22/CARRYB[59][33] ,
         \mult_22/CARRYB[59][34] , \mult_22/CARRYB[59][35] ,
         \mult_22/CARRYB[59][36] , \mult_22/CARRYB[59][37] ,
         \mult_22/CARRYB[59][38] , \mult_22/CARRYB[59][39] ,
         \mult_22/CARRYB[59][40] , \mult_22/CARRYB[59][41] ,
         \mult_22/CARRYB[59][42] , \mult_22/CARRYB[59][43] ,
         \mult_22/CARRYB[59][44] , \mult_22/CARRYB[59][45] ,
         \mult_22/CARRYB[59][46] , \mult_22/CARRYB[59][47] ,
         \mult_22/CARRYB[59][48] , \mult_22/CARRYB[59][49] ,
         \mult_22/CARRYB[59][50] , \mult_22/CARRYB[59][51] ,
         \mult_22/CARRYB[59][52] , \mult_22/CARRYB[59][53] ,
         \mult_22/CARRYB[59][54] , \mult_22/CARRYB[59][55] ,
         \mult_22/CARRYB[59][56] , \mult_22/CARRYB[59][57] ,
         \mult_22/CARRYB[59][58] , \mult_22/CARRYB[59][59] ,
         \mult_22/CARRYB[59][60] , \mult_22/CARRYB[59][61] ,
         \mult_22/CARRYB[59][62] , \mult_22/CARRYB[60][0] ,
         \mult_22/CARRYB[60][1] , \mult_22/CARRYB[60][2] ,
         \mult_22/CARRYB[60][3] , \mult_22/CARRYB[60][4] ,
         \mult_22/CARRYB[60][5] , \mult_22/CARRYB[60][6] ,
         \mult_22/CARRYB[60][7] , \mult_22/CARRYB[60][8] ,
         \mult_22/CARRYB[60][9] , \mult_22/CARRYB[60][10] ,
         \mult_22/CARRYB[60][11] , \mult_22/CARRYB[60][12] ,
         \mult_22/CARRYB[60][13] , \mult_22/CARRYB[60][14] ,
         \mult_22/CARRYB[60][15] , \mult_22/CARRYB[60][16] ,
         \mult_22/CARRYB[60][17] , \mult_22/CARRYB[60][18] ,
         \mult_22/CARRYB[60][19] , \mult_22/CARRYB[60][20] ,
         \mult_22/CARRYB[60][21] , \mult_22/CARRYB[60][22] ,
         \mult_22/CARRYB[60][23] , \mult_22/CARRYB[60][24] ,
         \mult_22/CARRYB[60][25] , \mult_22/CARRYB[60][26] ,
         \mult_22/CARRYB[60][27] , \mult_22/CARRYB[60][28] ,
         \mult_22/CARRYB[60][29] , \mult_22/CARRYB[60][30] ,
         \mult_22/CARRYB[60][31] , \mult_22/CARRYB[60][32] ,
         \mult_22/CARRYB[60][33] , \mult_22/CARRYB[60][34] ,
         \mult_22/CARRYB[60][35] , \mult_22/CARRYB[60][36] ,
         \mult_22/CARRYB[60][37] , \mult_22/CARRYB[60][38] ,
         \mult_22/CARRYB[60][39] , \mult_22/CARRYB[60][40] ,
         \mult_22/CARRYB[60][41] , \mult_22/CARRYB[60][42] ,
         \mult_22/CARRYB[60][43] , \mult_22/CARRYB[60][44] ,
         \mult_22/CARRYB[60][45] , \mult_22/CARRYB[60][46] ,
         \mult_22/CARRYB[60][47] , \mult_22/CARRYB[60][48] ,
         \mult_22/CARRYB[60][49] , \mult_22/CARRYB[60][50] ,
         \mult_22/CARRYB[60][51] , \mult_22/CARRYB[60][52] ,
         \mult_22/CARRYB[60][53] , \mult_22/CARRYB[60][54] ,
         \mult_22/CARRYB[60][55] , \mult_22/CARRYB[60][56] ,
         \mult_22/CARRYB[60][57] , \mult_22/CARRYB[60][58] ,
         \mult_22/CARRYB[60][59] , \mult_22/CARRYB[60][60] ,
         \mult_22/CARRYB[60][61] , \mult_22/CARRYB[60][62] ,
         \mult_22/CARRYB[61][0] , \mult_22/CARRYB[61][1] ,
         \mult_22/CARRYB[61][2] , \mult_22/CARRYB[61][3] ,
         \mult_22/CARRYB[61][4] , \mult_22/CARRYB[61][5] ,
         \mult_22/CARRYB[61][6] , \mult_22/CARRYB[61][7] ,
         \mult_22/CARRYB[61][8] , \mult_22/CARRYB[61][9] ,
         \mult_22/CARRYB[61][10] , \mult_22/CARRYB[61][11] ,
         \mult_22/CARRYB[61][12] , \mult_22/CARRYB[61][13] ,
         \mult_22/CARRYB[61][14] , \mult_22/CARRYB[61][15] ,
         \mult_22/CARRYB[61][16] , \mult_22/CARRYB[61][17] ,
         \mult_22/CARRYB[61][18] , \mult_22/CARRYB[61][19] ,
         \mult_22/CARRYB[61][20] , \mult_22/CARRYB[61][21] ,
         \mult_22/CARRYB[61][22] , \mult_22/CARRYB[61][23] ,
         \mult_22/CARRYB[61][24] , \mult_22/CARRYB[61][25] ,
         \mult_22/CARRYB[61][26] , \mult_22/CARRYB[61][27] ,
         \mult_22/CARRYB[61][28] , \mult_22/CARRYB[61][29] ,
         \mult_22/CARRYB[61][30] , \mult_22/CARRYB[61][31] ,
         \mult_22/CARRYB[61][32] , \mult_22/CARRYB[61][33] ,
         \mult_22/CARRYB[61][34] , \mult_22/CARRYB[61][35] ,
         \mult_22/CARRYB[61][36] , \mult_22/CARRYB[61][37] ,
         \mult_22/CARRYB[61][38] , \mult_22/CARRYB[61][39] ,
         \mult_22/CARRYB[61][40] , \mult_22/CARRYB[61][41] ,
         \mult_22/CARRYB[61][42] , \mult_22/CARRYB[61][43] ,
         \mult_22/CARRYB[61][44] , \mult_22/CARRYB[61][45] ,
         \mult_22/CARRYB[61][46] , \mult_22/CARRYB[61][47] ,
         \mult_22/CARRYB[61][48] , \mult_22/CARRYB[61][49] ,
         \mult_22/CARRYB[61][50] , \mult_22/CARRYB[61][51] ,
         \mult_22/CARRYB[61][52] , \mult_22/CARRYB[61][53] ,
         \mult_22/CARRYB[61][54] , \mult_22/CARRYB[61][55] ,
         \mult_22/CARRYB[61][56] , \mult_22/CARRYB[61][57] ,
         \mult_22/CARRYB[61][58] , \mult_22/CARRYB[61][59] ,
         \mult_22/CARRYB[61][60] , \mult_22/CARRYB[61][61] ,
         \mult_22/CARRYB[61][62] , \mult_22/CARRYB[62][0] ,
         \mult_22/CARRYB[62][1] , \mult_22/CARRYB[62][2] ,
         \mult_22/CARRYB[62][3] , \mult_22/CARRYB[62][4] ,
         \mult_22/CARRYB[62][5] , \mult_22/CARRYB[62][6] ,
         \mult_22/CARRYB[62][7] , \mult_22/CARRYB[62][8] ,
         \mult_22/CARRYB[62][9] , \mult_22/CARRYB[62][10] ,
         \mult_22/CARRYB[62][11] , \mult_22/CARRYB[62][12] ,
         \mult_22/CARRYB[62][13] , \mult_22/CARRYB[62][14] ,
         \mult_22/CARRYB[62][15] , \mult_22/CARRYB[62][16] ,
         \mult_22/CARRYB[62][17] , \mult_22/CARRYB[62][18] ,
         \mult_22/CARRYB[62][19] , \mult_22/CARRYB[62][20] ,
         \mult_22/CARRYB[62][21] , \mult_22/CARRYB[62][22] ,
         \mult_22/CARRYB[62][23] , \mult_22/CARRYB[62][24] ,
         \mult_22/CARRYB[62][25] , \mult_22/CARRYB[62][26] ,
         \mult_22/CARRYB[62][27] , \mult_22/CARRYB[62][28] ,
         \mult_22/CARRYB[62][29] , \mult_22/CARRYB[62][30] ,
         \mult_22/CARRYB[62][31] , \mult_22/CARRYB[62][32] ,
         \mult_22/CARRYB[62][33] , \mult_22/CARRYB[62][34] ,
         \mult_22/CARRYB[62][35] , \mult_22/CARRYB[62][36] ,
         \mult_22/CARRYB[62][37] , \mult_22/CARRYB[62][38] ,
         \mult_22/CARRYB[62][39] , \mult_22/CARRYB[62][40] ,
         \mult_22/CARRYB[62][41] , \mult_22/CARRYB[62][42] ,
         \mult_22/CARRYB[62][43] , \mult_22/CARRYB[62][44] ,
         \mult_22/CARRYB[62][45] , \mult_22/CARRYB[62][46] ,
         \mult_22/CARRYB[62][47] , \mult_22/CARRYB[62][48] ,
         \mult_22/CARRYB[62][49] , \mult_22/CARRYB[62][50] ,
         \mult_22/CARRYB[62][51] , \mult_22/CARRYB[62][52] ,
         \mult_22/CARRYB[62][53] , \mult_22/CARRYB[62][54] ,
         \mult_22/CARRYB[62][55] , \mult_22/CARRYB[62][56] ,
         \mult_22/CARRYB[62][57] , \mult_22/CARRYB[62][58] ,
         \mult_22/CARRYB[62][59] , \mult_22/CARRYB[62][60] ,
         \mult_22/CARRYB[62][61] , \mult_22/CARRYB[62][62] ,
         \mult_22/CARRYB[63][0] , \mult_22/CARRYB[63][1] ,
         \mult_22/CARRYB[63][2] , \mult_22/CARRYB[63][3] ,
         \mult_22/CARRYB[63][4] , \mult_22/CARRYB[63][5] ,
         \mult_22/CARRYB[63][6] , \mult_22/CARRYB[63][7] ,
         \mult_22/CARRYB[63][8] , \mult_22/CARRYB[63][9] ,
         \mult_22/CARRYB[63][10] , \mult_22/CARRYB[63][11] ,
         \mult_22/CARRYB[63][12] , \mult_22/CARRYB[63][13] ,
         \mult_22/CARRYB[63][14] , \mult_22/CARRYB[63][15] ,
         \mult_22/CARRYB[63][16] , \mult_22/CARRYB[63][17] ,
         \mult_22/CARRYB[63][18] , \mult_22/CARRYB[63][19] ,
         \mult_22/CARRYB[63][20] , \mult_22/CARRYB[63][21] ,
         \mult_22/CARRYB[63][22] , \mult_22/CARRYB[63][23] ,
         \mult_22/CARRYB[63][24] , \mult_22/CARRYB[63][25] ,
         \mult_22/CARRYB[63][26] , \mult_22/CARRYB[63][27] ,
         \mult_22/CARRYB[63][28] , \mult_22/CARRYB[63][29] ,
         \mult_22/CARRYB[63][30] , \mult_22/CARRYB[63][31] ,
         \mult_22/CARRYB[63][32] , \mult_22/CARRYB[63][33] ,
         \mult_22/CARRYB[63][34] , \mult_22/CARRYB[63][35] ,
         \mult_22/CARRYB[63][36] , \mult_22/CARRYB[63][37] ,
         \mult_22/CARRYB[63][38] , \mult_22/CARRYB[63][39] ,
         \mult_22/CARRYB[63][40] , \mult_22/CARRYB[63][41] ,
         \mult_22/CARRYB[63][42] , \mult_22/CARRYB[63][43] ,
         \mult_22/CARRYB[63][44] , \mult_22/CARRYB[63][45] ,
         \mult_22/CARRYB[63][46] , \mult_22/CARRYB[63][47] ,
         \mult_22/CARRYB[63][48] , \mult_22/CARRYB[63][49] ,
         \mult_22/CARRYB[63][50] , \mult_22/CARRYB[63][51] ,
         \mult_22/CARRYB[63][52] , \mult_22/CARRYB[63][53] ,
         \mult_22/CARRYB[63][54] , \mult_22/CARRYB[63][55] ,
         \mult_22/CARRYB[63][56] , \mult_22/CARRYB[63][57] ,
         \mult_22/CARRYB[63][58] , \mult_22/CARRYB[63][59] ,
         \mult_22/CARRYB[63][60] , \mult_22/CARRYB[63][61] ,
         \mult_22/CARRYB[63][62] , \mult_22/SUMB[48][1] ,
         \mult_22/SUMB[48][2] , \mult_22/SUMB[48][3] , \mult_22/SUMB[48][4] ,
         \mult_22/SUMB[48][5] , \mult_22/SUMB[48][6] , \mult_22/SUMB[48][7] ,
         \mult_22/SUMB[48][8] , \mult_22/SUMB[48][9] , \mult_22/SUMB[48][10] ,
         \mult_22/SUMB[48][11] , \mult_22/SUMB[48][12] ,
         \mult_22/SUMB[48][13] , \mult_22/SUMB[48][14] ,
         \mult_22/SUMB[48][15] , \mult_22/SUMB[48][16] ,
         \mult_22/SUMB[48][17] , \mult_22/SUMB[48][18] ,
         \mult_22/SUMB[48][19] , \mult_22/SUMB[48][20] ,
         \mult_22/SUMB[48][21] , \mult_22/SUMB[48][22] ,
         \mult_22/SUMB[48][23] , \mult_22/SUMB[48][24] ,
         \mult_22/SUMB[48][25] , \mult_22/SUMB[48][26] ,
         \mult_22/SUMB[48][27] , \mult_22/SUMB[48][28] ,
         \mult_22/SUMB[48][29] , \mult_22/SUMB[48][30] ,
         \mult_22/SUMB[48][31] , \mult_22/SUMB[48][32] ,
         \mult_22/SUMB[48][33] , \mult_22/SUMB[48][34] ,
         \mult_22/SUMB[48][35] , \mult_22/SUMB[48][36] ,
         \mult_22/SUMB[48][37] , \mult_22/SUMB[48][38] ,
         \mult_22/SUMB[48][39] , \mult_22/SUMB[48][40] ,
         \mult_22/SUMB[48][41] , \mult_22/SUMB[48][42] ,
         \mult_22/SUMB[48][43] , \mult_22/SUMB[48][44] ,
         \mult_22/SUMB[48][45] , \mult_22/SUMB[48][46] ,
         \mult_22/SUMB[48][47] , \mult_22/SUMB[48][48] ,
         \mult_22/SUMB[48][49] , \mult_22/SUMB[48][50] ,
         \mult_22/SUMB[48][51] , \mult_22/SUMB[48][52] ,
         \mult_22/SUMB[48][53] , \mult_22/SUMB[48][54] ,
         \mult_22/SUMB[48][55] , \mult_22/SUMB[48][56] ,
         \mult_22/SUMB[48][57] , \mult_22/SUMB[48][58] ,
         \mult_22/SUMB[48][59] , \mult_22/SUMB[48][60] ,
         \mult_22/SUMB[48][61] , \mult_22/SUMB[48][62] , \mult_22/SUMB[49][1] ,
         \mult_22/SUMB[49][2] , \mult_22/SUMB[49][3] , \mult_22/SUMB[49][4] ,
         \mult_22/SUMB[49][5] , \mult_22/SUMB[49][6] , \mult_22/SUMB[49][7] ,
         \mult_22/SUMB[49][8] , \mult_22/SUMB[49][9] , \mult_22/SUMB[49][10] ,
         \mult_22/SUMB[49][11] , \mult_22/SUMB[49][12] ,
         \mult_22/SUMB[49][13] , \mult_22/SUMB[49][14] ,
         \mult_22/SUMB[49][15] , \mult_22/SUMB[49][16] ,
         \mult_22/SUMB[49][17] , \mult_22/SUMB[49][18] ,
         \mult_22/SUMB[49][19] , \mult_22/SUMB[49][20] ,
         \mult_22/SUMB[49][21] , \mult_22/SUMB[49][22] ,
         \mult_22/SUMB[49][23] , \mult_22/SUMB[49][24] ,
         \mult_22/SUMB[49][25] , \mult_22/SUMB[49][26] ,
         \mult_22/SUMB[49][27] , \mult_22/SUMB[49][28] ,
         \mult_22/SUMB[49][29] , \mult_22/SUMB[49][30] ,
         \mult_22/SUMB[49][31] , \mult_22/SUMB[49][32] ,
         \mult_22/SUMB[49][33] , \mult_22/SUMB[49][34] ,
         \mult_22/SUMB[49][35] , \mult_22/SUMB[49][36] ,
         \mult_22/SUMB[49][37] , \mult_22/SUMB[49][38] ,
         \mult_22/SUMB[49][39] , \mult_22/SUMB[49][40] ,
         \mult_22/SUMB[49][41] , \mult_22/SUMB[49][42] ,
         \mult_22/SUMB[49][43] , \mult_22/SUMB[49][44] ,
         \mult_22/SUMB[49][45] , \mult_22/SUMB[49][46] ,
         \mult_22/SUMB[49][47] , \mult_22/SUMB[49][48] ,
         \mult_22/SUMB[49][49] , \mult_22/SUMB[49][50] ,
         \mult_22/SUMB[49][51] , \mult_22/SUMB[49][52] ,
         \mult_22/SUMB[49][53] , \mult_22/SUMB[49][54] ,
         \mult_22/SUMB[49][55] , \mult_22/SUMB[49][56] ,
         \mult_22/SUMB[49][57] , \mult_22/SUMB[49][58] ,
         \mult_22/SUMB[49][59] , \mult_22/SUMB[49][60] ,
         \mult_22/SUMB[49][61] , \mult_22/SUMB[49][62] , \mult_22/SUMB[50][1] ,
         \mult_22/SUMB[50][2] , \mult_22/SUMB[50][3] , \mult_22/SUMB[50][4] ,
         \mult_22/SUMB[50][5] , \mult_22/SUMB[50][6] , \mult_22/SUMB[50][7] ,
         \mult_22/SUMB[50][8] , \mult_22/SUMB[50][9] , \mult_22/SUMB[50][10] ,
         \mult_22/SUMB[50][11] , \mult_22/SUMB[50][12] ,
         \mult_22/SUMB[50][13] , \mult_22/SUMB[50][14] ,
         \mult_22/SUMB[50][15] , \mult_22/SUMB[50][16] ,
         \mult_22/SUMB[50][17] , \mult_22/SUMB[50][18] ,
         \mult_22/SUMB[50][19] , \mult_22/SUMB[50][20] ,
         \mult_22/SUMB[50][21] , \mult_22/SUMB[50][22] ,
         \mult_22/SUMB[50][23] , \mult_22/SUMB[50][24] ,
         \mult_22/SUMB[50][25] , \mult_22/SUMB[50][26] ,
         \mult_22/SUMB[50][27] , \mult_22/SUMB[50][28] ,
         \mult_22/SUMB[50][29] , \mult_22/SUMB[50][30] ,
         \mult_22/SUMB[50][31] , \mult_22/SUMB[50][32] ,
         \mult_22/SUMB[50][33] , \mult_22/SUMB[50][34] ,
         \mult_22/SUMB[50][35] , \mult_22/SUMB[50][36] ,
         \mult_22/SUMB[50][37] , \mult_22/SUMB[50][38] ,
         \mult_22/SUMB[50][39] , \mult_22/SUMB[50][40] ,
         \mult_22/SUMB[50][41] , \mult_22/SUMB[50][42] ,
         \mult_22/SUMB[50][43] , \mult_22/SUMB[50][44] ,
         \mult_22/SUMB[50][45] , \mult_22/SUMB[50][46] ,
         \mult_22/SUMB[50][47] , \mult_22/SUMB[50][48] ,
         \mult_22/SUMB[50][49] , \mult_22/SUMB[50][50] ,
         \mult_22/SUMB[50][51] , \mult_22/SUMB[50][52] ,
         \mult_22/SUMB[50][53] , \mult_22/SUMB[50][54] ,
         \mult_22/SUMB[50][55] , \mult_22/SUMB[50][56] ,
         \mult_22/SUMB[50][57] , \mult_22/SUMB[50][58] ,
         \mult_22/SUMB[50][59] , \mult_22/SUMB[50][60] ,
         \mult_22/SUMB[50][61] , \mult_22/SUMB[50][62] , \mult_22/SUMB[51][1] ,
         \mult_22/SUMB[51][2] , \mult_22/SUMB[51][3] , \mult_22/SUMB[51][4] ,
         \mult_22/SUMB[51][5] , \mult_22/SUMB[51][6] , \mult_22/SUMB[51][7] ,
         \mult_22/SUMB[51][8] , \mult_22/SUMB[51][9] , \mult_22/SUMB[51][10] ,
         \mult_22/SUMB[51][11] , \mult_22/SUMB[51][12] ,
         \mult_22/SUMB[51][13] , \mult_22/SUMB[51][14] ,
         \mult_22/SUMB[51][15] , \mult_22/SUMB[51][16] ,
         \mult_22/SUMB[51][17] , \mult_22/SUMB[51][18] ,
         \mult_22/SUMB[51][19] , \mult_22/SUMB[51][20] ,
         \mult_22/SUMB[51][21] , \mult_22/SUMB[51][22] ,
         \mult_22/SUMB[51][23] , \mult_22/SUMB[51][24] ,
         \mult_22/SUMB[51][25] , \mult_22/SUMB[51][26] ,
         \mult_22/SUMB[51][27] , \mult_22/SUMB[51][28] ,
         \mult_22/SUMB[51][29] , \mult_22/SUMB[51][30] ,
         \mult_22/SUMB[51][31] , \mult_22/SUMB[51][32] ,
         \mult_22/SUMB[51][33] , \mult_22/SUMB[51][34] ,
         \mult_22/SUMB[51][35] , \mult_22/SUMB[51][36] ,
         \mult_22/SUMB[51][37] , \mult_22/SUMB[51][38] ,
         \mult_22/SUMB[51][39] , \mult_22/SUMB[51][40] ,
         \mult_22/SUMB[51][41] , \mult_22/SUMB[51][42] ,
         \mult_22/SUMB[51][43] , \mult_22/SUMB[51][44] ,
         \mult_22/SUMB[51][45] , \mult_22/SUMB[51][46] ,
         \mult_22/SUMB[51][47] , \mult_22/SUMB[51][48] ,
         \mult_22/SUMB[51][49] , \mult_22/SUMB[51][50] ,
         \mult_22/SUMB[51][51] , \mult_22/SUMB[51][52] ,
         \mult_22/SUMB[51][53] , \mult_22/SUMB[51][54] ,
         \mult_22/SUMB[51][55] , \mult_22/SUMB[51][56] ,
         \mult_22/SUMB[51][57] , \mult_22/SUMB[51][58] ,
         \mult_22/SUMB[51][59] , \mult_22/SUMB[51][60] ,
         \mult_22/SUMB[51][61] , \mult_22/SUMB[51][62] , \mult_22/SUMB[52][1] ,
         \mult_22/SUMB[52][2] , \mult_22/SUMB[52][3] , \mult_22/SUMB[52][4] ,
         \mult_22/SUMB[52][5] , \mult_22/SUMB[52][6] , \mult_22/SUMB[52][7] ,
         \mult_22/SUMB[52][8] , \mult_22/SUMB[52][9] , \mult_22/SUMB[52][10] ,
         \mult_22/SUMB[52][11] , \mult_22/SUMB[52][12] ,
         \mult_22/SUMB[52][13] , \mult_22/SUMB[52][14] ,
         \mult_22/SUMB[52][15] , \mult_22/SUMB[52][16] ,
         \mult_22/SUMB[52][17] , \mult_22/SUMB[52][18] ,
         \mult_22/SUMB[52][19] , \mult_22/SUMB[52][20] ,
         \mult_22/SUMB[52][21] , \mult_22/SUMB[52][22] ,
         \mult_22/SUMB[52][23] , \mult_22/SUMB[52][24] ,
         \mult_22/SUMB[52][25] , \mult_22/SUMB[52][26] ,
         \mult_22/SUMB[52][27] , \mult_22/SUMB[52][28] ,
         \mult_22/SUMB[52][29] , \mult_22/SUMB[52][30] ,
         \mult_22/SUMB[52][31] , \mult_22/SUMB[52][32] ,
         \mult_22/SUMB[52][33] , \mult_22/SUMB[52][34] ,
         \mult_22/SUMB[52][35] , \mult_22/SUMB[52][36] ,
         \mult_22/SUMB[52][37] , \mult_22/SUMB[52][38] ,
         \mult_22/SUMB[52][39] , \mult_22/SUMB[52][40] ,
         \mult_22/SUMB[52][41] , \mult_22/SUMB[52][42] ,
         \mult_22/SUMB[52][43] , \mult_22/SUMB[52][44] ,
         \mult_22/SUMB[52][45] , \mult_22/SUMB[52][46] ,
         \mult_22/SUMB[52][47] , \mult_22/SUMB[52][48] ,
         \mult_22/SUMB[52][49] , \mult_22/SUMB[52][50] ,
         \mult_22/SUMB[52][51] , \mult_22/SUMB[52][52] ,
         \mult_22/SUMB[52][53] , \mult_22/SUMB[52][54] ,
         \mult_22/SUMB[52][55] , \mult_22/SUMB[52][56] ,
         \mult_22/SUMB[52][57] , \mult_22/SUMB[52][58] ,
         \mult_22/SUMB[52][59] , \mult_22/SUMB[52][60] ,
         \mult_22/SUMB[52][61] , \mult_22/SUMB[52][62] , \mult_22/SUMB[53][1] ,
         \mult_22/SUMB[53][2] , \mult_22/SUMB[53][3] , \mult_22/SUMB[53][4] ,
         \mult_22/SUMB[53][5] , \mult_22/SUMB[53][6] , \mult_22/SUMB[53][7] ,
         \mult_22/SUMB[53][8] , \mult_22/SUMB[53][9] , \mult_22/SUMB[53][10] ,
         \mult_22/SUMB[53][11] , \mult_22/SUMB[53][12] ,
         \mult_22/SUMB[53][13] , \mult_22/SUMB[53][14] ,
         \mult_22/SUMB[53][15] , \mult_22/SUMB[53][16] ,
         \mult_22/SUMB[53][17] , \mult_22/SUMB[53][18] ,
         \mult_22/SUMB[53][19] , \mult_22/SUMB[53][20] ,
         \mult_22/SUMB[53][21] , \mult_22/SUMB[53][22] ,
         \mult_22/SUMB[53][23] , \mult_22/SUMB[53][24] ,
         \mult_22/SUMB[53][25] , \mult_22/SUMB[53][26] ,
         \mult_22/SUMB[53][27] , \mult_22/SUMB[53][28] ,
         \mult_22/SUMB[53][29] , \mult_22/SUMB[53][30] ,
         \mult_22/SUMB[53][31] , \mult_22/SUMB[53][32] ,
         \mult_22/SUMB[53][33] , \mult_22/SUMB[53][34] ,
         \mult_22/SUMB[53][35] , \mult_22/SUMB[53][36] ,
         \mult_22/SUMB[53][37] , \mult_22/SUMB[53][38] ,
         \mult_22/SUMB[53][39] , \mult_22/SUMB[53][40] ,
         \mult_22/SUMB[53][41] , \mult_22/SUMB[53][42] ,
         \mult_22/SUMB[53][43] , \mult_22/SUMB[53][44] ,
         \mult_22/SUMB[53][45] , \mult_22/SUMB[53][46] ,
         \mult_22/SUMB[53][47] , \mult_22/SUMB[53][48] ,
         \mult_22/SUMB[53][49] , \mult_22/SUMB[53][50] ,
         \mult_22/SUMB[53][51] , \mult_22/SUMB[53][52] ,
         \mult_22/SUMB[53][53] , \mult_22/SUMB[53][54] ,
         \mult_22/SUMB[53][55] , \mult_22/SUMB[53][56] ,
         \mult_22/SUMB[53][57] , \mult_22/SUMB[53][58] ,
         \mult_22/SUMB[53][59] , \mult_22/SUMB[53][60] ,
         \mult_22/SUMB[53][61] , \mult_22/SUMB[53][62] , \mult_22/SUMB[54][1] ,
         \mult_22/SUMB[54][2] , \mult_22/SUMB[54][3] , \mult_22/SUMB[54][4] ,
         \mult_22/SUMB[54][5] , \mult_22/SUMB[54][6] , \mult_22/SUMB[54][7] ,
         \mult_22/SUMB[54][8] , \mult_22/SUMB[54][9] , \mult_22/SUMB[54][10] ,
         \mult_22/SUMB[54][11] , \mult_22/SUMB[54][12] ,
         \mult_22/SUMB[54][13] , \mult_22/SUMB[54][14] ,
         \mult_22/SUMB[54][15] , \mult_22/SUMB[54][16] ,
         \mult_22/SUMB[54][17] , \mult_22/SUMB[54][18] ,
         \mult_22/SUMB[54][19] , \mult_22/SUMB[54][20] ,
         \mult_22/SUMB[54][21] , \mult_22/SUMB[54][22] ,
         \mult_22/SUMB[54][23] , \mult_22/SUMB[54][24] ,
         \mult_22/SUMB[54][25] , \mult_22/SUMB[54][26] ,
         \mult_22/SUMB[54][27] , \mult_22/SUMB[54][28] ,
         \mult_22/SUMB[54][29] , \mult_22/SUMB[54][30] ,
         \mult_22/SUMB[54][31] , \mult_22/SUMB[54][32] ,
         \mult_22/SUMB[54][33] , \mult_22/SUMB[54][34] ,
         \mult_22/SUMB[54][35] , \mult_22/SUMB[54][36] ,
         \mult_22/SUMB[54][37] , \mult_22/SUMB[54][38] ,
         \mult_22/SUMB[54][39] , \mult_22/SUMB[54][40] ,
         \mult_22/SUMB[54][41] , \mult_22/SUMB[54][42] ,
         \mult_22/SUMB[54][43] , \mult_22/SUMB[54][44] ,
         \mult_22/SUMB[54][45] , \mult_22/SUMB[54][46] ,
         \mult_22/SUMB[54][47] , \mult_22/SUMB[54][48] ,
         \mult_22/SUMB[54][49] , \mult_22/SUMB[54][50] ,
         \mult_22/SUMB[54][51] , \mult_22/SUMB[54][52] ,
         \mult_22/SUMB[54][53] , \mult_22/SUMB[54][54] ,
         \mult_22/SUMB[54][55] , \mult_22/SUMB[54][56] ,
         \mult_22/SUMB[54][57] , \mult_22/SUMB[54][58] ,
         \mult_22/SUMB[54][59] , \mult_22/SUMB[54][60] ,
         \mult_22/SUMB[54][61] , \mult_22/SUMB[54][62] , \mult_22/SUMB[55][1] ,
         \mult_22/SUMB[55][2] , \mult_22/SUMB[55][3] , \mult_22/SUMB[55][4] ,
         \mult_22/SUMB[55][5] , \mult_22/SUMB[55][6] , \mult_22/SUMB[55][7] ,
         \mult_22/SUMB[55][8] , \mult_22/SUMB[55][9] , \mult_22/SUMB[55][10] ,
         \mult_22/SUMB[55][11] , \mult_22/SUMB[55][12] ,
         \mult_22/SUMB[55][13] , \mult_22/SUMB[55][14] ,
         \mult_22/SUMB[55][15] , \mult_22/SUMB[55][16] ,
         \mult_22/SUMB[55][17] , \mult_22/SUMB[55][18] ,
         \mult_22/SUMB[55][19] , \mult_22/SUMB[55][20] ,
         \mult_22/SUMB[55][21] , \mult_22/SUMB[55][22] ,
         \mult_22/SUMB[55][23] , \mult_22/SUMB[55][24] ,
         \mult_22/SUMB[55][25] , \mult_22/SUMB[55][26] ,
         \mult_22/SUMB[55][27] , \mult_22/SUMB[55][28] ,
         \mult_22/SUMB[55][29] , \mult_22/SUMB[55][30] ,
         \mult_22/SUMB[55][31] , \mult_22/SUMB[55][32] ,
         \mult_22/SUMB[55][33] , \mult_22/SUMB[55][34] ,
         \mult_22/SUMB[55][35] , \mult_22/SUMB[55][36] ,
         \mult_22/SUMB[55][37] , \mult_22/SUMB[55][38] ,
         \mult_22/SUMB[55][39] , \mult_22/SUMB[55][40] ,
         \mult_22/SUMB[55][41] , \mult_22/SUMB[55][42] ,
         \mult_22/SUMB[55][43] , \mult_22/SUMB[55][44] ,
         \mult_22/SUMB[55][45] , \mult_22/SUMB[55][46] ,
         \mult_22/SUMB[55][47] , \mult_22/SUMB[55][48] ,
         \mult_22/SUMB[55][49] , \mult_22/SUMB[55][50] ,
         \mult_22/SUMB[55][51] , \mult_22/SUMB[55][52] ,
         \mult_22/SUMB[55][53] , \mult_22/SUMB[55][54] ,
         \mult_22/SUMB[55][55] , \mult_22/SUMB[55][56] ,
         \mult_22/SUMB[55][57] , \mult_22/SUMB[55][58] ,
         \mult_22/SUMB[55][59] , \mult_22/SUMB[55][60] ,
         \mult_22/SUMB[55][61] , \mult_22/SUMB[55][62] ,
         \mult_22/CARRYB[48][0] , \mult_22/CARRYB[48][1] ,
         \mult_22/CARRYB[48][2] , \mult_22/CARRYB[48][3] ,
         \mult_22/CARRYB[48][4] , \mult_22/CARRYB[48][5] ,
         \mult_22/CARRYB[48][6] , \mult_22/CARRYB[48][7] ,
         \mult_22/CARRYB[48][8] , \mult_22/CARRYB[48][9] ,
         \mult_22/CARRYB[48][10] , \mult_22/CARRYB[48][11] ,
         \mult_22/CARRYB[48][12] , \mult_22/CARRYB[48][13] ,
         \mult_22/CARRYB[48][14] , \mult_22/CARRYB[48][15] ,
         \mult_22/CARRYB[48][16] , \mult_22/CARRYB[48][17] ,
         \mult_22/CARRYB[48][18] , \mult_22/CARRYB[48][19] ,
         \mult_22/CARRYB[48][20] , \mult_22/CARRYB[48][21] ,
         \mult_22/CARRYB[48][22] , \mult_22/CARRYB[48][23] ,
         \mult_22/CARRYB[48][24] , \mult_22/CARRYB[48][25] ,
         \mult_22/CARRYB[48][26] , \mult_22/CARRYB[48][27] ,
         \mult_22/CARRYB[48][28] , \mult_22/CARRYB[48][29] ,
         \mult_22/CARRYB[48][30] , \mult_22/CARRYB[48][31] ,
         \mult_22/CARRYB[48][32] , \mult_22/CARRYB[48][33] ,
         \mult_22/CARRYB[48][34] , \mult_22/CARRYB[48][35] ,
         \mult_22/CARRYB[48][36] , \mult_22/CARRYB[48][37] ,
         \mult_22/CARRYB[48][38] , \mult_22/CARRYB[48][39] ,
         \mult_22/CARRYB[48][40] , \mult_22/CARRYB[48][41] ,
         \mult_22/CARRYB[48][42] , \mult_22/CARRYB[48][43] ,
         \mult_22/CARRYB[48][44] , \mult_22/CARRYB[48][45] ,
         \mult_22/CARRYB[48][46] , \mult_22/CARRYB[48][47] ,
         \mult_22/CARRYB[48][48] , \mult_22/CARRYB[48][49] ,
         \mult_22/CARRYB[48][50] , \mult_22/CARRYB[48][51] ,
         \mult_22/CARRYB[48][52] , \mult_22/CARRYB[48][53] ,
         \mult_22/CARRYB[48][54] , \mult_22/CARRYB[48][55] ,
         \mult_22/CARRYB[48][56] , \mult_22/CARRYB[48][57] ,
         \mult_22/CARRYB[48][58] , \mult_22/CARRYB[48][59] ,
         \mult_22/CARRYB[48][60] , \mult_22/CARRYB[48][61] ,
         \mult_22/CARRYB[48][62] , \mult_22/CARRYB[49][0] ,
         \mult_22/CARRYB[49][1] , \mult_22/CARRYB[49][2] ,
         \mult_22/CARRYB[49][3] , \mult_22/CARRYB[49][4] ,
         \mult_22/CARRYB[49][5] , \mult_22/CARRYB[49][6] ,
         \mult_22/CARRYB[49][7] , \mult_22/CARRYB[49][8] ,
         \mult_22/CARRYB[49][9] , \mult_22/CARRYB[49][10] ,
         \mult_22/CARRYB[49][11] , \mult_22/CARRYB[49][12] ,
         \mult_22/CARRYB[49][13] , \mult_22/CARRYB[49][14] ,
         \mult_22/CARRYB[49][15] , \mult_22/CARRYB[49][16] ,
         \mult_22/CARRYB[49][17] , \mult_22/CARRYB[49][18] ,
         \mult_22/CARRYB[49][19] , \mult_22/CARRYB[49][20] ,
         \mult_22/CARRYB[49][21] , \mult_22/CARRYB[49][22] ,
         \mult_22/CARRYB[49][23] , \mult_22/CARRYB[49][24] ,
         \mult_22/CARRYB[49][25] , \mult_22/CARRYB[49][26] ,
         \mult_22/CARRYB[49][27] , \mult_22/CARRYB[49][28] ,
         \mult_22/CARRYB[49][29] , \mult_22/CARRYB[49][30] ,
         \mult_22/CARRYB[49][31] , \mult_22/CARRYB[49][32] ,
         \mult_22/CARRYB[49][33] , \mult_22/CARRYB[49][34] ,
         \mult_22/CARRYB[49][35] , \mult_22/CARRYB[49][36] ,
         \mult_22/CARRYB[49][37] , \mult_22/CARRYB[49][38] ,
         \mult_22/CARRYB[49][39] , \mult_22/CARRYB[49][40] ,
         \mult_22/CARRYB[49][41] , \mult_22/CARRYB[49][42] ,
         \mult_22/CARRYB[49][43] , \mult_22/CARRYB[49][44] ,
         \mult_22/CARRYB[49][45] , \mult_22/CARRYB[49][46] ,
         \mult_22/CARRYB[49][47] , \mult_22/CARRYB[49][48] ,
         \mult_22/CARRYB[49][49] , \mult_22/CARRYB[49][50] ,
         \mult_22/CARRYB[49][51] , \mult_22/CARRYB[49][52] ,
         \mult_22/CARRYB[49][53] , \mult_22/CARRYB[49][54] ,
         \mult_22/CARRYB[49][55] , \mult_22/CARRYB[49][56] ,
         \mult_22/CARRYB[49][57] , \mult_22/CARRYB[49][58] ,
         \mult_22/CARRYB[49][59] , \mult_22/CARRYB[49][60] ,
         \mult_22/CARRYB[49][61] , \mult_22/CARRYB[49][62] ,
         \mult_22/CARRYB[50][0] , \mult_22/CARRYB[50][1] ,
         \mult_22/CARRYB[50][2] , \mult_22/CARRYB[50][3] ,
         \mult_22/CARRYB[50][4] , \mult_22/CARRYB[50][5] ,
         \mult_22/CARRYB[50][6] , \mult_22/CARRYB[50][7] ,
         \mult_22/CARRYB[50][8] , \mult_22/CARRYB[50][9] ,
         \mult_22/CARRYB[50][10] , \mult_22/CARRYB[50][11] ,
         \mult_22/CARRYB[50][12] , \mult_22/CARRYB[50][13] ,
         \mult_22/CARRYB[50][14] , \mult_22/CARRYB[50][15] ,
         \mult_22/CARRYB[50][16] , \mult_22/CARRYB[50][17] ,
         \mult_22/CARRYB[50][18] , \mult_22/CARRYB[50][19] ,
         \mult_22/CARRYB[50][20] , \mult_22/CARRYB[50][21] ,
         \mult_22/CARRYB[50][22] , \mult_22/CARRYB[50][23] ,
         \mult_22/CARRYB[50][24] , \mult_22/CARRYB[50][25] ,
         \mult_22/CARRYB[50][26] , \mult_22/CARRYB[50][27] ,
         \mult_22/CARRYB[50][28] , \mult_22/CARRYB[50][29] ,
         \mult_22/CARRYB[50][30] , \mult_22/CARRYB[50][31] ,
         \mult_22/CARRYB[50][32] , \mult_22/CARRYB[50][33] ,
         \mult_22/CARRYB[50][34] , \mult_22/CARRYB[50][35] ,
         \mult_22/CARRYB[50][36] , \mult_22/CARRYB[50][37] ,
         \mult_22/CARRYB[50][38] , \mult_22/CARRYB[50][39] ,
         \mult_22/CARRYB[50][40] , \mult_22/CARRYB[50][41] ,
         \mult_22/CARRYB[50][42] , \mult_22/CARRYB[50][43] ,
         \mult_22/CARRYB[50][44] , \mult_22/CARRYB[50][45] ,
         \mult_22/CARRYB[50][46] , \mult_22/CARRYB[50][47] ,
         \mult_22/CARRYB[50][48] , \mult_22/CARRYB[50][49] ,
         \mult_22/CARRYB[50][50] , \mult_22/CARRYB[50][51] ,
         \mult_22/CARRYB[50][52] , \mult_22/CARRYB[50][53] ,
         \mult_22/CARRYB[50][54] , \mult_22/CARRYB[50][55] ,
         \mult_22/CARRYB[50][56] , \mult_22/CARRYB[50][57] ,
         \mult_22/CARRYB[50][58] , \mult_22/CARRYB[50][59] ,
         \mult_22/CARRYB[50][60] , \mult_22/CARRYB[50][61] ,
         \mult_22/CARRYB[50][62] , \mult_22/CARRYB[51][0] ,
         \mult_22/CARRYB[51][1] , \mult_22/CARRYB[51][2] ,
         \mult_22/CARRYB[51][3] , \mult_22/CARRYB[51][4] ,
         \mult_22/CARRYB[51][5] , \mult_22/CARRYB[51][6] ,
         \mult_22/CARRYB[51][7] , \mult_22/CARRYB[51][8] ,
         \mult_22/CARRYB[51][9] , \mult_22/CARRYB[51][10] ,
         \mult_22/CARRYB[51][11] , \mult_22/CARRYB[51][12] ,
         \mult_22/CARRYB[51][13] , \mult_22/CARRYB[51][14] ,
         \mult_22/CARRYB[51][15] , \mult_22/CARRYB[51][16] ,
         \mult_22/CARRYB[51][17] , \mult_22/CARRYB[51][18] ,
         \mult_22/CARRYB[51][19] , \mult_22/CARRYB[51][20] ,
         \mult_22/CARRYB[51][21] , \mult_22/CARRYB[51][22] ,
         \mult_22/CARRYB[51][23] , \mult_22/CARRYB[51][24] ,
         \mult_22/CARRYB[51][25] , \mult_22/CARRYB[51][26] ,
         \mult_22/CARRYB[51][27] , \mult_22/CARRYB[51][28] ,
         \mult_22/CARRYB[51][29] , \mult_22/CARRYB[51][30] ,
         \mult_22/CARRYB[51][31] , \mult_22/CARRYB[51][32] ,
         \mult_22/CARRYB[51][33] , \mult_22/CARRYB[51][34] ,
         \mult_22/CARRYB[51][35] , \mult_22/CARRYB[51][36] ,
         \mult_22/CARRYB[51][37] , \mult_22/CARRYB[51][38] ,
         \mult_22/CARRYB[51][39] , \mult_22/CARRYB[51][40] ,
         \mult_22/CARRYB[51][41] , \mult_22/CARRYB[51][42] ,
         \mult_22/CARRYB[51][43] , \mult_22/CARRYB[51][44] ,
         \mult_22/CARRYB[51][45] , \mult_22/CARRYB[51][46] ,
         \mult_22/CARRYB[51][47] , \mult_22/CARRYB[51][48] ,
         \mult_22/CARRYB[51][49] , \mult_22/CARRYB[51][50] ,
         \mult_22/CARRYB[51][51] , \mult_22/CARRYB[51][52] ,
         \mult_22/CARRYB[51][53] , \mult_22/CARRYB[51][54] ,
         \mult_22/CARRYB[51][55] , \mult_22/CARRYB[51][56] ,
         \mult_22/CARRYB[51][57] , \mult_22/CARRYB[51][58] ,
         \mult_22/CARRYB[51][59] , \mult_22/CARRYB[51][60] ,
         \mult_22/CARRYB[51][61] , \mult_22/CARRYB[51][62] ,
         \mult_22/CARRYB[52][0] , \mult_22/CARRYB[52][1] ,
         \mult_22/CARRYB[52][2] , \mult_22/CARRYB[52][3] ,
         \mult_22/CARRYB[52][4] , \mult_22/CARRYB[52][5] ,
         \mult_22/CARRYB[52][6] , \mult_22/CARRYB[52][7] ,
         \mult_22/CARRYB[52][8] , \mult_22/CARRYB[52][9] ,
         \mult_22/CARRYB[52][10] , \mult_22/CARRYB[52][11] ,
         \mult_22/CARRYB[52][12] , \mult_22/CARRYB[52][13] ,
         \mult_22/CARRYB[52][14] , \mult_22/CARRYB[52][15] ,
         \mult_22/CARRYB[52][16] , \mult_22/CARRYB[52][17] ,
         \mult_22/CARRYB[52][18] , \mult_22/CARRYB[52][19] ,
         \mult_22/CARRYB[52][20] , \mult_22/CARRYB[52][21] ,
         \mult_22/CARRYB[52][22] , \mult_22/CARRYB[52][23] ,
         \mult_22/CARRYB[52][24] , \mult_22/CARRYB[52][25] ,
         \mult_22/CARRYB[52][26] , \mult_22/CARRYB[52][27] ,
         \mult_22/CARRYB[52][28] , \mult_22/CARRYB[52][29] ,
         \mult_22/CARRYB[52][30] , \mult_22/CARRYB[52][31] ,
         \mult_22/CARRYB[52][32] , \mult_22/CARRYB[52][33] ,
         \mult_22/CARRYB[52][34] , \mult_22/CARRYB[52][35] ,
         \mult_22/CARRYB[52][36] , \mult_22/CARRYB[52][37] ,
         \mult_22/CARRYB[52][38] , \mult_22/CARRYB[52][39] ,
         \mult_22/CARRYB[52][40] , \mult_22/CARRYB[52][41] ,
         \mult_22/CARRYB[52][42] , \mult_22/CARRYB[52][43] ,
         \mult_22/CARRYB[52][44] , \mult_22/CARRYB[52][45] ,
         \mult_22/CARRYB[52][46] , \mult_22/CARRYB[52][47] ,
         \mult_22/CARRYB[52][48] , \mult_22/CARRYB[52][49] ,
         \mult_22/CARRYB[52][50] , \mult_22/CARRYB[52][51] ,
         \mult_22/CARRYB[52][52] , \mult_22/CARRYB[52][53] ,
         \mult_22/CARRYB[52][54] , \mult_22/CARRYB[52][55] ,
         \mult_22/CARRYB[52][56] , \mult_22/CARRYB[52][57] ,
         \mult_22/CARRYB[52][58] , \mult_22/CARRYB[52][59] ,
         \mult_22/CARRYB[52][60] , \mult_22/CARRYB[52][61] ,
         \mult_22/CARRYB[52][62] , \mult_22/CARRYB[53][0] ,
         \mult_22/CARRYB[53][1] , \mult_22/CARRYB[53][2] ,
         \mult_22/CARRYB[53][3] , \mult_22/CARRYB[53][4] ,
         \mult_22/CARRYB[53][5] , \mult_22/CARRYB[53][6] ,
         \mult_22/CARRYB[53][7] , \mult_22/CARRYB[53][8] ,
         \mult_22/CARRYB[53][9] , \mult_22/CARRYB[53][10] ,
         \mult_22/CARRYB[53][11] , \mult_22/CARRYB[53][12] ,
         \mult_22/CARRYB[53][13] , \mult_22/CARRYB[53][14] ,
         \mult_22/CARRYB[53][15] , \mult_22/CARRYB[53][16] ,
         \mult_22/CARRYB[53][17] , \mult_22/CARRYB[53][18] ,
         \mult_22/CARRYB[53][19] , \mult_22/CARRYB[53][20] ,
         \mult_22/CARRYB[53][21] , \mult_22/CARRYB[53][22] ,
         \mult_22/CARRYB[53][23] , \mult_22/CARRYB[53][24] ,
         \mult_22/CARRYB[53][25] , \mult_22/CARRYB[53][26] ,
         \mult_22/CARRYB[53][27] , \mult_22/CARRYB[53][28] ,
         \mult_22/CARRYB[53][29] , \mult_22/CARRYB[53][30] ,
         \mult_22/CARRYB[53][31] , \mult_22/CARRYB[53][32] ,
         \mult_22/CARRYB[53][33] , \mult_22/CARRYB[53][34] ,
         \mult_22/CARRYB[53][35] , \mult_22/CARRYB[53][36] ,
         \mult_22/CARRYB[53][37] , \mult_22/CARRYB[53][38] ,
         \mult_22/CARRYB[53][39] , \mult_22/CARRYB[53][40] ,
         \mult_22/CARRYB[53][41] , \mult_22/CARRYB[53][42] ,
         \mult_22/CARRYB[53][43] , \mult_22/CARRYB[53][44] ,
         \mult_22/CARRYB[53][45] , \mult_22/CARRYB[53][46] ,
         \mult_22/CARRYB[53][47] , \mult_22/CARRYB[53][48] ,
         \mult_22/CARRYB[53][49] , \mult_22/CARRYB[53][50] ,
         \mult_22/CARRYB[53][51] , \mult_22/CARRYB[53][52] ,
         \mult_22/CARRYB[53][53] , \mult_22/CARRYB[53][54] ,
         \mult_22/CARRYB[53][55] , \mult_22/CARRYB[53][56] ,
         \mult_22/CARRYB[53][57] , \mult_22/CARRYB[53][58] ,
         \mult_22/CARRYB[53][59] , \mult_22/CARRYB[53][60] ,
         \mult_22/CARRYB[53][61] , \mult_22/CARRYB[53][62] ,
         \mult_22/CARRYB[54][0] , \mult_22/CARRYB[54][1] ,
         \mult_22/CARRYB[54][2] , \mult_22/CARRYB[54][3] ,
         \mult_22/CARRYB[54][4] , \mult_22/CARRYB[54][5] ,
         \mult_22/CARRYB[54][6] , \mult_22/CARRYB[54][7] ,
         \mult_22/CARRYB[54][8] , \mult_22/CARRYB[54][9] ,
         \mult_22/CARRYB[54][10] , \mult_22/CARRYB[54][11] ,
         \mult_22/CARRYB[54][12] , \mult_22/CARRYB[54][13] ,
         \mult_22/CARRYB[54][14] , \mult_22/CARRYB[54][15] ,
         \mult_22/CARRYB[54][16] , \mult_22/CARRYB[54][17] ,
         \mult_22/CARRYB[54][18] , \mult_22/CARRYB[54][19] ,
         \mult_22/CARRYB[54][20] , \mult_22/CARRYB[54][21] ,
         \mult_22/CARRYB[54][22] , \mult_22/CARRYB[54][23] ,
         \mult_22/CARRYB[54][24] , \mult_22/CARRYB[54][25] ,
         \mult_22/CARRYB[54][26] , \mult_22/CARRYB[54][27] ,
         \mult_22/CARRYB[54][28] , \mult_22/CARRYB[54][29] ,
         \mult_22/CARRYB[54][30] , \mult_22/CARRYB[54][31] ,
         \mult_22/CARRYB[54][32] , \mult_22/CARRYB[54][33] ,
         \mult_22/CARRYB[54][34] , \mult_22/CARRYB[54][35] ,
         \mult_22/CARRYB[54][36] , \mult_22/CARRYB[54][37] ,
         \mult_22/CARRYB[54][38] , \mult_22/CARRYB[54][39] ,
         \mult_22/CARRYB[54][40] , \mult_22/CARRYB[54][41] ,
         \mult_22/CARRYB[54][42] , \mult_22/CARRYB[54][43] ,
         \mult_22/CARRYB[54][44] , \mult_22/CARRYB[54][45] ,
         \mult_22/CARRYB[54][46] , \mult_22/CARRYB[54][47] ,
         \mult_22/CARRYB[54][48] , \mult_22/CARRYB[54][49] ,
         \mult_22/CARRYB[54][50] , \mult_22/CARRYB[54][51] ,
         \mult_22/CARRYB[54][52] , \mult_22/CARRYB[54][53] ,
         \mult_22/CARRYB[54][54] , \mult_22/CARRYB[54][55] ,
         \mult_22/CARRYB[54][56] , \mult_22/CARRYB[54][57] ,
         \mult_22/CARRYB[54][58] , \mult_22/CARRYB[54][59] ,
         \mult_22/CARRYB[54][60] , \mult_22/CARRYB[54][61] ,
         \mult_22/CARRYB[54][62] , \mult_22/CARRYB[55][0] ,
         \mult_22/CARRYB[55][1] , \mult_22/CARRYB[55][2] ,
         \mult_22/CARRYB[55][3] , \mult_22/CARRYB[55][4] ,
         \mult_22/CARRYB[55][5] , \mult_22/CARRYB[55][6] ,
         \mult_22/CARRYB[55][7] , \mult_22/CARRYB[55][8] ,
         \mult_22/CARRYB[55][9] , \mult_22/CARRYB[55][10] ,
         \mult_22/CARRYB[55][11] , \mult_22/CARRYB[55][12] ,
         \mult_22/CARRYB[55][13] , \mult_22/CARRYB[55][14] ,
         \mult_22/CARRYB[55][15] , \mult_22/CARRYB[55][16] ,
         \mult_22/CARRYB[55][17] , \mult_22/CARRYB[55][18] ,
         \mult_22/CARRYB[55][19] , \mult_22/CARRYB[55][20] ,
         \mult_22/CARRYB[55][21] , \mult_22/CARRYB[55][22] ,
         \mult_22/CARRYB[55][23] , \mult_22/CARRYB[55][24] ,
         \mult_22/CARRYB[55][25] , \mult_22/CARRYB[55][26] ,
         \mult_22/CARRYB[55][27] , \mult_22/CARRYB[55][28] ,
         \mult_22/CARRYB[55][29] , \mult_22/CARRYB[55][30] ,
         \mult_22/CARRYB[55][31] , \mult_22/CARRYB[55][32] ,
         \mult_22/CARRYB[55][33] , \mult_22/CARRYB[55][34] ,
         \mult_22/CARRYB[55][35] , \mult_22/CARRYB[55][36] ,
         \mult_22/CARRYB[55][37] , \mult_22/CARRYB[55][38] ,
         \mult_22/CARRYB[55][39] , \mult_22/CARRYB[55][40] ,
         \mult_22/CARRYB[55][41] , \mult_22/CARRYB[55][42] ,
         \mult_22/CARRYB[55][43] , \mult_22/CARRYB[55][44] ,
         \mult_22/CARRYB[55][45] , \mult_22/CARRYB[55][46] ,
         \mult_22/CARRYB[55][47] , \mult_22/CARRYB[55][48] ,
         \mult_22/CARRYB[55][49] , \mult_22/CARRYB[55][50] ,
         \mult_22/CARRYB[55][51] , \mult_22/CARRYB[55][52] ,
         \mult_22/CARRYB[55][53] , \mult_22/CARRYB[55][54] ,
         \mult_22/CARRYB[55][55] , \mult_22/CARRYB[55][56] ,
         \mult_22/CARRYB[55][57] , \mult_22/CARRYB[55][58] ,
         \mult_22/CARRYB[55][59] , \mult_22/CARRYB[55][60] ,
         \mult_22/CARRYB[55][61] , \mult_22/CARRYB[55][62] ,
         \mult_22/SUMB[40][1] , \mult_22/SUMB[40][2] , \mult_22/SUMB[40][3] ,
         \mult_22/SUMB[40][4] , \mult_22/SUMB[40][5] , \mult_22/SUMB[40][6] ,
         \mult_22/SUMB[40][7] , \mult_22/SUMB[40][8] , \mult_22/SUMB[40][9] ,
         \mult_22/SUMB[40][10] , \mult_22/SUMB[40][11] ,
         \mult_22/SUMB[40][12] , \mult_22/SUMB[40][13] ,
         \mult_22/SUMB[40][14] , \mult_22/SUMB[40][15] ,
         \mult_22/SUMB[40][16] , \mult_22/SUMB[40][17] ,
         \mult_22/SUMB[40][18] , \mult_22/SUMB[40][19] ,
         \mult_22/SUMB[40][20] , \mult_22/SUMB[40][21] ,
         \mult_22/SUMB[40][22] , \mult_22/SUMB[40][23] ,
         \mult_22/SUMB[40][24] , \mult_22/SUMB[40][25] ,
         \mult_22/SUMB[40][26] , \mult_22/SUMB[40][27] ,
         \mult_22/SUMB[40][28] , \mult_22/SUMB[40][29] ,
         \mult_22/SUMB[40][30] , \mult_22/SUMB[40][31] ,
         \mult_22/SUMB[40][32] , \mult_22/SUMB[40][33] ,
         \mult_22/SUMB[40][34] , \mult_22/SUMB[40][35] ,
         \mult_22/SUMB[40][36] , \mult_22/SUMB[40][37] ,
         \mult_22/SUMB[40][38] , \mult_22/SUMB[40][39] ,
         \mult_22/SUMB[40][40] , \mult_22/SUMB[40][41] ,
         \mult_22/SUMB[40][42] , \mult_22/SUMB[40][43] ,
         \mult_22/SUMB[40][44] , \mult_22/SUMB[40][45] ,
         \mult_22/SUMB[40][46] , \mult_22/SUMB[40][47] ,
         \mult_22/SUMB[40][48] , \mult_22/SUMB[40][49] ,
         \mult_22/SUMB[40][50] , \mult_22/SUMB[40][51] ,
         \mult_22/SUMB[40][52] , \mult_22/SUMB[40][53] ,
         \mult_22/SUMB[40][54] , \mult_22/SUMB[40][55] ,
         \mult_22/SUMB[40][56] , \mult_22/SUMB[40][57] ,
         \mult_22/SUMB[40][58] , \mult_22/SUMB[40][59] ,
         \mult_22/SUMB[40][60] , \mult_22/SUMB[40][61] ,
         \mult_22/SUMB[40][62] , \mult_22/SUMB[41][1] , \mult_22/SUMB[41][2] ,
         \mult_22/SUMB[41][3] , \mult_22/SUMB[41][4] , \mult_22/SUMB[41][5] ,
         \mult_22/SUMB[41][6] , \mult_22/SUMB[41][7] , \mult_22/SUMB[41][8] ,
         \mult_22/SUMB[41][9] , \mult_22/SUMB[41][10] , \mult_22/SUMB[41][11] ,
         \mult_22/SUMB[41][12] , \mult_22/SUMB[41][13] ,
         \mult_22/SUMB[41][14] , \mult_22/SUMB[41][15] ,
         \mult_22/SUMB[41][16] , \mult_22/SUMB[41][17] ,
         \mult_22/SUMB[41][18] , \mult_22/SUMB[41][19] ,
         \mult_22/SUMB[41][20] , \mult_22/SUMB[41][21] ,
         \mult_22/SUMB[41][22] , \mult_22/SUMB[41][23] ,
         \mult_22/SUMB[41][24] , \mult_22/SUMB[41][25] ,
         \mult_22/SUMB[41][26] , \mult_22/SUMB[41][27] ,
         \mult_22/SUMB[41][28] , \mult_22/SUMB[41][29] ,
         \mult_22/SUMB[41][30] , \mult_22/SUMB[41][31] ,
         \mult_22/SUMB[41][32] , \mult_22/SUMB[41][33] ,
         \mult_22/SUMB[41][34] , \mult_22/SUMB[41][35] ,
         \mult_22/SUMB[41][36] , \mult_22/SUMB[41][37] ,
         \mult_22/SUMB[41][38] , \mult_22/SUMB[41][39] ,
         \mult_22/SUMB[41][40] , \mult_22/SUMB[41][41] ,
         \mult_22/SUMB[41][42] , \mult_22/SUMB[41][43] ,
         \mult_22/SUMB[41][44] , \mult_22/SUMB[41][45] ,
         \mult_22/SUMB[41][46] , \mult_22/SUMB[41][47] ,
         \mult_22/SUMB[41][48] , \mult_22/SUMB[41][49] ,
         \mult_22/SUMB[41][50] , \mult_22/SUMB[41][51] ,
         \mult_22/SUMB[41][52] , \mult_22/SUMB[41][53] ,
         \mult_22/SUMB[41][54] , \mult_22/SUMB[41][55] ,
         \mult_22/SUMB[41][56] , \mult_22/SUMB[41][57] ,
         \mult_22/SUMB[41][58] , \mult_22/SUMB[41][59] ,
         \mult_22/SUMB[41][60] , \mult_22/SUMB[41][61] ,
         \mult_22/SUMB[41][62] , \mult_22/SUMB[42][1] , \mult_22/SUMB[42][2] ,
         \mult_22/SUMB[42][3] , \mult_22/SUMB[42][4] , \mult_22/SUMB[42][5] ,
         \mult_22/SUMB[42][6] , \mult_22/SUMB[42][7] , \mult_22/SUMB[42][8] ,
         \mult_22/SUMB[42][9] , \mult_22/SUMB[42][10] , \mult_22/SUMB[42][11] ,
         \mult_22/SUMB[42][12] , \mult_22/SUMB[42][13] ,
         \mult_22/SUMB[42][14] , \mult_22/SUMB[42][15] ,
         \mult_22/SUMB[42][16] , \mult_22/SUMB[42][17] ,
         \mult_22/SUMB[42][18] , \mult_22/SUMB[42][19] ,
         \mult_22/SUMB[42][20] , \mult_22/SUMB[42][21] ,
         \mult_22/SUMB[42][22] , \mult_22/SUMB[42][23] ,
         \mult_22/SUMB[42][24] , \mult_22/SUMB[42][25] ,
         \mult_22/SUMB[42][26] , \mult_22/SUMB[42][27] ,
         \mult_22/SUMB[42][28] , \mult_22/SUMB[42][29] ,
         \mult_22/SUMB[42][30] , \mult_22/SUMB[42][31] ,
         \mult_22/SUMB[42][32] , \mult_22/SUMB[42][33] ,
         \mult_22/SUMB[42][34] , \mult_22/SUMB[42][35] ,
         \mult_22/SUMB[42][36] , \mult_22/SUMB[42][37] ,
         \mult_22/SUMB[42][38] , \mult_22/SUMB[42][39] ,
         \mult_22/SUMB[42][40] , \mult_22/SUMB[42][41] ,
         \mult_22/SUMB[42][42] , \mult_22/SUMB[42][43] ,
         \mult_22/SUMB[42][44] , \mult_22/SUMB[42][45] ,
         \mult_22/SUMB[42][46] , \mult_22/SUMB[42][47] ,
         \mult_22/SUMB[42][48] , \mult_22/SUMB[42][49] ,
         \mult_22/SUMB[42][50] , \mult_22/SUMB[42][51] ,
         \mult_22/SUMB[42][52] , \mult_22/SUMB[42][53] ,
         \mult_22/SUMB[42][54] , \mult_22/SUMB[42][55] ,
         \mult_22/SUMB[42][56] , \mult_22/SUMB[42][57] ,
         \mult_22/SUMB[42][58] , \mult_22/SUMB[42][59] ,
         \mult_22/SUMB[42][60] , \mult_22/SUMB[42][61] ,
         \mult_22/SUMB[42][62] , \mult_22/SUMB[43][1] , \mult_22/SUMB[43][2] ,
         \mult_22/SUMB[43][3] , \mult_22/SUMB[43][4] , \mult_22/SUMB[43][5] ,
         \mult_22/SUMB[43][6] , \mult_22/SUMB[43][7] , \mult_22/SUMB[43][8] ,
         \mult_22/SUMB[43][9] , \mult_22/SUMB[43][10] , \mult_22/SUMB[43][11] ,
         \mult_22/SUMB[43][12] , \mult_22/SUMB[43][13] ,
         \mult_22/SUMB[43][14] , \mult_22/SUMB[43][15] ,
         \mult_22/SUMB[43][16] , \mult_22/SUMB[43][17] ,
         \mult_22/SUMB[43][18] , \mult_22/SUMB[43][19] ,
         \mult_22/SUMB[43][20] , \mult_22/SUMB[43][21] ,
         \mult_22/SUMB[43][22] , \mult_22/SUMB[43][23] ,
         \mult_22/SUMB[43][24] , \mult_22/SUMB[43][25] ,
         \mult_22/SUMB[43][26] , \mult_22/SUMB[43][27] ,
         \mult_22/SUMB[43][28] , \mult_22/SUMB[43][29] ,
         \mult_22/SUMB[43][30] , \mult_22/SUMB[43][31] ,
         \mult_22/SUMB[43][32] , \mult_22/SUMB[43][33] ,
         \mult_22/SUMB[43][34] , \mult_22/SUMB[43][35] ,
         \mult_22/SUMB[43][36] , \mult_22/SUMB[43][37] ,
         \mult_22/SUMB[43][38] , \mult_22/SUMB[43][39] ,
         \mult_22/SUMB[43][40] , \mult_22/SUMB[43][41] ,
         \mult_22/SUMB[43][42] , \mult_22/SUMB[43][43] ,
         \mult_22/SUMB[43][44] , \mult_22/SUMB[43][45] ,
         \mult_22/SUMB[43][46] , \mult_22/SUMB[43][47] ,
         \mult_22/SUMB[43][48] , \mult_22/SUMB[43][49] ,
         \mult_22/SUMB[43][50] , \mult_22/SUMB[43][51] ,
         \mult_22/SUMB[43][52] , \mult_22/SUMB[43][53] ,
         \mult_22/SUMB[43][54] , \mult_22/SUMB[43][55] ,
         \mult_22/SUMB[43][56] , \mult_22/SUMB[43][57] ,
         \mult_22/SUMB[43][58] , \mult_22/SUMB[43][59] ,
         \mult_22/SUMB[43][60] , \mult_22/SUMB[43][61] ,
         \mult_22/SUMB[43][62] , \mult_22/SUMB[44][1] , \mult_22/SUMB[44][2] ,
         \mult_22/SUMB[44][3] , \mult_22/SUMB[44][4] , \mult_22/SUMB[44][5] ,
         \mult_22/SUMB[44][6] , \mult_22/SUMB[44][7] , \mult_22/SUMB[44][8] ,
         \mult_22/SUMB[44][9] , \mult_22/SUMB[44][10] , \mult_22/SUMB[44][11] ,
         \mult_22/SUMB[44][12] , \mult_22/SUMB[44][13] ,
         \mult_22/SUMB[44][14] , \mult_22/SUMB[44][15] ,
         \mult_22/SUMB[44][16] , \mult_22/SUMB[44][17] ,
         \mult_22/SUMB[44][18] , \mult_22/SUMB[44][19] ,
         \mult_22/SUMB[44][20] , \mult_22/SUMB[44][21] ,
         \mult_22/SUMB[44][22] , \mult_22/SUMB[44][23] ,
         \mult_22/SUMB[44][24] , \mult_22/SUMB[44][25] ,
         \mult_22/SUMB[44][26] , \mult_22/SUMB[44][27] ,
         \mult_22/SUMB[44][28] , \mult_22/SUMB[44][29] ,
         \mult_22/SUMB[44][30] , \mult_22/SUMB[44][31] ,
         \mult_22/SUMB[44][32] , \mult_22/SUMB[44][33] ,
         \mult_22/SUMB[44][34] , \mult_22/SUMB[44][35] ,
         \mult_22/SUMB[44][36] , \mult_22/SUMB[44][37] ,
         \mult_22/SUMB[44][38] , \mult_22/SUMB[44][39] ,
         \mult_22/SUMB[44][40] , \mult_22/SUMB[44][41] ,
         \mult_22/SUMB[44][42] , \mult_22/SUMB[44][43] ,
         \mult_22/SUMB[44][44] , \mult_22/SUMB[44][45] ,
         \mult_22/SUMB[44][46] , \mult_22/SUMB[44][47] ,
         \mult_22/SUMB[44][48] , \mult_22/SUMB[44][49] ,
         \mult_22/SUMB[44][50] , \mult_22/SUMB[44][51] ,
         \mult_22/SUMB[44][52] , \mult_22/SUMB[44][53] ,
         \mult_22/SUMB[44][54] , \mult_22/SUMB[44][55] ,
         \mult_22/SUMB[44][56] , \mult_22/SUMB[44][57] ,
         \mult_22/SUMB[44][58] , \mult_22/SUMB[44][59] ,
         \mult_22/SUMB[44][60] , \mult_22/SUMB[44][61] ,
         \mult_22/SUMB[44][62] , \mult_22/SUMB[45][1] , \mult_22/SUMB[45][2] ,
         \mult_22/SUMB[45][3] , \mult_22/SUMB[45][4] , \mult_22/SUMB[45][5] ,
         \mult_22/SUMB[45][6] , \mult_22/SUMB[45][7] , \mult_22/SUMB[45][8] ,
         \mult_22/SUMB[45][9] , \mult_22/SUMB[45][10] , \mult_22/SUMB[45][11] ,
         \mult_22/SUMB[45][12] , \mult_22/SUMB[45][13] ,
         \mult_22/SUMB[45][14] , \mult_22/SUMB[45][15] ,
         \mult_22/SUMB[45][16] , \mult_22/SUMB[45][17] ,
         \mult_22/SUMB[45][18] , \mult_22/SUMB[45][19] ,
         \mult_22/SUMB[45][20] , \mult_22/SUMB[45][21] ,
         \mult_22/SUMB[45][22] , \mult_22/SUMB[45][23] ,
         \mult_22/SUMB[45][24] , \mult_22/SUMB[45][25] ,
         \mult_22/SUMB[45][26] , \mult_22/SUMB[45][27] ,
         \mult_22/SUMB[45][28] , \mult_22/SUMB[45][29] ,
         \mult_22/SUMB[45][30] , \mult_22/SUMB[45][31] ,
         \mult_22/SUMB[45][32] , \mult_22/SUMB[45][33] ,
         \mult_22/SUMB[45][34] , \mult_22/SUMB[45][35] ,
         \mult_22/SUMB[45][36] , \mult_22/SUMB[45][37] ,
         \mult_22/SUMB[45][38] , \mult_22/SUMB[45][39] ,
         \mult_22/SUMB[45][40] , \mult_22/SUMB[45][41] ,
         \mult_22/SUMB[45][42] , \mult_22/SUMB[45][43] ,
         \mult_22/SUMB[45][44] , \mult_22/SUMB[45][45] ,
         \mult_22/SUMB[45][46] , \mult_22/SUMB[45][47] ,
         \mult_22/SUMB[45][48] , \mult_22/SUMB[45][49] ,
         \mult_22/SUMB[45][50] , \mult_22/SUMB[45][51] ,
         \mult_22/SUMB[45][52] , \mult_22/SUMB[45][53] ,
         \mult_22/SUMB[45][54] , \mult_22/SUMB[45][55] ,
         \mult_22/SUMB[45][56] , \mult_22/SUMB[45][57] ,
         \mult_22/SUMB[45][58] , \mult_22/SUMB[45][59] ,
         \mult_22/SUMB[45][60] , \mult_22/SUMB[45][61] ,
         \mult_22/SUMB[45][62] , \mult_22/SUMB[46][1] , \mult_22/SUMB[46][2] ,
         \mult_22/SUMB[46][3] , \mult_22/SUMB[46][4] , \mult_22/SUMB[46][5] ,
         \mult_22/SUMB[46][6] , \mult_22/SUMB[46][7] , \mult_22/SUMB[46][8] ,
         \mult_22/SUMB[46][9] , \mult_22/SUMB[46][10] , \mult_22/SUMB[46][11] ,
         \mult_22/SUMB[46][12] , \mult_22/SUMB[46][13] ,
         \mult_22/SUMB[46][14] , \mult_22/SUMB[46][15] ,
         \mult_22/SUMB[46][16] , \mult_22/SUMB[46][17] ,
         \mult_22/SUMB[46][18] , \mult_22/SUMB[46][19] ,
         \mult_22/SUMB[46][20] , \mult_22/SUMB[46][21] ,
         \mult_22/SUMB[46][22] , \mult_22/SUMB[46][23] ,
         \mult_22/SUMB[46][24] , \mult_22/SUMB[46][25] ,
         \mult_22/SUMB[46][26] , \mult_22/SUMB[46][27] ,
         \mult_22/SUMB[46][28] , \mult_22/SUMB[46][29] ,
         \mult_22/SUMB[46][30] , \mult_22/SUMB[46][31] ,
         \mult_22/SUMB[46][32] , \mult_22/SUMB[46][33] ,
         \mult_22/SUMB[46][34] , \mult_22/SUMB[46][35] ,
         \mult_22/SUMB[46][36] , \mult_22/SUMB[46][37] ,
         \mult_22/SUMB[46][38] , \mult_22/SUMB[46][39] ,
         \mult_22/SUMB[46][40] , \mult_22/SUMB[46][41] ,
         \mult_22/SUMB[46][42] , \mult_22/SUMB[46][43] ,
         \mult_22/SUMB[46][44] , \mult_22/SUMB[46][45] ,
         \mult_22/SUMB[46][46] , \mult_22/SUMB[46][47] ,
         \mult_22/SUMB[46][48] , \mult_22/SUMB[46][49] ,
         \mult_22/SUMB[46][50] , \mult_22/SUMB[46][51] ,
         \mult_22/SUMB[46][52] , \mult_22/SUMB[46][53] ,
         \mult_22/SUMB[46][54] , \mult_22/SUMB[46][55] ,
         \mult_22/SUMB[46][56] , \mult_22/SUMB[46][57] ,
         \mult_22/SUMB[46][58] , \mult_22/SUMB[46][59] ,
         \mult_22/SUMB[46][60] , \mult_22/SUMB[46][61] ,
         \mult_22/SUMB[46][62] , \mult_22/SUMB[47][1] , \mult_22/SUMB[47][2] ,
         \mult_22/SUMB[47][3] , \mult_22/SUMB[47][4] , \mult_22/SUMB[47][5] ,
         \mult_22/SUMB[47][6] , \mult_22/SUMB[47][7] , \mult_22/SUMB[47][8] ,
         \mult_22/SUMB[47][9] , \mult_22/SUMB[47][10] , \mult_22/SUMB[47][11] ,
         \mult_22/SUMB[47][12] , \mult_22/SUMB[47][13] ,
         \mult_22/SUMB[47][14] , \mult_22/SUMB[47][15] ,
         \mult_22/SUMB[47][16] , \mult_22/SUMB[47][17] ,
         \mult_22/SUMB[47][18] , \mult_22/SUMB[47][19] ,
         \mult_22/SUMB[47][20] , \mult_22/SUMB[47][21] ,
         \mult_22/SUMB[47][22] , \mult_22/SUMB[47][23] ,
         \mult_22/SUMB[47][24] , \mult_22/SUMB[47][25] ,
         \mult_22/SUMB[47][26] , \mult_22/SUMB[47][27] ,
         \mult_22/SUMB[47][28] , \mult_22/SUMB[47][29] ,
         \mult_22/SUMB[47][30] , \mult_22/SUMB[47][31] ,
         \mult_22/SUMB[47][32] , \mult_22/SUMB[47][33] ,
         \mult_22/SUMB[47][34] , \mult_22/SUMB[47][35] ,
         \mult_22/SUMB[47][36] , \mult_22/SUMB[47][37] ,
         \mult_22/SUMB[47][38] , \mult_22/SUMB[47][39] ,
         \mult_22/SUMB[47][40] , \mult_22/SUMB[47][41] ,
         \mult_22/SUMB[47][42] , \mult_22/SUMB[47][43] ,
         \mult_22/SUMB[47][44] , \mult_22/SUMB[47][45] ,
         \mult_22/SUMB[47][46] , \mult_22/SUMB[47][47] ,
         \mult_22/SUMB[47][48] , \mult_22/SUMB[47][49] ,
         \mult_22/SUMB[47][50] , \mult_22/SUMB[47][51] ,
         \mult_22/SUMB[47][52] , \mult_22/SUMB[47][53] ,
         \mult_22/SUMB[47][54] , \mult_22/SUMB[47][55] ,
         \mult_22/SUMB[47][56] , \mult_22/SUMB[47][57] ,
         \mult_22/SUMB[47][58] , \mult_22/SUMB[47][59] ,
         \mult_22/SUMB[47][60] , \mult_22/SUMB[47][61] ,
         \mult_22/SUMB[47][62] , \mult_22/CARRYB[40][0] ,
         \mult_22/CARRYB[40][1] , \mult_22/CARRYB[40][2] ,
         \mult_22/CARRYB[40][3] , \mult_22/CARRYB[40][4] ,
         \mult_22/CARRYB[40][5] , \mult_22/CARRYB[40][6] ,
         \mult_22/CARRYB[40][7] , \mult_22/CARRYB[40][8] ,
         \mult_22/CARRYB[40][9] , \mult_22/CARRYB[40][10] ,
         \mult_22/CARRYB[40][11] , \mult_22/CARRYB[40][12] ,
         \mult_22/CARRYB[40][13] , \mult_22/CARRYB[40][14] ,
         \mult_22/CARRYB[40][15] , \mult_22/CARRYB[40][16] ,
         \mult_22/CARRYB[40][17] , \mult_22/CARRYB[40][18] ,
         \mult_22/CARRYB[40][19] , \mult_22/CARRYB[40][20] ,
         \mult_22/CARRYB[40][21] , \mult_22/CARRYB[40][22] ,
         \mult_22/CARRYB[40][23] , \mult_22/CARRYB[40][24] ,
         \mult_22/CARRYB[40][25] , \mult_22/CARRYB[40][26] ,
         \mult_22/CARRYB[40][27] , \mult_22/CARRYB[40][28] ,
         \mult_22/CARRYB[40][29] , \mult_22/CARRYB[40][30] ,
         \mult_22/CARRYB[40][31] , \mult_22/CARRYB[40][32] ,
         \mult_22/CARRYB[40][33] , \mult_22/CARRYB[40][34] ,
         \mult_22/CARRYB[40][35] , \mult_22/CARRYB[40][36] ,
         \mult_22/CARRYB[40][37] , \mult_22/CARRYB[40][38] ,
         \mult_22/CARRYB[40][39] , \mult_22/CARRYB[40][40] ,
         \mult_22/CARRYB[40][41] , \mult_22/CARRYB[40][42] ,
         \mult_22/CARRYB[40][43] , \mult_22/CARRYB[40][44] ,
         \mult_22/CARRYB[40][45] , \mult_22/CARRYB[40][46] ,
         \mult_22/CARRYB[40][47] , \mult_22/CARRYB[40][48] ,
         \mult_22/CARRYB[40][49] , \mult_22/CARRYB[40][50] ,
         \mult_22/CARRYB[40][51] , \mult_22/CARRYB[40][52] ,
         \mult_22/CARRYB[40][53] , \mult_22/CARRYB[40][54] ,
         \mult_22/CARRYB[40][55] , \mult_22/CARRYB[40][56] ,
         \mult_22/CARRYB[40][57] , \mult_22/CARRYB[40][58] ,
         \mult_22/CARRYB[40][59] , \mult_22/CARRYB[40][60] ,
         \mult_22/CARRYB[40][61] , \mult_22/CARRYB[40][62] ,
         \mult_22/CARRYB[41][0] , \mult_22/CARRYB[41][1] ,
         \mult_22/CARRYB[41][2] , \mult_22/CARRYB[41][3] ,
         \mult_22/CARRYB[41][4] , \mult_22/CARRYB[41][5] ,
         \mult_22/CARRYB[41][6] , \mult_22/CARRYB[41][7] ,
         \mult_22/CARRYB[41][8] , \mult_22/CARRYB[41][9] ,
         \mult_22/CARRYB[41][10] , \mult_22/CARRYB[41][11] ,
         \mult_22/CARRYB[41][12] , \mult_22/CARRYB[41][13] ,
         \mult_22/CARRYB[41][14] , \mult_22/CARRYB[41][15] ,
         \mult_22/CARRYB[41][16] , \mult_22/CARRYB[41][17] ,
         \mult_22/CARRYB[41][18] , \mult_22/CARRYB[41][19] ,
         \mult_22/CARRYB[41][20] , \mult_22/CARRYB[41][21] ,
         \mult_22/CARRYB[41][22] , \mult_22/CARRYB[41][23] ,
         \mult_22/CARRYB[41][24] , \mult_22/CARRYB[41][25] ,
         \mult_22/CARRYB[41][26] , \mult_22/CARRYB[41][27] ,
         \mult_22/CARRYB[41][28] , \mult_22/CARRYB[41][29] ,
         \mult_22/CARRYB[41][30] , \mult_22/CARRYB[41][31] ,
         \mult_22/CARRYB[41][32] , \mult_22/CARRYB[41][33] ,
         \mult_22/CARRYB[41][34] , \mult_22/CARRYB[41][35] ,
         \mult_22/CARRYB[41][36] , \mult_22/CARRYB[41][37] ,
         \mult_22/CARRYB[41][38] , \mult_22/CARRYB[41][39] ,
         \mult_22/CARRYB[41][40] , \mult_22/CARRYB[41][41] ,
         \mult_22/CARRYB[41][42] , \mult_22/CARRYB[41][43] ,
         \mult_22/CARRYB[41][44] , \mult_22/CARRYB[41][45] ,
         \mult_22/CARRYB[41][46] , \mult_22/CARRYB[41][47] ,
         \mult_22/CARRYB[41][48] , \mult_22/CARRYB[41][49] ,
         \mult_22/CARRYB[41][50] , \mult_22/CARRYB[41][51] ,
         \mult_22/CARRYB[41][52] , \mult_22/CARRYB[41][53] ,
         \mult_22/CARRYB[41][54] , \mult_22/CARRYB[41][55] ,
         \mult_22/CARRYB[41][56] , \mult_22/CARRYB[41][57] ,
         \mult_22/CARRYB[41][58] , \mult_22/CARRYB[41][59] ,
         \mult_22/CARRYB[41][60] , \mult_22/CARRYB[41][61] ,
         \mult_22/CARRYB[41][62] , \mult_22/CARRYB[42][0] ,
         \mult_22/CARRYB[42][1] , \mult_22/CARRYB[42][2] ,
         \mult_22/CARRYB[42][3] , \mult_22/CARRYB[42][4] ,
         \mult_22/CARRYB[42][5] , \mult_22/CARRYB[42][6] ,
         \mult_22/CARRYB[42][7] , \mult_22/CARRYB[42][8] ,
         \mult_22/CARRYB[42][9] , \mult_22/CARRYB[42][10] ,
         \mult_22/CARRYB[42][11] , \mult_22/CARRYB[42][12] ,
         \mult_22/CARRYB[42][13] , \mult_22/CARRYB[42][14] ,
         \mult_22/CARRYB[42][15] , \mult_22/CARRYB[42][16] ,
         \mult_22/CARRYB[42][17] , \mult_22/CARRYB[42][18] ,
         \mult_22/CARRYB[42][19] , \mult_22/CARRYB[42][20] ,
         \mult_22/CARRYB[42][21] , \mult_22/CARRYB[42][22] ,
         \mult_22/CARRYB[42][23] , \mult_22/CARRYB[42][24] ,
         \mult_22/CARRYB[42][25] , \mult_22/CARRYB[42][26] ,
         \mult_22/CARRYB[42][27] , \mult_22/CARRYB[42][28] ,
         \mult_22/CARRYB[42][29] , \mult_22/CARRYB[42][30] ,
         \mult_22/CARRYB[42][31] , \mult_22/CARRYB[42][32] ,
         \mult_22/CARRYB[42][33] , \mult_22/CARRYB[42][34] ,
         \mult_22/CARRYB[42][35] , \mult_22/CARRYB[42][36] ,
         \mult_22/CARRYB[42][37] , \mult_22/CARRYB[42][38] ,
         \mult_22/CARRYB[42][39] , \mult_22/CARRYB[42][40] ,
         \mult_22/CARRYB[42][41] , \mult_22/CARRYB[42][42] ,
         \mult_22/CARRYB[42][43] , \mult_22/CARRYB[42][44] ,
         \mult_22/CARRYB[42][45] , \mult_22/CARRYB[42][46] ,
         \mult_22/CARRYB[42][47] , \mult_22/CARRYB[42][48] ,
         \mult_22/CARRYB[42][49] , \mult_22/CARRYB[42][50] ,
         \mult_22/CARRYB[42][51] , \mult_22/CARRYB[42][52] ,
         \mult_22/CARRYB[42][53] , \mult_22/CARRYB[42][54] ,
         \mult_22/CARRYB[42][55] , \mult_22/CARRYB[42][56] ,
         \mult_22/CARRYB[42][57] , \mult_22/CARRYB[42][58] ,
         \mult_22/CARRYB[42][59] , \mult_22/CARRYB[42][60] ,
         \mult_22/CARRYB[42][61] , \mult_22/CARRYB[42][62] ,
         \mult_22/CARRYB[43][0] , \mult_22/CARRYB[43][1] ,
         \mult_22/CARRYB[43][2] , \mult_22/CARRYB[43][3] ,
         \mult_22/CARRYB[43][4] , \mult_22/CARRYB[43][5] ,
         \mult_22/CARRYB[43][6] , \mult_22/CARRYB[43][7] ,
         \mult_22/CARRYB[43][8] , \mult_22/CARRYB[43][9] ,
         \mult_22/CARRYB[43][10] , \mult_22/CARRYB[43][11] ,
         \mult_22/CARRYB[43][12] , \mult_22/CARRYB[43][13] ,
         \mult_22/CARRYB[43][14] , \mult_22/CARRYB[43][15] ,
         \mult_22/CARRYB[43][16] , \mult_22/CARRYB[43][17] ,
         \mult_22/CARRYB[43][18] , \mult_22/CARRYB[43][19] ,
         \mult_22/CARRYB[43][20] , \mult_22/CARRYB[43][21] ,
         \mult_22/CARRYB[43][22] , \mult_22/CARRYB[43][23] ,
         \mult_22/CARRYB[43][24] , \mult_22/CARRYB[43][25] ,
         \mult_22/CARRYB[43][26] , \mult_22/CARRYB[43][27] ,
         \mult_22/CARRYB[43][28] , \mult_22/CARRYB[43][29] ,
         \mult_22/CARRYB[43][30] , \mult_22/CARRYB[43][31] ,
         \mult_22/CARRYB[43][32] , \mult_22/CARRYB[43][33] ,
         \mult_22/CARRYB[43][34] , \mult_22/CARRYB[43][35] ,
         \mult_22/CARRYB[43][36] , \mult_22/CARRYB[43][37] ,
         \mult_22/CARRYB[43][38] , \mult_22/CARRYB[43][39] ,
         \mult_22/CARRYB[43][40] , \mult_22/CARRYB[43][41] ,
         \mult_22/CARRYB[43][42] , \mult_22/CARRYB[43][43] ,
         \mult_22/CARRYB[43][44] , \mult_22/CARRYB[43][45] ,
         \mult_22/CARRYB[43][46] , \mult_22/CARRYB[43][47] ,
         \mult_22/CARRYB[43][48] , \mult_22/CARRYB[43][49] ,
         \mult_22/CARRYB[43][50] , \mult_22/CARRYB[43][51] ,
         \mult_22/CARRYB[43][52] , \mult_22/CARRYB[43][53] ,
         \mult_22/CARRYB[43][54] , \mult_22/CARRYB[43][55] ,
         \mult_22/CARRYB[43][56] , \mult_22/CARRYB[43][57] ,
         \mult_22/CARRYB[43][58] , \mult_22/CARRYB[43][59] ,
         \mult_22/CARRYB[43][60] , \mult_22/CARRYB[43][61] ,
         \mult_22/CARRYB[43][62] , \mult_22/CARRYB[44][0] ,
         \mult_22/CARRYB[44][1] , \mult_22/CARRYB[44][2] ,
         \mult_22/CARRYB[44][3] , \mult_22/CARRYB[44][4] ,
         \mult_22/CARRYB[44][5] , \mult_22/CARRYB[44][6] ,
         \mult_22/CARRYB[44][7] , \mult_22/CARRYB[44][8] ,
         \mult_22/CARRYB[44][9] , \mult_22/CARRYB[44][10] ,
         \mult_22/CARRYB[44][11] , \mult_22/CARRYB[44][12] ,
         \mult_22/CARRYB[44][13] , \mult_22/CARRYB[44][14] ,
         \mult_22/CARRYB[44][15] , \mult_22/CARRYB[44][16] ,
         \mult_22/CARRYB[44][17] , \mult_22/CARRYB[44][18] ,
         \mult_22/CARRYB[44][19] , \mult_22/CARRYB[44][20] ,
         \mult_22/CARRYB[44][21] , \mult_22/CARRYB[44][22] ,
         \mult_22/CARRYB[44][23] , \mult_22/CARRYB[44][24] ,
         \mult_22/CARRYB[44][25] , \mult_22/CARRYB[44][26] ,
         \mult_22/CARRYB[44][27] , \mult_22/CARRYB[44][28] ,
         \mult_22/CARRYB[44][29] , \mult_22/CARRYB[44][30] ,
         \mult_22/CARRYB[44][31] , \mult_22/CARRYB[44][32] ,
         \mult_22/CARRYB[44][33] , \mult_22/CARRYB[44][34] ,
         \mult_22/CARRYB[44][35] , \mult_22/CARRYB[44][36] ,
         \mult_22/CARRYB[44][37] , \mult_22/CARRYB[44][38] ,
         \mult_22/CARRYB[44][39] , \mult_22/CARRYB[44][40] ,
         \mult_22/CARRYB[44][41] , \mult_22/CARRYB[44][42] ,
         \mult_22/CARRYB[44][43] , \mult_22/CARRYB[44][44] ,
         \mult_22/CARRYB[44][45] , \mult_22/CARRYB[44][46] ,
         \mult_22/CARRYB[44][47] , \mult_22/CARRYB[44][48] ,
         \mult_22/CARRYB[44][49] , \mult_22/CARRYB[44][50] ,
         \mult_22/CARRYB[44][51] , \mult_22/CARRYB[44][52] ,
         \mult_22/CARRYB[44][53] , \mult_22/CARRYB[44][54] ,
         \mult_22/CARRYB[44][55] , \mult_22/CARRYB[44][56] ,
         \mult_22/CARRYB[44][57] , \mult_22/CARRYB[44][58] ,
         \mult_22/CARRYB[44][59] , \mult_22/CARRYB[44][60] ,
         \mult_22/CARRYB[44][61] , \mult_22/CARRYB[44][62] ,
         \mult_22/CARRYB[45][0] , \mult_22/CARRYB[45][1] ,
         \mult_22/CARRYB[45][2] , \mult_22/CARRYB[45][3] ,
         \mult_22/CARRYB[45][4] , \mult_22/CARRYB[45][5] ,
         \mult_22/CARRYB[45][6] , \mult_22/CARRYB[45][7] ,
         \mult_22/CARRYB[45][8] , \mult_22/CARRYB[45][9] ,
         \mult_22/CARRYB[45][10] , \mult_22/CARRYB[45][11] ,
         \mult_22/CARRYB[45][12] , \mult_22/CARRYB[45][13] ,
         \mult_22/CARRYB[45][14] , \mult_22/CARRYB[45][15] ,
         \mult_22/CARRYB[45][16] , \mult_22/CARRYB[45][17] ,
         \mult_22/CARRYB[45][18] , \mult_22/CARRYB[45][19] ,
         \mult_22/CARRYB[45][20] , \mult_22/CARRYB[45][21] ,
         \mult_22/CARRYB[45][22] , \mult_22/CARRYB[45][23] ,
         \mult_22/CARRYB[45][24] , \mult_22/CARRYB[45][25] ,
         \mult_22/CARRYB[45][26] , \mult_22/CARRYB[45][27] ,
         \mult_22/CARRYB[45][28] , \mult_22/CARRYB[45][29] ,
         \mult_22/CARRYB[45][30] , \mult_22/CARRYB[45][31] ,
         \mult_22/CARRYB[45][32] , \mult_22/CARRYB[45][33] ,
         \mult_22/CARRYB[45][34] , \mult_22/CARRYB[45][35] ,
         \mult_22/CARRYB[45][36] , \mult_22/CARRYB[45][37] ,
         \mult_22/CARRYB[45][38] , \mult_22/CARRYB[45][39] ,
         \mult_22/CARRYB[45][40] , \mult_22/CARRYB[45][41] ,
         \mult_22/CARRYB[45][42] , \mult_22/CARRYB[45][43] ,
         \mult_22/CARRYB[45][44] , \mult_22/CARRYB[45][45] ,
         \mult_22/CARRYB[45][46] , \mult_22/CARRYB[45][47] ,
         \mult_22/CARRYB[45][48] , \mult_22/CARRYB[45][49] ,
         \mult_22/CARRYB[45][50] , \mult_22/CARRYB[45][51] ,
         \mult_22/CARRYB[45][52] , \mult_22/CARRYB[45][53] ,
         \mult_22/CARRYB[45][54] , \mult_22/CARRYB[45][55] ,
         \mult_22/CARRYB[45][56] , \mult_22/CARRYB[45][57] ,
         \mult_22/CARRYB[45][58] , \mult_22/CARRYB[45][59] ,
         \mult_22/CARRYB[45][60] , \mult_22/CARRYB[45][61] ,
         \mult_22/CARRYB[45][62] , \mult_22/CARRYB[46][0] ,
         \mult_22/CARRYB[46][1] , \mult_22/CARRYB[46][2] ,
         \mult_22/CARRYB[46][3] , \mult_22/CARRYB[46][4] ,
         \mult_22/CARRYB[46][5] , \mult_22/CARRYB[46][6] ,
         \mult_22/CARRYB[46][7] , \mult_22/CARRYB[46][8] ,
         \mult_22/CARRYB[46][9] , \mult_22/CARRYB[46][10] ,
         \mult_22/CARRYB[46][11] , \mult_22/CARRYB[46][12] ,
         \mult_22/CARRYB[46][13] , \mult_22/CARRYB[46][14] ,
         \mult_22/CARRYB[46][15] , \mult_22/CARRYB[46][16] ,
         \mult_22/CARRYB[46][17] , \mult_22/CARRYB[46][18] ,
         \mult_22/CARRYB[46][19] , \mult_22/CARRYB[46][20] ,
         \mult_22/CARRYB[46][21] , \mult_22/CARRYB[46][22] ,
         \mult_22/CARRYB[46][23] , \mult_22/CARRYB[46][24] ,
         \mult_22/CARRYB[46][25] , \mult_22/CARRYB[46][26] ,
         \mult_22/CARRYB[46][27] , \mult_22/CARRYB[46][28] ,
         \mult_22/CARRYB[46][29] , \mult_22/CARRYB[46][30] ,
         \mult_22/CARRYB[46][31] , \mult_22/CARRYB[46][32] ,
         \mult_22/CARRYB[46][33] , \mult_22/CARRYB[46][34] ,
         \mult_22/CARRYB[46][35] , \mult_22/CARRYB[46][36] ,
         \mult_22/CARRYB[46][37] , \mult_22/CARRYB[46][38] ,
         \mult_22/CARRYB[46][39] , \mult_22/CARRYB[46][40] ,
         \mult_22/CARRYB[46][41] , \mult_22/CARRYB[46][42] ,
         \mult_22/CARRYB[46][43] , \mult_22/CARRYB[46][44] ,
         \mult_22/CARRYB[46][45] , \mult_22/CARRYB[46][46] ,
         \mult_22/CARRYB[46][47] , \mult_22/CARRYB[46][48] ,
         \mult_22/CARRYB[46][49] , \mult_22/CARRYB[46][50] ,
         \mult_22/CARRYB[46][51] , \mult_22/CARRYB[46][52] ,
         \mult_22/CARRYB[46][53] , \mult_22/CARRYB[46][54] ,
         \mult_22/CARRYB[46][55] , \mult_22/CARRYB[46][56] ,
         \mult_22/CARRYB[46][57] , \mult_22/CARRYB[46][58] ,
         \mult_22/CARRYB[46][59] , \mult_22/CARRYB[46][60] ,
         \mult_22/CARRYB[46][61] , \mult_22/CARRYB[46][62] ,
         \mult_22/CARRYB[47][0] , \mult_22/CARRYB[47][1] ,
         \mult_22/CARRYB[47][2] , \mult_22/CARRYB[47][3] ,
         \mult_22/CARRYB[47][4] , \mult_22/CARRYB[47][5] ,
         \mult_22/CARRYB[47][6] , \mult_22/CARRYB[47][7] ,
         \mult_22/CARRYB[47][8] , \mult_22/CARRYB[47][9] ,
         \mult_22/CARRYB[47][10] , \mult_22/CARRYB[47][11] ,
         \mult_22/CARRYB[47][12] , \mult_22/CARRYB[47][13] ,
         \mult_22/CARRYB[47][14] , \mult_22/CARRYB[47][15] ,
         \mult_22/CARRYB[47][16] , \mult_22/CARRYB[47][17] ,
         \mult_22/CARRYB[47][18] , \mult_22/CARRYB[47][19] ,
         \mult_22/CARRYB[47][20] , \mult_22/CARRYB[47][21] ,
         \mult_22/CARRYB[47][22] , \mult_22/CARRYB[47][23] ,
         \mult_22/CARRYB[47][24] , \mult_22/CARRYB[47][25] ,
         \mult_22/CARRYB[47][26] , \mult_22/CARRYB[47][27] ,
         \mult_22/CARRYB[47][28] , \mult_22/CARRYB[47][29] ,
         \mult_22/CARRYB[47][30] , \mult_22/CARRYB[47][31] ,
         \mult_22/CARRYB[47][32] , \mult_22/CARRYB[47][33] ,
         \mult_22/CARRYB[47][34] , \mult_22/CARRYB[47][35] ,
         \mult_22/CARRYB[47][36] , \mult_22/CARRYB[47][37] ,
         \mult_22/CARRYB[47][38] , \mult_22/CARRYB[47][39] ,
         \mult_22/CARRYB[47][40] , \mult_22/CARRYB[47][41] ,
         \mult_22/CARRYB[47][42] , \mult_22/CARRYB[47][43] ,
         \mult_22/CARRYB[47][44] , \mult_22/CARRYB[47][45] ,
         \mult_22/CARRYB[47][46] , \mult_22/CARRYB[47][47] ,
         \mult_22/CARRYB[47][48] , \mult_22/CARRYB[47][49] ,
         \mult_22/CARRYB[47][50] , \mult_22/CARRYB[47][51] ,
         \mult_22/CARRYB[47][52] , \mult_22/CARRYB[47][53] ,
         \mult_22/CARRYB[47][54] , \mult_22/CARRYB[47][55] ,
         \mult_22/CARRYB[47][56] , \mult_22/CARRYB[47][57] ,
         \mult_22/CARRYB[47][58] , \mult_22/CARRYB[47][59] ,
         \mult_22/CARRYB[47][60] , \mult_22/CARRYB[47][61] ,
         \mult_22/CARRYB[47][62] , \mult_22/SUMB[32][1] ,
         \mult_22/SUMB[32][2] , \mult_22/SUMB[32][3] , \mult_22/SUMB[32][4] ,
         \mult_22/SUMB[32][5] , \mult_22/SUMB[32][6] , \mult_22/SUMB[32][7] ,
         \mult_22/SUMB[32][8] , \mult_22/SUMB[32][9] , \mult_22/SUMB[32][10] ,
         \mult_22/SUMB[32][11] , \mult_22/SUMB[32][12] ,
         \mult_22/SUMB[32][13] , \mult_22/SUMB[32][14] ,
         \mult_22/SUMB[32][15] , \mult_22/SUMB[32][16] ,
         \mult_22/SUMB[32][17] , \mult_22/SUMB[32][18] ,
         \mult_22/SUMB[32][19] , \mult_22/SUMB[32][20] ,
         \mult_22/SUMB[32][21] , \mult_22/SUMB[32][22] ,
         \mult_22/SUMB[32][23] , \mult_22/SUMB[32][24] ,
         \mult_22/SUMB[32][25] , \mult_22/SUMB[32][26] ,
         \mult_22/SUMB[32][27] , \mult_22/SUMB[32][28] ,
         \mult_22/SUMB[32][29] , \mult_22/SUMB[32][30] ,
         \mult_22/SUMB[32][31] , \mult_22/SUMB[32][32] ,
         \mult_22/SUMB[32][33] , \mult_22/SUMB[32][34] ,
         \mult_22/SUMB[32][35] , \mult_22/SUMB[32][36] ,
         \mult_22/SUMB[32][37] , \mult_22/SUMB[32][38] ,
         \mult_22/SUMB[32][39] , \mult_22/SUMB[32][40] ,
         \mult_22/SUMB[32][41] , \mult_22/SUMB[32][42] ,
         \mult_22/SUMB[32][43] , \mult_22/SUMB[32][44] ,
         \mult_22/SUMB[32][45] , \mult_22/SUMB[32][46] ,
         \mult_22/SUMB[32][47] , \mult_22/SUMB[32][48] ,
         \mult_22/SUMB[32][49] , \mult_22/SUMB[32][50] ,
         \mult_22/SUMB[32][51] , \mult_22/SUMB[32][52] ,
         \mult_22/SUMB[32][53] , \mult_22/SUMB[32][54] ,
         \mult_22/SUMB[32][55] , \mult_22/SUMB[32][56] ,
         \mult_22/SUMB[32][57] , \mult_22/SUMB[32][58] ,
         \mult_22/SUMB[32][59] , \mult_22/SUMB[32][60] ,
         \mult_22/SUMB[32][61] , \mult_22/SUMB[32][62] , \mult_22/SUMB[33][1] ,
         \mult_22/SUMB[33][2] , \mult_22/SUMB[33][3] , \mult_22/SUMB[33][4] ,
         \mult_22/SUMB[33][5] , \mult_22/SUMB[33][6] , \mult_22/SUMB[33][7] ,
         \mult_22/SUMB[33][8] , \mult_22/SUMB[33][9] , \mult_22/SUMB[33][10] ,
         \mult_22/SUMB[33][11] , \mult_22/SUMB[33][12] ,
         \mult_22/SUMB[33][13] , \mult_22/SUMB[33][14] ,
         \mult_22/SUMB[33][15] , \mult_22/SUMB[33][16] ,
         \mult_22/SUMB[33][17] , \mult_22/SUMB[33][18] ,
         \mult_22/SUMB[33][19] , \mult_22/SUMB[33][20] ,
         \mult_22/SUMB[33][21] , \mult_22/SUMB[33][22] ,
         \mult_22/SUMB[33][23] , \mult_22/SUMB[33][24] ,
         \mult_22/SUMB[33][25] , \mult_22/SUMB[33][26] ,
         \mult_22/SUMB[33][27] , \mult_22/SUMB[33][28] ,
         \mult_22/SUMB[33][29] , \mult_22/SUMB[33][30] ,
         \mult_22/SUMB[33][31] , \mult_22/SUMB[33][32] ,
         \mult_22/SUMB[33][33] , \mult_22/SUMB[33][34] ,
         \mult_22/SUMB[33][35] , \mult_22/SUMB[33][36] ,
         \mult_22/SUMB[33][37] , \mult_22/SUMB[33][38] ,
         \mult_22/SUMB[33][39] , \mult_22/SUMB[33][40] ,
         \mult_22/SUMB[33][41] , \mult_22/SUMB[33][42] ,
         \mult_22/SUMB[33][43] , \mult_22/SUMB[33][44] ,
         \mult_22/SUMB[33][45] , \mult_22/SUMB[33][46] ,
         \mult_22/SUMB[33][47] , \mult_22/SUMB[33][48] ,
         \mult_22/SUMB[33][49] , \mult_22/SUMB[33][50] ,
         \mult_22/SUMB[33][51] , \mult_22/SUMB[33][52] ,
         \mult_22/SUMB[33][53] , \mult_22/SUMB[33][54] ,
         \mult_22/SUMB[33][55] , \mult_22/SUMB[33][56] ,
         \mult_22/SUMB[33][57] , \mult_22/SUMB[33][58] ,
         \mult_22/SUMB[33][59] , \mult_22/SUMB[33][60] ,
         \mult_22/SUMB[33][61] , \mult_22/SUMB[33][62] , \mult_22/SUMB[34][1] ,
         \mult_22/SUMB[34][2] , \mult_22/SUMB[34][3] , \mult_22/SUMB[34][4] ,
         \mult_22/SUMB[34][5] , \mult_22/SUMB[34][6] , \mult_22/SUMB[34][7] ,
         \mult_22/SUMB[34][8] , \mult_22/SUMB[34][9] , \mult_22/SUMB[34][10] ,
         \mult_22/SUMB[34][11] , \mult_22/SUMB[34][12] ,
         \mult_22/SUMB[34][13] , \mult_22/SUMB[34][14] ,
         \mult_22/SUMB[34][15] , \mult_22/SUMB[34][16] ,
         \mult_22/SUMB[34][17] , \mult_22/SUMB[34][18] ,
         \mult_22/SUMB[34][19] , \mult_22/SUMB[34][20] ,
         \mult_22/SUMB[34][21] , \mult_22/SUMB[34][22] ,
         \mult_22/SUMB[34][23] , \mult_22/SUMB[34][24] ,
         \mult_22/SUMB[34][25] , \mult_22/SUMB[34][26] ,
         \mult_22/SUMB[34][27] , \mult_22/SUMB[34][28] ,
         \mult_22/SUMB[34][29] , \mult_22/SUMB[34][30] ,
         \mult_22/SUMB[34][31] , \mult_22/SUMB[34][32] ,
         \mult_22/SUMB[34][33] , \mult_22/SUMB[34][34] ,
         \mult_22/SUMB[34][35] , \mult_22/SUMB[34][36] ,
         \mult_22/SUMB[34][37] , \mult_22/SUMB[34][38] ,
         \mult_22/SUMB[34][39] , \mult_22/SUMB[34][40] ,
         \mult_22/SUMB[34][41] , \mult_22/SUMB[34][42] ,
         \mult_22/SUMB[34][43] , \mult_22/SUMB[34][44] ,
         \mult_22/SUMB[34][45] , \mult_22/SUMB[34][46] ,
         \mult_22/SUMB[34][47] , \mult_22/SUMB[34][48] ,
         \mult_22/SUMB[34][49] , \mult_22/SUMB[34][50] ,
         \mult_22/SUMB[34][51] , \mult_22/SUMB[34][52] ,
         \mult_22/SUMB[34][53] , \mult_22/SUMB[34][54] ,
         \mult_22/SUMB[34][55] , \mult_22/SUMB[34][56] ,
         \mult_22/SUMB[34][57] , \mult_22/SUMB[34][58] ,
         \mult_22/SUMB[34][59] , \mult_22/SUMB[34][60] ,
         \mult_22/SUMB[34][61] , \mult_22/SUMB[34][62] , \mult_22/SUMB[35][1] ,
         \mult_22/SUMB[35][2] , \mult_22/SUMB[35][3] , \mult_22/SUMB[35][4] ,
         \mult_22/SUMB[35][5] , \mult_22/SUMB[35][6] , \mult_22/SUMB[35][7] ,
         \mult_22/SUMB[35][8] , \mult_22/SUMB[35][9] , \mult_22/SUMB[35][10] ,
         \mult_22/SUMB[35][11] , \mult_22/SUMB[35][12] ,
         \mult_22/SUMB[35][13] , \mult_22/SUMB[35][14] ,
         \mult_22/SUMB[35][15] , \mult_22/SUMB[35][16] ,
         \mult_22/SUMB[35][17] , \mult_22/SUMB[35][18] ,
         \mult_22/SUMB[35][19] , \mult_22/SUMB[35][20] ,
         \mult_22/SUMB[35][21] , \mult_22/SUMB[35][22] ,
         \mult_22/SUMB[35][23] , \mult_22/SUMB[35][24] ,
         \mult_22/SUMB[35][25] , \mult_22/SUMB[35][26] ,
         \mult_22/SUMB[35][27] , \mult_22/SUMB[35][28] ,
         \mult_22/SUMB[35][29] , \mult_22/SUMB[35][30] ,
         \mult_22/SUMB[35][31] , \mult_22/SUMB[35][32] ,
         \mult_22/SUMB[35][33] , \mult_22/SUMB[35][34] ,
         \mult_22/SUMB[35][35] , \mult_22/SUMB[35][36] ,
         \mult_22/SUMB[35][37] , \mult_22/SUMB[35][38] ,
         \mult_22/SUMB[35][39] , \mult_22/SUMB[35][40] ,
         \mult_22/SUMB[35][41] , \mult_22/SUMB[35][42] ,
         \mult_22/SUMB[35][43] , \mult_22/SUMB[35][44] ,
         \mult_22/SUMB[35][45] , \mult_22/SUMB[35][46] ,
         \mult_22/SUMB[35][47] , \mult_22/SUMB[35][48] ,
         \mult_22/SUMB[35][49] , \mult_22/SUMB[35][50] ,
         \mult_22/SUMB[35][51] , \mult_22/SUMB[35][52] ,
         \mult_22/SUMB[35][53] , \mult_22/SUMB[35][54] ,
         \mult_22/SUMB[35][55] , \mult_22/SUMB[35][56] ,
         \mult_22/SUMB[35][57] , \mult_22/SUMB[35][58] ,
         \mult_22/SUMB[35][59] , \mult_22/SUMB[35][60] ,
         \mult_22/SUMB[35][61] , \mult_22/SUMB[35][62] , \mult_22/SUMB[36][1] ,
         \mult_22/SUMB[36][2] , \mult_22/SUMB[36][3] , \mult_22/SUMB[36][4] ,
         \mult_22/SUMB[36][5] , \mult_22/SUMB[36][6] , \mult_22/SUMB[36][7] ,
         \mult_22/SUMB[36][8] , \mult_22/SUMB[36][9] , \mult_22/SUMB[36][10] ,
         \mult_22/SUMB[36][11] , \mult_22/SUMB[36][12] ,
         \mult_22/SUMB[36][13] , \mult_22/SUMB[36][14] ,
         \mult_22/SUMB[36][15] , \mult_22/SUMB[36][16] ,
         \mult_22/SUMB[36][17] , \mult_22/SUMB[36][18] ,
         \mult_22/SUMB[36][19] , \mult_22/SUMB[36][20] ,
         \mult_22/SUMB[36][21] , \mult_22/SUMB[36][22] ,
         \mult_22/SUMB[36][23] , \mult_22/SUMB[36][24] ,
         \mult_22/SUMB[36][25] , \mult_22/SUMB[36][26] ,
         \mult_22/SUMB[36][27] , \mult_22/SUMB[36][28] ,
         \mult_22/SUMB[36][29] , \mult_22/SUMB[36][30] ,
         \mult_22/SUMB[36][31] , \mult_22/SUMB[36][32] ,
         \mult_22/SUMB[36][33] , \mult_22/SUMB[36][34] ,
         \mult_22/SUMB[36][35] , \mult_22/SUMB[36][36] ,
         \mult_22/SUMB[36][37] , \mult_22/SUMB[36][38] ,
         \mult_22/SUMB[36][39] , \mult_22/SUMB[36][40] ,
         \mult_22/SUMB[36][41] , \mult_22/SUMB[36][42] ,
         \mult_22/SUMB[36][43] , \mult_22/SUMB[36][44] ,
         \mult_22/SUMB[36][45] , \mult_22/SUMB[36][46] ,
         \mult_22/SUMB[36][47] , \mult_22/SUMB[36][48] ,
         \mult_22/SUMB[36][49] , \mult_22/SUMB[36][50] ,
         \mult_22/SUMB[36][51] , \mult_22/SUMB[36][52] ,
         \mult_22/SUMB[36][53] , \mult_22/SUMB[36][54] ,
         \mult_22/SUMB[36][55] , \mult_22/SUMB[36][56] ,
         \mult_22/SUMB[36][57] , \mult_22/SUMB[36][58] ,
         \mult_22/SUMB[36][59] , \mult_22/SUMB[36][60] ,
         \mult_22/SUMB[36][61] , \mult_22/SUMB[36][62] , \mult_22/SUMB[37][1] ,
         \mult_22/SUMB[37][2] , \mult_22/SUMB[37][3] , \mult_22/SUMB[37][4] ,
         \mult_22/SUMB[37][5] , \mult_22/SUMB[37][6] , \mult_22/SUMB[37][7] ,
         \mult_22/SUMB[37][8] , \mult_22/SUMB[37][9] , \mult_22/SUMB[37][10] ,
         \mult_22/SUMB[37][11] , \mult_22/SUMB[37][12] ,
         \mult_22/SUMB[37][13] , \mult_22/SUMB[37][14] ,
         \mult_22/SUMB[37][15] , \mult_22/SUMB[37][16] ,
         \mult_22/SUMB[37][17] , \mult_22/SUMB[37][18] ,
         \mult_22/SUMB[37][19] , \mult_22/SUMB[37][20] ,
         \mult_22/SUMB[37][21] , \mult_22/SUMB[37][22] ,
         \mult_22/SUMB[37][23] , \mult_22/SUMB[37][24] ,
         \mult_22/SUMB[37][25] , \mult_22/SUMB[37][26] ,
         \mult_22/SUMB[37][27] , \mult_22/SUMB[37][28] ,
         \mult_22/SUMB[37][29] , \mult_22/SUMB[37][30] ,
         \mult_22/SUMB[37][31] , \mult_22/SUMB[37][32] ,
         \mult_22/SUMB[37][33] , \mult_22/SUMB[37][34] ,
         \mult_22/SUMB[37][35] , \mult_22/SUMB[37][36] ,
         \mult_22/SUMB[37][37] , \mult_22/SUMB[37][38] ,
         \mult_22/SUMB[37][39] , \mult_22/SUMB[37][40] ,
         \mult_22/SUMB[37][41] , \mult_22/SUMB[37][42] ,
         \mult_22/SUMB[37][43] , \mult_22/SUMB[37][44] ,
         \mult_22/SUMB[37][45] , \mult_22/SUMB[37][46] ,
         \mult_22/SUMB[37][47] , \mult_22/SUMB[37][48] ,
         \mult_22/SUMB[37][49] , \mult_22/SUMB[37][50] ,
         \mult_22/SUMB[37][51] , \mult_22/SUMB[37][52] ,
         \mult_22/SUMB[37][53] , \mult_22/SUMB[37][54] ,
         \mult_22/SUMB[37][55] , \mult_22/SUMB[37][56] ,
         \mult_22/SUMB[37][57] , \mult_22/SUMB[37][58] ,
         \mult_22/SUMB[37][59] , \mult_22/SUMB[37][60] ,
         \mult_22/SUMB[37][61] , \mult_22/SUMB[37][62] , \mult_22/SUMB[38][1] ,
         \mult_22/SUMB[38][2] , \mult_22/SUMB[38][3] , \mult_22/SUMB[38][4] ,
         \mult_22/SUMB[38][5] , \mult_22/SUMB[38][6] , \mult_22/SUMB[38][7] ,
         \mult_22/SUMB[38][8] , \mult_22/SUMB[38][9] , \mult_22/SUMB[38][10] ,
         \mult_22/SUMB[38][11] , \mult_22/SUMB[38][12] ,
         \mult_22/SUMB[38][13] , \mult_22/SUMB[38][14] ,
         \mult_22/SUMB[38][15] , \mult_22/SUMB[38][16] ,
         \mult_22/SUMB[38][17] , \mult_22/SUMB[38][18] ,
         \mult_22/SUMB[38][19] , \mult_22/SUMB[38][20] ,
         \mult_22/SUMB[38][21] , \mult_22/SUMB[38][22] ,
         \mult_22/SUMB[38][23] , \mult_22/SUMB[38][24] ,
         \mult_22/SUMB[38][25] , \mult_22/SUMB[38][26] ,
         \mult_22/SUMB[38][27] , \mult_22/SUMB[38][28] ,
         \mult_22/SUMB[38][29] , \mult_22/SUMB[38][30] ,
         \mult_22/SUMB[38][31] , \mult_22/SUMB[38][32] ,
         \mult_22/SUMB[38][33] , \mult_22/SUMB[38][34] ,
         \mult_22/SUMB[38][35] , \mult_22/SUMB[38][36] ,
         \mult_22/SUMB[38][37] , \mult_22/SUMB[38][38] ,
         \mult_22/SUMB[38][39] , \mult_22/SUMB[38][40] ,
         \mult_22/SUMB[38][41] , \mult_22/SUMB[38][42] ,
         \mult_22/SUMB[38][43] , \mult_22/SUMB[38][44] ,
         \mult_22/SUMB[38][45] , \mult_22/SUMB[38][46] ,
         \mult_22/SUMB[38][47] , \mult_22/SUMB[38][48] ,
         \mult_22/SUMB[38][49] , \mult_22/SUMB[38][50] ,
         \mult_22/SUMB[38][51] , \mult_22/SUMB[38][52] ,
         \mult_22/SUMB[38][53] , \mult_22/SUMB[38][54] ,
         \mult_22/SUMB[38][55] , \mult_22/SUMB[38][56] ,
         \mult_22/SUMB[38][57] , \mult_22/SUMB[38][58] ,
         \mult_22/SUMB[38][59] , \mult_22/SUMB[38][60] ,
         \mult_22/SUMB[38][61] , \mult_22/SUMB[38][62] , \mult_22/SUMB[39][1] ,
         \mult_22/SUMB[39][2] , \mult_22/SUMB[39][3] , \mult_22/SUMB[39][4] ,
         \mult_22/SUMB[39][5] , \mult_22/SUMB[39][6] , \mult_22/SUMB[39][7] ,
         \mult_22/SUMB[39][8] , \mult_22/SUMB[39][9] , \mult_22/SUMB[39][10] ,
         \mult_22/SUMB[39][11] , \mult_22/SUMB[39][12] ,
         \mult_22/SUMB[39][13] , \mult_22/SUMB[39][14] ,
         \mult_22/SUMB[39][15] , \mult_22/SUMB[39][16] ,
         \mult_22/SUMB[39][17] , \mult_22/SUMB[39][18] ,
         \mult_22/SUMB[39][19] , \mult_22/SUMB[39][20] ,
         \mult_22/SUMB[39][21] , \mult_22/SUMB[39][22] ,
         \mult_22/SUMB[39][23] , \mult_22/SUMB[39][24] ,
         \mult_22/SUMB[39][25] , \mult_22/SUMB[39][26] ,
         \mult_22/SUMB[39][27] , \mult_22/SUMB[39][28] ,
         \mult_22/SUMB[39][29] , \mult_22/SUMB[39][30] ,
         \mult_22/SUMB[39][31] , \mult_22/SUMB[39][32] ,
         \mult_22/SUMB[39][33] , \mult_22/SUMB[39][34] ,
         \mult_22/SUMB[39][35] , \mult_22/SUMB[39][36] ,
         \mult_22/SUMB[39][37] , \mult_22/SUMB[39][38] ,
         \mult_22/SUMB[39][39] , \mult_22/SUMB[39][40] ,
         \mult_22/SUMB[39][41] , \mult_22/SUMB[39][42] ,
         \mult_22/SUMB[39][43] , \mult_22/SUMB[39][44] ,
         \mult_22/SUMB[39][45] , \mult_22/SUMB[39][46] ,
         \mult_22/SUMB[39][47] , \mult_22/SUMB[39][48] ,
         \mult_22/SUMB[39][49] , \mult_22/SUMB[39][50] ,
         \mult_22/SUMB[39][51] , \mult_22/SUMB[39][52] ,
         \mult_22/SUMB[39][53] , \mult_22/SUMB[39][54] ,
         \mult_22/SUMB[39][55] , \mult_22/SUMB[39][56] ,
         \mult_22/SUMB[39][57] , \mult_22/SUMB[39][58] ,
         \mult_22/SUMB[39][59] , \mult_22/SUMB[39][60] ,
         \mult_22/SUMB[39][61] , \mult_22/SUMB[39][62] ,
         \mult_22/CARRYB[32][0] , \mult_22/CARRYB[32][1] ,
         \mult_22/CARRYB[32][2] , \mult_22/CARRYB[32][3] ,
         \mult_22/CARRYB[32][4] , \mult_22/CARRYB[32][5] ,
         \mult_22/CARRYB[32][6] , \mult_22/CARRYB[32][7] ,
         \mult_22/CARRYB[32][8] , \mult_22/CARRYB[32][9] ,
         \mult_22/CARRYB[32][10] , \mult_22/CARRYB[32][11] ,
         \mult_22/CARRYB[32][12] , \mult_22/CARRYB[32][13] ,
         \mult_22/CARRYB[32][14] , \mult_22/CARRYB[32][15] ,
         \mult_22/CARRYB[32][16] , \mult_22/CARRYB[32][17] ,
         \mult_22/CARRYB[32][18] , \mult_22/CARRYB[32][19] ,
         \mult_22/CARRYB[32][20] , \mult_22/CARRYB[32][21] ,
         \mult_22/CARRYB[32][22] , \mult_22/CARRYB[32][23] ,
         \mult_22/CARRYB[32][24] , \mult_22/CARRYB[32][25] ,
         \mult_22/CARRYB[32][26] , \mult_22/CARRYB[32][27] ,
         \mult_22/CARRYB[32][28] , \mult_22/CARRYB[32][29] ,
         \mult_22/CARRYB[32][30] , \mult_22/CARRYB[32][31] ,
         \mult_22/CARRYB[32][32] , \mult_22/CARRYB[32][33] ,
         \mult_22/CARRYB[32][34] , \mult_22/CARRYB[32][35] ,
         \mult_22/CARRYB[32][36] , \mult_22/CARRYB[32][37] ,
         \mult_22/CARRYB[32][38] , \mult_22/CARRYB[32][39] ,
         \mult_22/CARRYB[32][40] , \mult_22/CARRYB[32][41] ,
         \mult_22/CARRYB[32][42] , \mult_22/CARRYB[32][43] ,
         \mult_22/CARRYB[32][44] , \mult_22/CARRYB[32][45] ,
         \mult_22/CARRYB[32][46] , \mult_22/CARRYB[32][47] ,
         \mult_22/CARRYB[32][48] , \mult_22/CARRYB[32][49] ,
         \mult_22/CARRYB[32][50] , \mult_22/CARRYB[32][51] ,
         \mult_22/CARRYB[32][52] , \mult_22/CARRYB[32][53] ,
         \mult_22/CARRYB[32][54] , \mult_22/CARRYB[32][55] ,
         \mult_22/CARRYB[32][56] , \mult_22/CARRYB[32][57] ,
         \mult_22/CARRYB[32][58] , \mult_22/CARRYB[32][59] ,
         \mult_22/CARRYB[32][60] , \mult_22/CARRYB[32][61] ,
         \mult_22/CARRYB[32][62] , \mult_22/CARRYB[33][0] ,
         \mult_22/CARRYB[33][1] , \mult_22/CARRYB[33][2] ,
         \mult_22/CARRYB[33][3] , \mult_22/CARRYB[33][4] ,
         \mult_22/CARRYB[33][5] , \mult_22/CARRYB[33][6] ,
         \mult_22/CARRYB[33][7] , \mult_22/CARRYB[33][8] ,
         \mult_22/CARRYB[33][9] , \mult_22/CARRYB[33][10] ,
         \mult_22/CARRYB[33][11] , \mult_22/CARRYB[33][12] ,
         \mult_22/CARRYB[33][13] , \mult_22/CARRYB[33][14] ,
         \mult_22/CARRYB[33][15] , \mult_22/CARRYB[33][16] ,
         \mult_22/CARRYB[33][17] , \mult_22/CARRYB[33][18] ,
         \mult_22/CARRYB[33][19] , \mult_22/CARRYB[33][20] ,
         \mult_22/CARRYB[33][21] , \mult_22/CARRYB[33][22] ,
         \mult_22/CARRYB[33][23] , \mult_22/CARRYB[33][24] ,
         \mult_22/CARRYB[33][25] , \mult_22/CARRYB[33][26] ,
         \mult_22/CARRYB[33][27] , \mult_22/CARRYB[33][28] ,
         \mult_22/CARRYB[33][29] , \mult_22/CARRYB[33][30] ,
         \mult_22/CARRYB[33][31] , \mult_22/CARRYB[33][32] ,
         \mult_22/CARRYB[33][33] , \mult_22/CARRYB[33][34] ,
         \mult_22/CARRYB[33][35] , \mult_22/CARRYB[33][36] ,
         \mult_22/CARRYB[33][37] , \mult_22/CARRYB[33][38] ,
         \mult_22/CARRYB[33][39] , \mult_22/CARRYB[33][40] ,
         \mult_22/CARRYB[33][41] , \mult_22/CARRYB[33][42] ,
         \mult_22/CARRYB[33][43] , \mult_22/CARRYB[33][44] ,
         \mult_22/CARRYB[33][45] , \mult_22/CARRYB[33][46] ,
         \mult_22/CARRYB[33][47] , \mult_22/CARRYB[33][48] ,
         \mult_22/CARRYB[33][49] , \mult_22/CARRYB[33][50] ,
         \mult_22/CARRYB[33][51] , \mult_22/CARRYB[33][52] ,
         \mult_22/CARRYB[33][53] , \mult_22/CARRYB[33][54] ,
         \mult_22/CARRYB[33][55] , \mult_22/CARRYB[33][56] ,
         \mult_22/CARRYB[33][57] , \mult_22/CARRYB[33][58] ,
         \mult_22/CARRYB[33][59] , \mult_22/CARRYB[33][60] ,
         \mult_22/CARRYB[33][61] , \mult_22/CARRYB[33][62] ,
         \mult_22/CARRYB[34][0] , \mult_22/CARRYB[34][1] ,
         \mult_22/CARRYB[34][2] , \mult_22/CARRYB[34][3] ,
         \mult_22/CARRYB[34][4] , \mult_22/CARRYB[34][5] ,
         \mult_22/CARRYB[34][6] , \mult_22/CARRYB[34][7] ,
         \mult_22/CARRYB[34][8] , \mult_22/CARRYB[34][9] ,
         \mult_22/CARRYB[34][10] , \mult_22/CARRYB[34][11] ,
         \mult_22/CARRYB[34][12] , \mult_22/CARRYB[34][13] ,
         \mult_22/CARRYB[34][14] , \mult_22/CARRYB[34][15] ,
         \mult_22/CARRYB[34][16] , \mult_22/CARRYB[34][17] ,
         \mult_22/CARRYB[34][18] , \mult_22/CARRYB[34][19] ,
         \mult_22/CARRYB[34][20] , \mult_22/CARRYB[34][21] ,
         \mult_22/CARRYB[34][22] , \mult_22/CARRYB[34][23] ,
         \mult_22/CARRYB[34][24] , \mult_22/CARRYB[34][25] ,
         \mult_22/CARRYB[34][26] , \mult_22/CARRYB[34][27] ,
         \mult_22/CARRYB[34][28] , \mult_22/CARRYB[34][29] ,
         \mult_22/CARRYB[34][30] , \mult_22/CARRYB[34][31] ,
         \mult_22/CARRYB[34][32] , \mult_22/CARRYB[34][33] ,
         \mult_22/CARRYB[34][34] , \mult_22/CARRYB[34][35] ,
         \mult_22/CARRYB[34][36] , \mult_22/CARRYB[34][37] ,
         \mult_22/CARRYB[34][38] , \mult_22/CARRYB[34][39] ,
         \mult_22/CARRYB[34][40] , \mult_22/CARRYB[34][41] ,
         \mult_22/CARRYB[34][42] , \mult_22/CARRYB[34][43] ,
         \mult_22/CARRYB[34][44] , \mult_22/CARRYB[34][45] ,
         \mult_22/CARRYB[34][46] , \mult_22/CARRYB[34][47] ,
         \mult_22/CARRYB[34][48] , \mult_22/CARRYB[34][49] ,
         \mult_22/CARRYB[34][50] , \mult_22/CARRYB[34][51] ,
         \mult_22/CARRYB[34][52] , \mult_22/CARRYB[34][53] ,
         \mult_22/CARRYB[34][54] , \mult_22/CARRYB[34][55] ,
         \mult_22/CARRYB[34][56] , \mult_22/CARRYB[34][57] ,
         \mult_22/CARRYB[34][58] , \mult_22/CARRYB[34][59] ,
         \mult_22/CARRYB[34][60] , \mult_22/CARRYB[34][61] ,
         \mult_22/CARRYB[34][62] , \mult_22/CARRYB[35][0] ,
         \mult_22/CARRYB[35][1] , \mult_22/CARRYB[35][2] ,
         \mult_22/CARRYB[35][3] , \mult_22/CARRYB[35][4] ,
         \mult_22/CARRYB[35][5] , \mult_22/CARRYB[35][6] ,
         \mult_22/CARRYB[35][7] , \mult_22/CARRYB[35][8] ,
         \mult_22/CARRYB[35][9] , \mult_22/CARRYB[35][10] ,
         \mult_22/CARRYB[35][11] , \mult_22/CARRYB[35][12] ,
         \mult_22/CARRYB[35][13] , \mult_22/CARRYB[35][14] ,
         \mult_22/CARRYB[35][15] , \mult_22/CARRYB[35][16] ,
         \mult_22/CARRYB[35][17] , \mult_22/CARRYB[35][18] ,
         \mult_22/CARRYB[35][19] , \mult_22/CARRYB[35][20] ,
         \mult_22/CARRYB[35][21] , \mult_22/CARRYB[35][22] ,
         \mult_22/CARRYB[35][23] , \mult_22/CARRYB[35][24] ,
         \mult_22/CARRYB[35][25] , \mult_22/CARRYB[35][26] ,
         \mult_22/CARRYB[35][27] , \mult_22/CARRYB[35][28] ,
         \mult_22/CARRYB[35][29] , \mult_22/CARRYB[35][30] ,
         \mult_22/CARRYB[35][31] , \mult_22/CARRYB[35][32] ,
         \mult_22/CARRYB[35][33] , \mult_22/CARRYB[35][34] ,
         \mult_22/CARRYB[35][35] , \mult_22/CARRYB[35][36] ,
         \mult_22/CARRYB[35][37] , \mult_22/CARRYB[35][38] ,
         \mult_22/CARRYB[35][39] , \mult_22/CARRYB[35][40] ,
         \mult_22/CARRYB[35][41] , \mult_22/CARRYB[35][42] ,
         \mult_22/CARRYB[35][43] , \mult_22/CARRYB[35][44] ,
         \mult_22/CARRYB[35][45] , \mult_22/CARRYB[35][46] ,
         \mult_22/CARRYB[35][47] , \mult_22/CARRYB[35][48] ,
         \mult_22/CARRYB[35][49] , \mult_22/CARRYB[35][50] ,
         \mult_22/CARRYB[35][51] , \mult_22/CARRYB[35][52] ,
         \mult_22/CARRYB[35][53] , \mult_22/CARRYB[35][54] ,
         \mult_22/CARRYB[35][55] , \mult_22/CARRYB[35][56] ,
         \mult_22/CARRYB[35][57] , \mult_22/CARRYB[35][58] ,
         \mult_22/CARRYB[35][59] , \mult_22/CARRYB[35][60] ,
         \mult_22/CARRYB[35][61] , \mult_22/CARRYB[35][62] ,
         \mult_22/CARRYB[36][0] , \mult_22/CARRYB[36][1] ,
         \mult_22/CARRYB[36][2] , \mult_22/CARRYB[36][3] ,
         \mult_22/CARRYB[36][4] , \mult_22/CARRYB[36][5] ,
         \mult_22/CARRYB[36][6] , \mult_22/CARRYB[36][7] ,
         \mult_22/CARRYB[36][8] , \mult_22/CARRYB[36][9] ,
         \mult_22/CARRYB[36][10] , \mult_22/CARRYB[36][11] ,
         \mult_22/CARRYB[36][12] , \mult_22/CARRYB[36][13] ,
         \mult_22/CARRYB[36][14] , \mult_22/CARRYB[36][15] ,
         \mult_22/CARRYB[36][16] , \mult_22/CARRYB[36][17] ,
         \mult_22/CARRYB[36][18] , \mult_22/CARRYB[36][19] ,
         \mult_22/CARRYB[36][20] , \mult_22/CARRYB[36][21] ,
         \mult_22/CARRYB[36][22] , \mult_22/CARRYB[36][23] ,
         \mult_22/CARRYB[36][24] , \mult_22/CARRYB[36][25] ,
         \mult_22/CARRYB[36][26] , \mult_22/CARRYB[36][27] ,
         \mult_22/CARRYB[36][28] , \mult_22/CARRYB[36][29] ,
         \mult_22/CARRYB[36][30] , \mult_22/CARRYB[36][31] ,
         \mult_22/CARRYB[36][32] , \mult_22/CARRYB[36][33] ,
         \mult_22/CARRYB[36][34] , \mult_22/CARRYB[36][35] ,
         \mult_22/CARRYB[36][36] , \mult_22/CARRYB[36][37] ,
         \mult_22/CARRYB[36][38] , \mult_22/CARRYB[36][39] ,
         \mult_22/CARRYB[36][40] , \mult_22/CARRYB[36][41] ,
         \mult_22/CARRYB[36][42] , \mult_22/CARRYB[36][43] ,
         \mult_22/CARRYB[36][44] , \mult_22/CARRYB[36][45] ,
         \mult_22/CARRYB[36][46] , \mult_22/CARRYB[36][47] ,
         \mult_22/CARRYB[36][48] , \mult_22/CARRYB[36][49] ,
         \mult_22/CARRYB[36][50] , \mult_22/CARRYB[36][51] ,
         \mult_22/CARRYB[36][52] , \mult_22/CARRYB[36][53] ,
         \mult_22/CARRYB[36][54] , \mult_22/CARRYB[36][55] ,
         \mult_22/CARRYB[36][56] , \mult_22/CARRYB[36][57] ,
         \mult_22/CARRYB[36][58] , \mult_22/CARRYB[36][59] ,
         \mult_22/CARRYB[36][60] , \mult_22/CARRYB[36][61] ,
         \mult_22/CARRYB[36][62] , \mult_22/CARRYB[37][0] ,
         \mult_22/CARRYB[37][1] , \mult_22/CARRYB[37][2] ,
         \mult_22/CARRYB[37][3] , \mult_22/CARRYB[37][4] ,
         \mult_22/CARRYB[37][5] , \mult_22/CARRYB[37][6] ,
         \mult_22/CARRYB[37][7] , \mult_22/CARRYB[37][8] ,
         \mult_22/CARRYB[37][9] , \mult_22/CARRYB[37][10] ,
         \mult_22/CARRYB[37][11] , \mult_22/CARRYB[37][12] ,
         \mult_22/CARRYB[37][13] , \mult_22/CARRYB[37][14] ,
         \mult_22/CARRYB[37][15] , \mult_22/CARRYB[37][16] ,
         \mult_22/CARRYB[37][17] , \mult_22/CARRYB[37][18] ,
         \mult_22/CARRYB[37][19] , \mult_22/CARRYB[37][20] ,
         \mult_22/CARRYB[37][21] , \mult_22/CARRYB[37][22] ,
         \mult_22/CARRYB[37][23] , \mult_22/CARRYB[37][24] ,
         \mult_22/CARRYB[37][25] , \mult_22/CARRYB[37][26] ,
         \mult_22/CARRYB[37][27] , \mult_22/CARRYB[37][28] ,
         \mult_22/CARRYB[37][29] , \mult_22/CARRYB[37][30] ,
         \mult_22/CARRYB[37][31] , \mult_22/CARRYB[37][32] ,
         \mult_22/CARRYB[37][33] , \mult_22/CARRYB[37][34] ,
         \mult_22/CARRYB[37][35] , \mult_22/CARRYB[37][36] ,
         \mult_22/CARRYB[37][37] , \mult_22/CARRYB[37][38] ,
         \mult_22/CARRYB[37][39] , \mult_22/CARRYB[37][40] ,
         \mult_22/CARRYB[37][41] , \mult_22/CARRYB[37][42] ,
         \mult_22/CARRYB[37][43] , \mult_22/CARRYB[37][44] ,
         \mult_22/CARRYB[37][45] , \mult_22/CARRYB[37][46] ,
         \mult_22/CARRYB[37][47] , \mult_22/CARRYB[37][48] ,
         \mult_22/CARRYB[37][49] , \mult_22/CARRYB[37][50] ,
         \mult_22/CARRYB[37][51] , \mult_22/CARRYB[37][52] ,
         \mult_22/CARRYB[37][53] , \mult_22/CARRYB[37][54] ,
         \mult_22/CARRYB[37][55] , \mult_22/CARRYB[37][56] ,
         \mult_22/CARRYB[37][57] , \mult_22/CARRYB[37][58] ,
         \mult_22/CARRYB[37][59] , \mult_22/CARRYB[37][60] ,
         \mult_22/CARRYB[37][61] , \mult_22/CARRYB[37][62] ,
         \mult_22/CARRYB[38][0] , \mult_22/CARRYB[38][1] ,
         \mult_22/CARRYB[38][2] , \mult_22/CARRYB[38][3] ,
         \mult_22/CARRYB[38][4] , \mult_22/CARRYB[38][5] ,
         \mult_22/CARRYB[38][6] , \mult_22/CARRYB[38][7] ,
         \mult_22/CARRYB[38][8] , \mult_22/CARRYB[38][9] ,
         \mult_22/CARRYB[38][10] , \mult_22/CARRYB[38][11] ,
         \mult_22/CARRYB[38][12] , \mult_22/CARRYB[38][13] ,
         \mult_22/CARRYB[38][14] , \mult_22/CARRYB[38][15] ,
         \mult_22/CARRYB[38][16] , \mult_22/CARRYB[38][17] ,
         \mult_22/CARRYB[38][18] , \mult_22/CARRYB[38][19] ,
         \mult_22/CARRYB[38][20] , \mult_22/CARRYB[38][21] ,
         \mult_22/CARRYB[38][22] , \mult_22/CARRYB[38][23] ,
         \mult_22/CARRYB[38][24] , \mult_22/CARRYB[38][25] ,
         \mult_22/CARRYB[38][26] , \mult_22/CARRYB[38][27] ,
         \mult_22/CARRYB[38][28] , \mult_22/CARRYB[38][29] ,
         \mult_22/CARRYB[38][30] , \mult_22/CARRYB[38][31] ,
         \mult_22/CARRYB[38][32] , \mult_22/CARRYB[38][33] ,
         \mult_22/CARRYB[38][34] , \mult_22/CARRYB[38][35] ,
         \mult_22/CARRYB[38][36] , \mult_22/CARRYB[38][37] ,
         \mult_22/CARRYB[38][38] , \mult_22/CARRYB[38][39] ,
         \mult_22/CARRYB[38][40] , \mult_22/CARRYB[38][41] ,
         \mult_22/CARRYB[38][42] , \mult_22/CARRYB[38][43] ,
         \mult_22/CARRYB[38][44] , \mult_22/CARRYB[38][45] ,
         \mult_22/CARRYB[38][46] , \mult_22/CARRYB[38][47] ,
         \mult_22/CARRYB[38][48] , \mult_22/CARRYB[38][49] ,
         \mult_22/CARRYB[38][50] , \mult_22/CARRYB[38][51] ,
         \mult_22/CARRYB[38][52] , \mult_22/CARRYB[38][53] ,
         \mult_22/CARRYB[38][54] , \mult_22/CARRYB[38][55] ,
         \mult_22/CARRYB[38][56] , \mult_22/CARRYB[38][57] ,
         \mult_22/CARRYB[38][58] , \mult_22/CARRYB[38][59] ,
         \mult_22/CARRYB[38][60] , \mult_22/CARRYB[38][61] ,
         \mult_22/CARRYB[38][62] , \mult_22/CARRYB[39][0] ,
         \mult_22/CARRYB[39][1] , \mult_22/CARRYB[39][2] ,
         \mult_22/CARRYB[39][3] , \mult_22/CARRYB[39][4] ,
         \mult_22/CARRYB[39][5] , \mult_22/CARRYB[39][6] ,
         \mult_22/CARRYB[39][7] , \mult_22/CARRYB[39][8] ,
         \mult_22/CARRYB[39][9] , \mult_22/CARRYB[39][10] ,
         \mult_22/CARRYB[39][11] , \mult_22/CARRYB[39][12] ,
         \mult_22/CARRYB[39][13] , \mult_22/CARRYB[39][14] ,
         \mult_22/CARRYB[39][15] , \mult_22/CARRYB[39][16] ,
         \mult_22/CARRYB[39][17] , \mult_22/CARRYB[39][18] ,
         \mult_22/CARRYB[39][19] , \mult_22/CARRYB[39][20] ,
         \mult_22/CARRYB[39][21] , \mult_22/CARRYB[39][22] ,
         \mult_22/CARRYB[39][23] , \mult_22/CARRYB[39][24] ,
         \mult_22/CARRYB[39][25] , \mult_22/CARRYB[39][26] ,
         \mult_22/CARRYB[39][27] , \mult_22/CARRYB[39][28] ,
         \mult_22/CARRYB[39][29] , \mult_22/CARRYB[39][30] ,
         \mult_22/CARRYB[39][31] , \mult_22/CARRYB[39][32] ,
         \mult_22/CARRYB[39][33] , \mult_22/CARRYB[39][34] ,
         \mult_22/CARRYB[39][35] , \mult_22/CARRYB[39][36] ,
         \mult_22/CARRYB[39][37] , \mult_22/CARRYB[39][38] ,
         \mult_22/CARRYB[39][39] , \mult_22/CARRYB[39][40] ,
         \mult_22/CARRYB[39][41] , \mult_22/CARRYB[39][42] ,
         \mult_22/CARRYB[39][43] , \mult_22/CARRYB[39][44] ,
         \mult_22/CARRYB[39][45] , \mult_22/CARRYB[39][46] ,
         \mult_22/CARRYB[39][47] , \mult_22/CARRYB[39][48] ,
         \mult_22/CARRYB[39][49] , \mult_22/CARRYB[39][50] ,
         \mult_22/CARRYB[39][51] , \mult_22/CARRYB[39][52] ,
         \mult_22/CARRYB[39][53] , \mult_22/CARRYB[39][54] ,
         \mult_22/CARRYB[39][55] , \mult_22/CARRYB[39][56] ,
         \mult_22/CARRYB[39][57] , \mult_22/CARRYB[39][58] ,
         \mult_22/CARRYB[39][59] , \mult_22/CARRYB[39][60] ,
         \mult_22/CARRYB[39][61] , \mult_22/CARRYB[39][62] ,
         \mult_22/SUMB[24][1] , \mult_22/SUMB[24][2] , \mult_22/SUMB[24][3] ,
         \mult_22/SUMB[24][4] , \mult_22/SUMB[24][5] , \mult_22/SUMB[24][6] ,
         \mult_22/SUMB[24][7] , \mult_22/SUMB[24][8] , \mult_22/SUMB[24][9] ,
         \mult_22/SUMB[24][10] , \mult_22/SUMB[24][11] ,
         \mult_22/SUMB[24][12] , \mult_22/SUMB[24][13] ,
         \mult_22/SUMB[24][14] , \mult_22/SUMB[24][15] ,
         \mult_22/SUMB[24][16] , \mult_22/SUMB[24][17] ,
         \mult_22/SUMB[24][18] , \mult_22/SUMB[24][19] ,
         \mult_22/SUMB[24][20] , \mult_22/SUMB[24][21] ,
         \mult_22/SUMB[24][22] , \mult_22/SUMB[24][23] ,
         \mult_22/SUMB[24][24] , \mult_22/SUMB[24][25] ,
         \mult_22/SUMB[24][26] , \mult_22/SUMB[24][27] ,
         \mult_22/SUMB[24][28] , \mult_22/SUMB[24][29] ,
         \mult_22/SUMB[24][30] , \mult_22/SUMB[24][31] ,
         \mult_22/SUMB[24][32] , \mult_22/SUMB[24][33] ,
         \mult_22/SUMB[24][34] , \mult_22/SUMB[24][35] ,
         \mult_22/SUMB[24][36] , \mult_22/SUMB[24][37] ,
         \mult_22/SUMB[24][38] , \mult_22/SUMB[24][39] ,
         \mult_22/SUMB[24][40] , \mult_22/SUMB[24][41] ,
         \mult_22/SUMB[24][42] , \mult_22/SUMB[24][43] ,
         \mult_22/SUMB[24][44] , \mult_22/SUMB[24][45] ,
         \mult_22/SUMB[24][46] , \mult_22/SUMB[24][47] ,
         \mult_22/SUMB[24][48] , \mult_22/SUMB[24][49] ,
         \mult_22/SUMB[24][50] , \mult_22/SUMB[24][51] ,
         \mult_22/SUMB[24][52] , \mult_22/SUMB[24][53] ,
         \mult_22/SUMB[24][54] , \mult_22/SUMB[24][55] ,
         \mult_22/SUMB[24][56] , \mult_22/SUMB[24][57] ,
         \mult_22/SUMB[24][58] , \mult_22/SUMB[24][59] ,
         \mult_22/SUMB[24][60] , \mult_22/SUMB[24][61] ,
         \mult_22/SUMB[24][62] , \mult_22/SUMB[25][1] , \mult_22/SUMB[25][2] ,
         \mult_22/SUMB[25][3] , \mult_22/SUMB[25][4] , \mult_22/SUMB[25][5] ,
         \mult_22/SUMB[25][6] , \mult_22/SUMB[25][7] , \mult_22/SUMB[25][8] ,
         \mult_22/SUMB[25][9] , \mult_22/SUMB[25][10] , \mult_22/SUMB[25][11] ,
         \mult_22/SUMB[25][12] , \mult_22/SUMB[25][13] ,
         \mult_22/SUMB[25][14] , \mult_22/SUMB[25][15] ,
         \mult_22/SUMB[25][16] , \mult_22/SUMB[25][17] ,
         \mult_22/SUMB[25][18] , \mult_22/SUMB[25][19] ,
         \mult_22/SUMB[25][20] , \mult_22/SUMB[25][21] ,
         \mult_22/SUMB[25][22] , \mult_22/SUMB[25][23] ,
         \mult_22/SUMB[25][24] , \mult_22/SUMB[25][25] ,
         \mult_22/SUMB[25][26] , \mult_22/SUMB[25][27] ,
         \mult_22/SUMB[25][28] , \mult_22/SUMB[25][29] ,
         \mult_22/SUMB[25][30] , \mult_22/SUMB[25][31] ,
         \mult_22/SUMB[25][32] , \mult_22/SUMB[25][33] ,
         \mult_22/SUMB[25][34] , \mult_22/SUMB[25][36] ,
         \mult_22/SUMB[25][37] , \mult_22/SUMB[25][38] ,
         \mult_22/SUMB[25][39] , \mult_22/SUMB[25][40] ,
         \mult_22/SUMB[25][41] , \mult_22/SUMB[25][42] ,
         \mult_22/SUMB[25][43] , \mult_22/SUMB[25][44] ,
         \mult_22/SUMB[25][45] , \mult_22/SUMB[25][46] ,
         \mult_22/SUMB[25][47] , \mult_22/SUMB[25][48] ,
         \mult_22/SUMB[25][49] , \mult_22/SUMB[25][50] ,
         \mult_22/SUMB[25][51] , \mult_22/SUMB[25][52] ,
         \mult_22/SUMB[25][53] , \mult_22/SUMB[25][54] ,
         \mult_22/SUMB[25][55] , \mult_22/SUMB[25][56] ,
         \mult_22/SUMB[25][57] , \mult_22/SUMB[25][58] ,
         \mult_22/SUMB[25][59] , \mult_22/SUMB[25][60] ,
         \mult_22/SUMB[25][61] , \mult_22/SUMB[25][62] , \mult_22/SUMB[26][1] ,
         \mult_22/SUMB[26][2] , \mult_22/SUMB[26][3] , \mult_22/SUMB[26][4] ,
         \mult_22/SUMB[26][5] , \mult_22/SUMB[26][6] , \mult_22/SUMB[26][7] ,
         \mult_22/SUMB[26][8] , \mult_22/SUMB[26][9] , \mult_22/SUMB[26][10] ,
         \mult_22/SUMB[26][11] , \mult_22/SUMB[26][12] ,
         \mult_22/SUMB[26][13] , \mult_22/SUMB[26][14] ,
         \mult_22/SUMB[26][15] , \mult_22/SUMB[26][16] ,
         \mult_22/SUMB[26][17] , \mult_22/SUMB[26][18] ,
         \mult_22/SUMB[26][19] , \mult_22/SUMB[26][20] ,
         \mult_22/SUMB[26][21] , \mult_22/SUMB[26][22] ,
         \mult_22/SUMB[26][23] , \mult_22/SUMB[26][24] ,
         \mult_22/SUMB[26][25] , \mult_22/SUMB[26][26] ,
         \mult_22/SUMB[26][27] , \mult_22/SUMB[26][28] ,
         \mult_22/SUMB[26][29] , \mult_22/SUMB[26][30] ,
         \mult_22/SUMB[26][31] , \mult_22/SUMB[26][32] ,
         \mult_22/SUMB[26][33] , \mult_22/SUMB[26][34] ,
         \mult_22/SUMB[26][35] , \mult_22/SUMB[26][36] ,
         \mult_22/SUMB[26][37] , \mult_22/SUMB[26][38] ,
         \mult_22/SUMB[26][39] , \mult_22/SUMB[26][40] ,
         \mult_22/SUMB[26][41] , \mult_22/SUMB[26][42] ,
         \mult_22/SUMB[26][43] , \mult_22/SUMB[26][44] ,
         \mult_22/SUMB[26][45] , \mult_22/SUMB[26][46] ,
         \mult_22/SUMB[26][47] , \mult_22/SUMB[26][48] ,
         \mult_22/SUMB[26][49] , \mult_22/SUMB[26][50] ,
         \mult_22/SUMB[26][51] , \mult_22/SUMB[26][52] ,
         \mult_22/SUMB[26][53] , \mult_22/SUMB[26][54] ,
         \mult_22/SUMB[26][55] , \mult_22/SUMB[26][56] ,
         \mult_22/SUMB[26][57] , \mult_22/SUMB[26][58] ,
         \mult_22/SUMB[26][59] , \mult_22/SUMB[26][60] ,
         \mult_22/SUMB[26][61] , \mult_22/SUMB[26][62] , \mult_22/SUMB[27][1] ,
         \mult_22/SUMB[27][2] , \mult_22/SUMB[27][3] , \mult_22/SUMB[27][4] ,
         \mult_22/SUMB[27][5] , \mult_22/SUMB[27][6] , \mult_22/SUMB[27][7] ,
         \mult_22/SUMB[27][8] , \mult_22/SUMB[27][9] , \mult_22/SUMB[27][10] ,
         \mult_22/SUMB[27][11] , \mult_22/SUMB[27][12] ,
         \mult_22/SUMB[27][13] , \mult_22/SUMB[27][14] ,
         \mult_22/SUMB[27][15] , \mult_22/SUMB[27][16] ,
         \mult_22/SUMB[27][17] , \mult_22/SUMB[27][18] ,
         \mult_22/SUMB[27][19] , \mult_22/SUMB[27][20] ,
         \mult_22/SUMB[27][21] , \mult_22/SUMB[27][22] ,
         \mult_22/SUMB[27][23] , \mult_22/SUMB[27][24] ,
         \mult_22/SUMB[27][25] , \mult_22/SUMB[27][26] ,
         \mult_22/SUMB[27][27] , \mult_22/SUMB[27][28] ,
         \mult_22/SUMB[27][29] , \mult_22/SUMB[27][30] ,
         \mult_22/SUMB[27][31] , \mult_22/SUMB[27][32] ,
         \mult_22/SUMB[27][33] , \mult_22/SUMB[27][34] ,
         \mult_22/SUMB[27][35] , \mult_22/SUMB[27][36] ,
         \mult_22/SUMB[27][37] , \mult_22/SUMB[27][38] ,
         \mult_22/SUMB[27][39] , \mult_22/SUMB[27][40] ,
         \mult_22/SUMB[27][41] , \mult_22/SUMB[27][42] ,
         \mult_22/SUMB[27][43] , \mult_22/SUMB[27][44] ,
         \mult_22/SUMB[27][45] , \mult_22/SUMB[27][46] ,
         \mult_22/SUMB[27][47] , \mult_22/SUMB[27][48] ,
         \mult_22/SUMB[27][49] , \mult_22/SUMB[27][50] ,
         \mult_22/SUMB[27][51] , \mult_22/SUMB[27][52] ,
         \mult_22/SUMB[27][53] , \mult_22/SUMB[27][54] ,
         \mult_22/SUMB[27][55] , \mult_22/SUMB[27][56] ,
         \mult_22/SUMB[27][57] , \mult_22/SUMB[27][58] ,
         \mult_22/SUMB[27][59] , \mult_22/SUMB[27][60] ,
         \mult_22/SUMB[27][61] , \mult_22/SUMB[27][62] , \mult_22/SUMB[28][1] ,
         \mult_22/SUMB[28][2] , \mult_22/SUMB[28][3] , \mult_22/SUMB[28][4] ,
         \mult_22/SUMB[28][5] , \mult_22/SUMB[28][6] , \mult_22/SUMB[28][7] ,
         \mult_22/SUMB[28][8] , \mult_22/SUMB[28][9] , \mult_22/SUMB[28][10] ,
         \mult_22/SUMB[28][11] , \mult_22/SUMB[28][12] ,
         \mult_22/SUMB[28][13] , \mult_22/SUMB[28][14] ,
         \mult_22/SUMB[28][15] , \mult_22/SUMB[28][16] ,
         \mult_22/SUMB[28][17] , \mult_22/SUMB[28][18] ,
         \mult_22/SUMB[28][19] , \mult_22/SUMB[28][20] ,
         \mult_22/SUMB[28][21] , \mult_22/SUMB[28][22] ,
         \mult_22/SUMB[28][23] , \mult_22/SUMB[28][24] ,
         \mult_22/SUMB[28][25] , \mult_22/SUMB[28][26] ,
         \mult_22/SUMB[28][27] , \mult_22/SUMB[28][28] ,
         \mult_22/SUMB[28][29] , \mult_22/SUMB[28][30] ,
         \mult_22/SUMB[28][31] , \mult_22/SUMB[28][32] ,
         \mult_22/SUMB[28][33] , \mult_22/SUMB[28][34] ,
         \mult_22/SUMB[28][35] , \mult_22/SUMB[28][36] ,
         \mult_22/SUMB[28][37] , \mult_22/SUMB[28][38] ,
         \mult_22/SUMB[28][39] , \mult_22/SUMB[28][40] ,
         \mult_22/SUMB[28][41] , \mult_22/SUMB[28][42] ,
         \mult_22/SUMB[28][43] , \mult_22/SUMB[28][44] ,
         \mult_22/SUMB[28][45] , \mult_22/SUMB[28][46] ,
         \mult_22/SUMB[28][47] , \mult_22/SUMB[28][48] ,
         \mult_22/SUMB[28][49] , \mult_22/SUMB[28][50] ,
         \mult_22/SUMB[28][51] , \mult_22/SUMB[28][52] ,
         \mult_22/SUMB[28][53] , \mult_22/SUMB[28][54] ,
         \mult_22/SUMB[28][55] , \mult_22/SUMB[28][56] ,
         \mult_22/SUMB[28][57] , \mult_22/SUMB[28][58] ,
         \mult_22/SUMB[28][59] , \mult_22/SUMB[28][60] ,
         \mult_22/SUMB[28][61] , \mult_22/SUMB[28][62] , \mult_22/SUMB[29][1] ,
         \mult_22/SUMB[29][2] , \mult_22/SUMB[29][3] , \mult_22/SUMB[29][4] ,
         \mult_22/SUMB[29][5] , \mult_22/SUMB[29][6] , \mult_22/SUMB[29][7] ,
         \mult_22/SUMB[29][8] , \mult_22/SUMB[29][9] , \mult_22/SUMB[29][10] ,
         \mult_22/SUMB[29][11] , \mult_22/SUMB[29][12] ,
         \mult_22/SUMB[29][13] , \mult_22/SUMB[29][14] ,
         \mult_22/SUMB[29][15] , \mult_22/SUMB[29][16] ,
         \mult_22/SUMB[29][17] , \mult_22/SUMB[29][18] ,
         \mult_22/SUMB[29][19] , \mult_22/SUMB[29][20] ,
         \mult_22/SUMB[29][21] , \mult_22/SUMB[29][22] ,
         \mult_22/SUMB[29][23] , \mult_22/SUMB[29][24] ,
         \mult_22/SUMB[29][25] , \mult_22/SUMB[29][26] ,
         \mult_22/SUMB[29][27] , \mult_22/SUMB[29][28] ,
         \mult_22/SUMB[29][29] , \mult_22/SUMB[29][30] ,
         \mult_22/SUMB[29][31] , \mult_22/SUMB[29][32] ,
         \mult_22/SUMB[29][33] , \mult_22/SUMB[29][34] ,
         \mult_22/SUMB[29][35] , \mult_22/SUMB[29][36] ,
         \mult_22/SUMB[29][37] , \mult_22/SUMB[29][38] ,
         \mult_22/SUMB[29][39] , \mult_22/SUMB[29][40] ,
         \mult_22/SUMB[29][41] , \mult_22/SUMB[29][42] ,
         \mult_22/SUMB[29][43] , \mult_22/SUMB[29][44] ,
         \mult_22/SUMB[29][45] , \mult_22/SUMB[29][46] ,
         \mult_22/SUMB[29][47] , \mult_22/SUMB[29][48] ,
         \mult_22/SUMB[29][49] , \mult_22/SUMB[29][50] ,
         \mult_22/SUMB[29][51] , \mult_22/SUMB[29][52] ,
         \mult_22/SUMB[29][53] , \mult_22/SUMB[29][54] ,
         \mult_22/SUMB[29][55] , \mult_22/SUMB[29][56] ,
         \mult_22/SUMB[29][57] , \mult_22/SUMB[29][58] ,
         \mult_22/SUMB[29][59] , \mult_22/SUMB[29][60] ,
         \mult_22/SUMB[29][61] , \mult_22/SUMB[29][62] , \mult_22/SUMB[30][1] ,
         \mult_22/SUMB[30][2] , \mult_22/SUMB[30][3] , \mult_22/SUMB[30][4] ,
         \mult_22/SUMB[30][5] , \mult_22/SUMB[30][6] , \mult_22/SUMB[30][7] ,
         \mult_22/SUMB[30][8] , \mult_22/SUMB[30][9] , \mult_22/SUMB[30][10] ,
         \mult_22/SUMB[30][11] , \mult_22/SUMB[30][12] ,
         \mult_22/SUMB[30][13] , \mult_22/SUMB[30][14] ,
         \mult_22/SUMB[30][15] , \mult_22/SUMB[30][16] ,
         \mult_22/SUMB[30][17] , \mult_22/SUMB[30][18] ,
         \mult_22/SUMB[30][19] , \mult_22/SUMB[30][20] ,
         \mult_22/SUMB[30][21] , \mult_22/SUMB[30][22] ,
         \mult_22/SUMB[30][23] , \mult_22/SUMB[30][24] ,
         \mult_22/SUMB[30][25] , \mult_22/SUMB[30][26] ,
         \mult_22/SUMB[30][27] , \mult_22/SUMB[30][28] ,
         \mult_22/SUMB[30][29] , \mult_22/SUMB[30][30] ,
         \mult_22/SUMB[30][31] , \mult_22/SUMB[30][32] ,
         \mult_22/SUMB[30][33] , \mult_22/SUMB[30][34] ,
         \mult_22/SUMB[30][35] , \mult_22/SUMB[30][36] ,
         \mult_22/SUMB[30][37] , \mult_22/SUMB[30][38] ,
         \mult_22/SUMB[30][39] , \mult_22/SUMB[30][40] ,
         \mult_22/SUMB[30][41] , \mult_22/SUMB[30][42] ,
         \mult_22/SUMB[30][43] , \mult_22/SUMB[30][44] ,
         \mult_22/SUMB[30][45] , \mult_22/SUMB[30][46] ,
         \mult_22/SUMB[30][47] , \mult_22/SUMB[30][48] ,
         \mult_22/SUMB[30][49] , \mult_22/SUMB[30][50] ,
         \mult_22/SUMB[30][51] , \mult_22/SUMB[30][52] ,
         \mult_22/SUMB[30][53] , \mult_22/SUMB[30][54] ,
         \mult_22/SUMB[30][55] , \mult_22/SUMB[30][56] ,
         \mult_22/SUMB[30][57] , \mult_22/SUMB[30][58] ,
         \mult_22/SUMB[30][59] , \mult_22/SUMB[30][60] ,
         \mult_22/SUMB[30][61] , \mult_22/SUMB[30][62] , \mult_22/SUMB[31][1] ,
         \mult_22/SUMB[31][2] , \mult_22/SUMB[31][3] , \mult_22/SUMB[31][4] ,
         \mult_22/SUMB[31][5] , \mult_22/SUMB[31][6] , \mult_22/SUMB[31][7] ,
         \mult_22/SUMB[31][8] , \mult_22/SUMB[31][9] , \mult_22/SUMB[31][10] ,
         \mult_22/SUMB[31][11] , \mult_22/SUMB[31][12] ,
         \mult_22/SUMB[31][13] , \mult_22/SUMB[31][14] ,
         \mult_22/SUMB[31][15] , \mult_22/SUMB[31][16] ,
         \mult_22/SUMB[31][17] , \mult_22/SUMB[31][18] ,
         \mult_22/SUMB[31][19] , \mult_22/SUMB[31][20] ,
         \mult_22/SUMB[31][21] , \mult_22/SUMB[31][22] ,
         \mult_22/SUMB[31][23] , \mult_22/SUMB[31][24] ,
         \mult_22/SUMB[31][25] , \mult_22/SUMB[31][26] ,
         \mult_22/SUMB[31][27] , \mult_22/SUMB[31][28] ,
         \mult_22/SUMB[31][29] , \mult_22/SUMB[31][30] ,
         \mult_22/SUMB[31][31] , \mult_22/SUMB[31][32] ,
         \mult_22/SUMB[31][33] , \mult_22/SUMB[31][34] ,
         \mult_22/SUMB[31][35] , \mult_22/SUMB[31][36] ,
         \mult_22/SUMB[31][37] , \mult_22/SUMB[31][38] ,
         \mult_22/SUMB[31][39] , \mult_22/SUMB[31][40] ,
         \mult_22/SUMB[31][41] , \mult_22/SUMB[31][42] ,
         \mult_22/SUMB[31][43] , \mult_22/SUMB[31][44] ,
         \mult_22/SUMB[31][45] , \mult_22/SUMB[31][46] ,
         \mult_22/SUMB[31][47] , \mult_22/SUMB[31][48] ,
         \mult_22/SUMB[31][49] , \mult_22/SUMB[31][50] ,
         \mult_22/SUMB[31][51] , \mult_22/SUMB[31][52] ,
         \mult_22/SUMB[31][53] , \mult_22/SUMB[31][54] ,
         \mult_22/SUMB[31][55] , \mult_22/SUMB[31][56] ,
         \mult_22/SUMB[31][57] , \mult_22/SUMB[31][58] ,
         \mult_22/SUMB[31][59] , \mult_22/SUMB[31][60] ,
         \mult_22/SUMB[31][61] , \mult_22/SUMB[31][62] ,
         \mult_22/CARRYB[24][0] , \mult_22/CARRYB[24][1] ,
         \mult_22/CARRYB[24][2] , \mult_22/CARRYB[24][3] ,
         \mult_22/CARRYB[24][4] , \mult_22/CARRYB[24][5] ,
         \mult_22/CARRYB[24][6] , \mult_22/CARRYB[24][7] ,
         \mult_22/CARRYB[24][8] , \mult_22/CARRYB[24][9] ,
         \mult_22/CARRYB[24][10] , \mult_22/CARRYB[24][11] ,
         \mult_22/CARRYB[24][12] , \mult_22/CARRYB[24][13] ,
         \mult_22/CARRYB[24][14] , \mult_22/CARRYB[24][15] ,
         \mult_22/CARRYB[24][16] , \mult_22/CARRYB[24][17] ,
         \mult_22/CARRYB[24][18] , \mult_22/CARRYB[24][19] ,
         \mult_22/CARRYB[24][20] , \mult_22/CARRYB[24][21] ,
         \mult_22/CARRYB[24][22] , \mult_22/CARRYB[24][23] ,
         \mult_22/CARRYB[24][24] , \mult_22/CARRYB[24][25] ,
         \mult_22/CARRYB[24][26] , \mult_22/CARRYB[24][27] ,
         \mult_22/CARRYB[24][28] , \mult_22/CARRYB[24][29] ,
         \mult_22/CARRYB[24][30] , \mult_22/CARRYB[24][31] ,
         \mult_22/CARRYB[24][32] , \mult_22/CARRYB[24][33] ,
         \mult_22/CARRYB[24][34] , \mult_22/CARRYB[24][35] ,
         \mult_22/CARRYB[24][36] , \mult_22/CARRYB[24][37] ,
         \mult_22/CARRYB[24][38] , \mult_22/CARRYB[24][39] ,
         \mult_22/CARRYB[24][40] , \mult_22/CARRYB[24][41] ,
         \mult_22/CARRYB[24][42] , \mult_22/CARRYB[24][43] ,
         \mult_22/CARRYB[24][44] , \mult_22/CARRYB[24][45] ,
         \mult_22/CARRYB[24][46] , \mult_22/CARRYB[24][47] ,
         \mult_22/CARRYB[24][48] , \mult_22/CARRYB[24][49] ,
         \mult_22/CARRYB[24][50] , \mult_22/CARRYB[24][51] ,
         \mult_22/CARRYB[24][52] , \mult_22/CARRYB[24][53] ,
         \mult_22/CARRYB[24][54] , \mult_22/CARRYB[24][55] ,
         \mult_22/CARRYB[24][56] , \mult_22/CARRYB[24][57] ,
         \mult_22/CARRYB[24][58] , \mult_22/CARRYB[24][59] ,
         \mult_22/CARRYB[24][60] , \mult_22/CARRYB[24][61] ,
         \mult_22/CARRYB[24][62] , \mult_22/CARRYB[25][0] ,
         \mult_22/CARRYB[25][1] , \mult_22/CARRYB[25][2] ,
         \mult_22/CARRYB[25][3] , \mult_22/CARRYB[25][4] ,
         \mult_22/CARRYB[25][5] , \mult_22/CARRYB[25][6] ,
         \mult_22/CARRYB[25][7] , \mult_22/CARRYB[25][8] ,
         \mult_22/CARRYB[25][9] , \mult_22/CARRYB[25][10] ,
         \mult_22/CARRYB[25][11] , \mult_22/CARRYB[25][12] ,
         \mult_22/CARRYB[25][13] , \mult_22/CARRYB[25][14] ,
         \mult_22/CARRYB[25][15] , \mult_22/CARRYB[25][16] ,
         \mult_22/CARRYB[25][17] , \mult_22/CARRYB[25][18] ,
         \mult_22/CARRYB[25][19] , \mult_22/CARRYB[25][20] ,
         \mult_22/CARRYB[25][21] , \mult_22/CARRYB[25][22] ,
         \mult_22/CARRYB[25][23] , \mult_22/CARRYB[25][24] ,
         \mult_22/CARRYB[25][25] , \mult_22/CARRYB[25][26] ,
         \mult_22/CARRYB[25][27] , \mult_22/CARRYB[25][28] ,
         \mult_22/CARRYB[25][29] , \mult_22/CARRYB[25][30] ,
         \mult_22/CARRYB[25][31] , \mult_22/CARRYB[25][32] ,
         \mult_22/CARRYB[25][33] , \mult_22/CARRYB[25][34] ,
         \mult_22/CARRYB[25][35] , \mult_22/CARRYB[25][36] ,
         \mult_22/CARRYB[25][37] , \mult_22/CARRYB[25][38] ,
         \mult_22/CARRYB[25][39] , \mult_22/CARRYB[25][40] ,
         \mult_22/CARRYB[25][41] , \mult_22/CARRYB[25][42] ,
         \mult_22/CARRYB[25][43] , \mult_22/CARRYB[25][44] ,
         \mult_22/CARRYB[25][45] , \mult_22/CARRYB[25][46] ,
         \mult_22/CARRYB[25][47] , \mult_22/CARRYB[25][48] ,
         \mult_22/CARRYB[25][49] , \mult_22/CARRYB[25][50] ,
         \mult_22/CARRYB[25][51] , \mult_22/CARRYB[25][52] ,
         \mult_22/CARRYB[25][53] , \mult_22/CARRYB[25][54] ,
         \mult_22/CARRYB[25][55] , \mult_22/CARRYB[25][56] ,
         \mult_22/CARRYB[25][57] , \mult_22/CARRYB[25][58] ,
         \mult_22/CARRYB[25][59] , \mult_22/CARRYB[25][60] ,
         \mult_22/CARRYB[25][61] , \mult_22/CARRYB[25][62] ,
         \mult_22/CARRYB[26][0] , \mult_22/CARRYB[26][1] ,
         \mult_22/CARRYB[26][2] , \mult_22/CARRYB[26][3] ,
         \mult_22/CARRYB[26][4] , \mult_22/CARRYB[26][5] ,
         \mult_22/CARRYB[26][6] , \mult_22/CARRYB[26][7] ,
         \mult_22/CARRYB[26][8] , \mult_22/CARRYB[26][9] ,
         \mult_22/CARRYB[26][10] , \mult_22/CARRYB[26][11] ,
         \mult_22/CARRYB[26][12] , \mult_22/CARRYB[26][13] ,
         \mult_22/CARRYB[26][14] , \mult_22/CARRYB[26][15] ,
         \mult_22/CARRYB[26][16] , \mult_22/CARRYB[26][17] ,
         \mult_22/CARRYB[26][18] , \mult_22/CARRYB[26][19] ,
         \mult_22/CARRYB[26][20] , \mult_22/CARRYB[26][21] ,
         \mult_22/CARRYB[26][22] , \mult_22/CARRYB[26][23] ,
         \mult_22/CARRYB[26][24] , \mult_22/CARRYB[26][25] ,
         \mult_22/CARRYB[26][26] , \mult_22/CARRYB[26][27] ,
         \mult_22/CARRYB[26][28] , \mult_22/CARRYB[26][29] ,
         \mult_22/CARRYB[26][30] , \mult_22/CARRYB[26][31] ,
         \mult_22/CARRYB[26][32] , \mult_22/CARRYB[26][33] ,
         \mult_22/CARRYB[26][34] , \mult_22/CARRYB[26][35] ,
         \mult_22/CARRYB[26][36] , \mult_22/CARRYB[26][37] ,
         \mult_22/CARRYB[26][38] , \mult_22/CARRYB[26][39] ,
         \mult_22/CARRYB[26][40] , \mult_22/CARRYB[26][41] ,
         \mult_22/CARRYB[26][42] , \mult_22/CARRYB[26][43] ,
         \mult_22/CARRYB[26][44] , \mult_22/CARRYB[26][45] ,
         \mult_22/CARRYB[26][46] , \mult_22/CARRYB[26][47] ,
         \mult_22/CARRYB[26][48] , \mult_22/CARRYB[26][49] ,
         \mult_22/CARRYB[26][50] , \mult_22/CARRYB[26][51] ,
         \mult_22/CARRYB[26][52] , \mult_22/CARRYB[26][53] ,
         \mult_22/CARRYB[26][54] , \mult_22/CARRYB[26][55] ,
         \mult_22/CARRYB[26][56] , \mult_22/CARRYB[26][57] ,
         \mult_22/CARRYB[26][58] , \mult_22/CARRYB[26][59] ,
         \mult_22/CARRYB[26][60] , \mult_22/CARRYB[26][61] ,
         \mult_22/CARRYB[26][62] , \mult_22/CARRYB[27][0] ,
         \mult_22/CARRYB[27][1] , \mult_22/CARRYB[27][2] ,
         \mult_22/CARRYB[27][3] , \mult_22/CARRYB[27][4] ,
         \mult_22/CARRYB[27][5] , \mult_22/CARRYB[27][6] ,
         \mult_22/CARRYB[27][7] , \mult_22/CARRYB[27][8] ,
         \mult_22/CARRYB[27][9] , \mult_22/CARRYB[27][10] ,
         \mult_22/CARRYB[27][11] , \mult_22/CARRYB[27][12] ,
         \mult_22/CARRYB[27][13] , \mult_22/CARRYB[27][14] ,
         \mult_22/CARRYB[27][15] , \mult_22/CARRYB[27][16] ,
         \mult_22/CARRYB[27][17] , \mult_22/CARRYB[27][18] ,
         \mult_22/CARRYB[27][19] , \mult_22/CARRYB[27][20] ,
         \mult_22/CARRYB[27][21] , \mult_22/CARRYB[27][22] ,
         \mult_22/CARRYB[27][23] , \mult_22/CARRYB[27][24] ,
         \mult_22/CARRYB[27][25] , \mult_22/CARRYB[27][26] ,
         \mult_22/CARRYB[27][27] , \mult_22/CARRYB[27][28] ,
         \mult_22/CARRYB[27][29] , \mult_22/CARRYB[27][30] ,
         \mult_22/CARRYB[27][31] , \mult_22/CARRYB[27][32] ,
         \mult_22/CARRYB[27][33] , \mult_22/CARRYB[27][34] ,
         \mult_22/CARRYB[27][35] , \mult_22/CARRYB[27][36] ,
         \mult_22/CARRYB[27][37] , \mult_22/CARRYB[27][38] ,
         \mult_22/CARRYB[27][39] , \mult_22/CARRYB[27][40] ,
         \mult_22/CARRYB[27][41] , \mult_22/CARRYB[27][42] ,
         \mult_22/CARRYB[27][43] , \mult_22/CARRYB[27][44] ,
         \mult_22/CARRYB[27][45] , \mult_22/CARRYB[27][46] ,
         \mult_22/CARRYB[27][47] , \mult_22/CARRYB[27][48] ,
         \mult_22/CARRYB[27][49] , \mult_22/CARRYB[27][50] ,
         \mult_22/CARRYB[27][51] , \mult_22/CARRYB[27][52] ,
         \mult_22/CARRYB[27][53] , \mult_22/CARRYB[27][54] ,
         \mult_22/CARRYB[27][55] , \mult_22/CARRYB[27][56] ,
         \mult_22/CARRYB[27][57] , \mult_22/CARRYB[27][58] ,
         \mult_22/CARRYB[27][59] , \mult_22/CARRYB[27][60] ,
         \mult_22/CARRYB[27][61] , \mult_22/CARRYB[27][62] ,
         \mult_22/CARRYB[28][0] , \mult_22/CARRYB[28][1] ,
         \mult_22/CARRYB[28][2] , \mult_22/CARRYB[28][3] ,
         \mult_22/CARRYB[28][4] , \mult_22/CARRYB[28][5] ,
         \mult_22/CARRYB[28][6] , \mult_22/CARRYB[28][7] ,
         \mult_22/CARRYB[28][8] , \mult_22/CARRYB[28][9] ,
         \mult_22/CARRYB[28][10] , \mult_22/CARRYB[28][11] ,
         \mult_22/CARRYB[28][12] , \mult_22/CARRYB[28][13] ,
         \mult_22/CARRYB[28][14] , \mult_22/CARRYB[28][15] ,
         \mult_22/CARRYB[28][16] , \mult_22/CARRYB[28][17] ,
         \mult_22/CARRYB[28][18] , \mult_22/CARRYB[28][19] ,
         \mult_22/CARRYB[28][20] , \mult_22/CARRYB[28][21] ,
         \mult_22/CARRYB[28][22] , \mult_22/CARRYB[28][23] ,
         \mult_22/CARRYB[28][24] , \mult_22/CARRYB[28][25] ,
         \mult_22/CARRYB[28][26] , \mult_22/CARRYB[28][27] ,
         \mult_22/CARRYB[28][28] , \mult_22/CARRYB[28][29] ,
         \mult_22/CARRYB[28][30] , \mult_22/CARRYB[28][31] ,
         \mult_22/CARRYB[28][32] , \mult_22/CARRYB[28][33] ,
         \mult_22/CARRYB[28][34] , \mult_22/CARRYB[28][35] ,
         \mult_22/CARRYB[28][36] , \mult_22/CARRYB[28][37] ,
         \mult_22/CARRYB[28][38] , \mult_22/CARRYB[28][39] ,
         \mult_22/CARRYB[28][40] , \mult_22/CARRYB[28][41] ,
         \mult_22/CARRYB[28][42] , \mult_22/CARRYB[28][43] ,
         \mult_22/CARRYB[28][44] , \mult_22/CARRYB[28][45] ,
         \mult_22/CARRYB[28][46] , \mult_22/CARRYB[28][47] ,
         \mult_22/CARRYB[28][48] , \mult_22/CARRYB[28][49] ,
         \mult_22/CARRYB[28][50] , \mult_22/CARRYB[28][51] ,
         \mult_22/CARRYB[28][52] , \mult_22/CARRYB[28][53] ,
         \mult_22/CARRYB[28][54] , \mult_22/CARRYB[28][55] ,
         \mult_22/CARRYB[28][56] , \mult_22/CARRYB[28][57] ,
         \mult_22/CARRYB[28][58] , \mult_22/CARRYB[28][59] ,
         \mult_22/CARRYB[28][60] , \mult_22/CARRYB[28][61] ,
         \mult_22/CARRYB[28][62] , \mult_22/CARRYB[29][0] ,
         \mult_22/CARRYB[29][1] , \mult_22/CARRYB[29][2] ,
         \mult_22/CARRYB[29][3] , \mult_22/CARRYB[29][4] ,
         \mult_22/CARRYB[29][5] , \mult_22/CARRYB[29][6] ,
         \mult_22/CARRYB[29][7] , \mult_22/CARRYB[29][8] ,
         \mult_22/CARRYB[29][9] , \mult_22/CARRYB[29][10] ,
         \mult_22/CARRYB[29][11] , \mult_22/CARRYB[29][12] ,
         \mult_22/CARRYB[29][13] , \mult_22/CARRYB[29][14] ,
         \mult_22/CARRYB[29][15] , \mult_22/CARRYB[29][16] ,
         \mult_22/CARRYB[29][17] , \mult_22/CARRYB[29][18] ,
         \mult_22/CARRYB[29][19] , \mult_22/CARRYB[29][20] ,
         \mult_22/CARRYB[29][21] , \mult_22/CARRYB[29][22] ,
         \mult_22/CARRYB[29][23] , \mult_22/CARRYB[29][24] ,
         \mult_22/CARRYB[29][25] , \mult_22/CARRYB[29][26] ,
         \mult_22/CARRYB[29][27] , \mult_22/CARRYB[29][28] ,
         \mult_22/CARRYB[29][29] , \mult_22/CARRYB[29][30] ,
         \mult_22/CARRYB[29][31] , \mult_22/CARRYB[29][32] ,
         \mult_22/CARRYB[29][33] , \mult_22/CARRYB[29][34] ,
         \mult_22/CARRYB[29][35] , \mult_22/CARRYB[29][36] ,
         \mult_22/CARRYB[29][37] , \mult_22/CARRYB[29][38] ,
         \mult_22/CARRYB[29][39] , \mult_22/CARRYB[29][40] ,
         \mult_22/CARRYB[29][41] , \mult_22/CARRYB[29][42] ,
         \mult_22/CARRYB[29][43] , \mult_22/CARRYB[29][44] ,
         \mult_22/CARRYB[29][45] , \mult_22/CARRYB[29][46] ,
         \mult_22/CARRYB[29][47] , \mult_22/CARRYB[29][48] ,
         \mult_22/CARRYB[29][49] , \mult_22/CARRYB[29][50] ,
         \mult_22/CARRYB[29][51] , \mult_22/CARRYB[29][52] ,
         \mult_22/CARRYB[29][53] , \mult_22/CARRYB[29][54] ,
         \mult_22/CARRYB[29][55] , \mult_22/CARRYB[29][56] ,
         \mult_22/CARRYB[29][57] , \mult_22/CARRYB[29][58] ,
         \mult_22/CARRYB[29][59] , \mult_22/CARRYB[29][60] ,
         \mult_22/CARRYB[29][61] , \mult_22/CARRYB[29][62] ,
         \mult_22/CARRYB[30][0] , \mult_22/CARRYB[30][1] ,
         \mult_22/CARRYB[30][2] , \mult_22/CARRYB[30][3] ,
         \mult_22/CARRYB[30][4] , \mult_22/CARRYB[30][5] ,
         \mult_22/CARRYB[30][6] , \mult_22/CARRYB[30][7] ,
         \mult_22/CARRYB[30][8] , \mult_22/CARRYB[30][9] ,
         \mult_22/CARRYB[30][10] , \mult_22/CARRYB[30][11] ,
         \mult_22/CARRYB[30][12] , \mult_22/CARRYB[30][13] ,
         \mult_22/CARRYB[30][14] , \mult_22/CARRYB[30][15] ,
         \mult_22/CARRYB[30][16] , \mult_22/CARRYB[30][17] ,
         \mult_22/CARRYB[30][18] , \mult_22/CARRYB[30][19] ,
         \mult_22/CARRYB[30][20] , \mult_22/CARRYB[30][21] ,
         \mult_22/CARRYB[30][22] , \mult_22/CARRYB[30][23] ,
         \mult_22/CARRYB[30][24] , \mult_22/CARRYB[30][25] ,
         \mult_22/CARRYB[30][26] , \mult_22/CARRYB[30][27] ,
         \mult_22/CARRYB[30][28] , \mult_22/CARRYB[30][29] ,
         \mult_22/CARRYB[30][30] , \mult_22/CARRYB[30][31] ,
         \mult_22/CARRYB[30][32] , \mult_22/CARRYB[30][33] ,
         \mult_22/CARRYB[30][34] , \mult_22/CARRYB[30][35] ,
         \mult_22/CARRYB[30][36] , \mult_22/CARRYB[30][37] ,
         \mult_22/CARRYB[30][38] , \mult_22/CARRYB[30][39] ,
         \mult_22/CARRYB[30][40] , \mult_22/CARRYB[30][41] ,
         \mult_22/CARRYB[30][42] , \mult_22/CARRYB[30][43] ,
         \mult_22/CARRYB[30][44] , \mult_22/CARRYB[30][45] ,
         \mult_22/CARRYB[30][46] , \mult_22/CARRYB[30][47] ,
         \mult_22/CARRYB[30][48] , \mult_22/CARRYB[30][49] ,
         \mult_22/CARRYB[30][50] , \mult_22/CARRYB[30][51] ,
         \mult_22/CARRYB[30][52] , \mult_22/CARRYB[30][53] ,
         \mult_22/CARRYB[30][54] , \mult_22/CARRYB[30][55] ,
         \mult_22/CARRYB[30][56] , \mult_22/CARRYB[30][57] ,
         \mult_22/CARRYB[30][58] , \mult_22/CARRYB[30][59] ,
         \mult_22/CARRYB[30][60] , \mult_22/CARRYB[30][61] ,
         \mult_22/CARRYB[30][62] , \mult_22/CARRYB[31][0] ,
         \mult_22/CARRYB[31][1] , \mult_22/CARRYB[31][2] ,
         \mult_22/CARRYB[31][3] , \mult_22/CARRYB[31][4] ,
         \mult_22/CARRYB[31][5] , \mult_22/CARRYB[31][6] ,
         \mult_22/CARRYB[31][7] , \mult_22/CARRYB[31][8] ,
         \mult_22/CARRYB[31][9] , \mult_22/CARRYB[31][10] ,
         \mult_22/CARRYB[31][11] , \mult_22/CARRYB[31][12] ,
         \mult_22/CARRYB[31][13] , \mult_22/CARRYB[31][14] ,
         \mult_22/CARRYB[31][15] , \mult_22/CARRYB[31][16] ,
         \mult_22/CARRYB[31][17] , \mult_22/CARRYB[31][18] ,
         \mult_22/CARRYB[31][19] , \mult_22/CARRYB[31][20] ,
         \mult_22/CARRYB[31][21] , \mult_22/CARRYB[31][22] ,
         \mult_22/CARRYB[31][23] , \mult_22/CARRYB[31][24] ,
         \mult_22/CARRYB[31][25] , \mult_22/CARRYB[31][26] ,
         \mult_22/CARRYB[31][27] , \mult_22/CARRYB[31][28] ,
         \mult_22/CARRYB[31][29] , \mult_22/CARRYB[31][30] ,
         \mult_22/CARRYB[31][31] , \mult_22/CARRYB[31][32] ,
         \mult_22/CARRYB[31][33] , \mult_22/CARRYB[31][34] ,
         \mult_22/CARRYB[31][35] , \mult_22/CARRYB[31][36] ,
         \mult_22/CARRYB[31][37] , \mult_22/CARRYB[31][38] ,
         \mult_22/CARRYB[31][39] , \mult_22/CARRYB[31][40] ,
         \mult_22/CARRYB[31][41] , \mult_22/CARRYB[31][42] ,
         \mult_22/CARRYB[31][43] , \mult_22/CARRYB[31][44] ,
         \mult_22/CARRYB[31][45] , \mult_22/CARRYB[31][46] ,
         \mult_22/CARRYB[31][47] , \mult_22/CARRYB[31][48] ,
         \mult_22/CARRYB[31][49] , \mult_22/CARRYB[31][50] ,
         \mult_22/CARRYB[31][51] , \mult_22/CARRYB[31][52] ,
         \mult_22/CARRYB[31][53] , \mult_22/CARRYB[31][54] ,
         \mult_22/CARRYB[31][55] , \mult_22/CARRYB[31][56] ,
         \mult_22/CARRYB[31][57] , \mult_22/CARRYB[31][58] ,
         \mult_22/CARRYB[31][59] , \mult_22/CARRYB[31][60] ,
         \mult_22/CARRYB[31][61] , \mult_22/CARRYB[31][62] ,
         \mult_22/SUMB[16][1] , \mult_22/SUMB[16][2] , \mult_22/SUMB[16][3] ,
         \mult_22/SUMB[16][4] , \mult_22/SUMB[16][5] , \mult_22/SUMB[16][6] ,
         \mult_22/SUMB[16][7] , \mult_22/SUMB[16][8] , \mult_22/SUMB[16][9] ,
         \mult_22/SUMB[16][10] , \mult_22/SUMB[16][11] ,
         \mult_22/SUMB[16][12] , \mult_22/SUMB[16][13] ,
         \mult_22/SUMB[16][14] , \mult_22/SUMB[16][15] ,
         \mult_22/SUMB[16][16] , \mult_22/SUMB[16][17] ,
         \mult_22/SUMB[16][18] , \mult_22/SUMB[16][19] ,
         \mult_22/SUMB[16][20] , \mult_22/SUMB[16][21] ,
         \mult_22/SUMB[16][22] , \mult_22/SUMB[16][23] ,
         \mult_22/SUMB[16][24] , \mult_22/SUMB[16][25] ,
         \mult_22/SUMB[16][26] , \mult_22/SUMB[16][27] ,
         \mult_22/SUMB[16][28] , \mult_22/SUMB[16][29] ,
         \mult_22/SUMB[16][30] , \mult_22/SUMB[16][31] ,
         \mult_22/SUMB[16][32] , \mult_22/SUMB[16][33] ,
         \mult_22/SUMB[16][34] , \mult_22/SUMB[16][35] ,
         \mult_22/SUMB[16][36] , \mult_22/SUMB[16][37] ,
         \mult_22/SUMB[16][38] , \mult_22/SUMB[16][39] ,
         \mult_22/SUMB[16][40] , \mult_22/SUMB[16][41] ,
         \mult_22/SUMB[16][42] , \mult_22/SUMB[16][43] ,
         \mult_22/SUMB[16][44] , \mult_22/SUMB[16][45] ,
         \mult_22/SUMB[16][46] , \mult_22/SUMB[16][47] ,
         \mult_22/SUMB[16][48] , \mult_22/SUMB[16][49] ,
         \mult_22/SUMB[16][50] , \mult_22/SUMB[16][51] ,
         \mult_22/SUMB[16][52] , \mult_22/SUMB[16][53] ,
         \mult_22/SUMB[16][54] , \mult_22/SUMB[16][55] ,
         \mult_22/SUMB[16][56] , \mult_22/SUMB[16][57] ,
         \mult_22/SUMB[16][58] , \mult_22/SUMB[16][59] ,
         \mult_22/SUMB[16][60] , \mult_22/SUMB[16][61] ,
         \mult_22/SUMB[16][62] , \mult_22/SUMB[17][1] , \mult_22/SUMB[17][2] ,
         \mult_22/SUMB[17][3] , \mult_22/SUMB[17][4] , \mult_22/SUMB[17][5] ,
         \mult_22/SUMB[17][6] , \mult_22/SUMB[17][7] , \mult_22/SUMB[17][8] ,
         \mult_22/SUMB[17][9] , \mult_22/SUMB[17][10] , \mult_22/SUMB[17][11] ,
         \mult_22/SUMB[17][12] , \mult_22/SUMB[17][13] ,
         \mult_22/SUMB[17][14] , \mult_22/SUMB[17][15] ,
         \mult_22/SUMB[17][16] , \mult_22/SUMB[17][17] ,
         \mult_22/SUMB[17][18] , \mult_22/SUMB[17][19] ,
         \mult_22/SUMB[17][20] , \mult_22/SUMB[17][21] ,
         \mult_22/SUMB[17][22] , \mult_22/SUMB[17][23] ,
         \mult_22/SUMB[17][24] , \mult_22/SUMB[17][25] ,
         \mult_22/SUMB[17][26] , \mult_22/SUMB[17][27] ,
         \mult_22/SUMB[17][28] , \mult_22/SUMB[17][29] ,
         \mult_22/SUMB[17][30] , \mult_22/SUMB[17][31] ,
         \mult_22/SUMB[17][32] , \mult_22/SUMB[17][33] ,
         \mult_22/SUMB[17][34] , \mult_22/SUMB[17][35] ,
         \mult_22/SUMB[17][36] , \mult_22/SUMB[17][37] ,
         \mult_22/SUMB[17][38] , \mult_22/SUMB[17][39] ,
         \mult_22/SUMB[17][40] , \mult_22/SUMB[17][41] ,
         \mult_22/SUMB[17][42] , \mult_22/SUMB[17][43] ,
         \mult_22/SUMB[17][44] , \mult_22/SUMB[17][45] ,
         \mult_22/SUMB[17][46] , \mult_22/SUMB[17][47] ,
         \mult_22/SUMB[17][48] , \mult_22/SUMB[17][49] ,
         \mult_22/SUMB[17][50] , \mult_22/SUMB[17][51] ,
         \mult_22/SUMB[17][52] , \mult_22/SUMB[17][53] ,
         \mult_22/SUMB[17][54] , \mult_22/SUMB[17][55] ,
         \mult_22/SUMB[17][56] , \mult_22/SUMB[17][57] ,
         \mult_22/SUMB[17][58] , \mult_22/SUMB[17][59] ,
         \mult_22/SUMB[17][60] , \mult_22/SUMB[17][61] ,
         \mult_22/SUMB[17][62] , \mult_22/SUMB[18][1] , \mult_22/SUMB[18][2] ,
         \mult_22/SUMB[18][3] , \mult_22/SUMB[18][4] , \mult_22/SUMB[18][5] ,
         \mult_22/SUMB[18][6] , \mult_22/SUMB[18][7] , \mult_22/SUMB[18][8] ,
         \mult_22/SUMB[18][9] , \mult_22/SUMB[18][10] , \mult_22/SUMB[18][11] ,
         \mult_22/SUMB[18][12] , \mult_22/SUMB[18][13] ,
         \mult_22/SUMB[18][14] , \mult_22/SUMB[18][15] ,
         \mult_22/SUMB[18][16] , \mult_22/SUMB[18][17] ,
         \mult_22/SUMB[18][18] , \mult_22/SUMB[18][19] ,
         \mult_22/SUMB[18][20] , \mult_22/SUMB[18][21] ,
         \mult_22/SUMB[18][22] , \mult_22/SUMB[18][23] ,
         \mult_22/SUMB[18][24] , \mult_22/SUMB[18][25] ,
         \mult_22/SUMB[18][26] , \mult_22/SUMB[18][27] ,
         \mult_22/SUMB[18][28] , \mult_22/SUMB[18][29] ,
         \mult_22/SUMB[18][30] , \mult_22/SUMB[18][31] ,
         \mult_22/SUMB[18][32] , \mult_22/SUMB[18][33] ,
         \mult_22/SUMB[18][34] , \mult_22/SUMB[18][35] ,
         \mult_22/SUMB[18][36] , \mult_22/SUMB[18][37] ,
         \mult_22/SUMB[18][38] , \mult_22/SUMB[18][39] ,
         \mult_22/SUMB[18][40] , \mult_22/SUMB[18][41] ,
         \mult_22/SUMB[18][42] , \mult_22/SUMB[18][43] ,
         \mult_22/SUMB[18][44] , \mult_22/SUMB[18][45] ,
         \mult_22/SUMB[18][46] , \mult_22/SUMB[18][47] ,
         \mult_22/SUMB[18][48] , \mult_22/SUMB[18][49] ,
         \mult_22/SUMB[18][50] , \mult_22/SUMB[18][51] ,
         \mult_22/SUMB[18][52] , \mult_22/SUMB[18][53] ,
         \mult_22/SUMB[18][54] , \mult_22/SUMB[18][55] ,
         \mult_22/SUMB[18][56] , \mult_22/SUMB[18][57] ,
         \mult_22/SUMB[18][58] , \mult_22/SUMB[18][59] ,
         \mult_22/SUMB[18][60] , \mult_22/SUMB[18][61] ,
         \mult_22/SUMB[18][62] , \mult_22/SUMB[19][1] , \mult_22/SUMB[19][2] ,
         \mult_22/SUMB[19][3] , \mult_22/SUMB[19][4] , \mult_22/SUMB[19][5] ,
         \mult_22/SUMB[19][6] , \mult_22/SUMB[19][7] , \mult_22/SUMB[19][8] ,
         \mult_22/SUMB[19][9] , \mult_22/SUMB[19][10] , \mult_22/SUMB[19][11] ,
         \mult_22/SUMB[19][12] , \mult_22/SUMB[19][13] ,
         \mult_22/SUMB[19][14] , \mult_22/SUMB[19][15] ,
         \mult_22/SUMB[19][16] , \mult_22/SUMB[19][17] ,
         \mult_22/SUMB[19][18] , \mult_22/SUMB[19][19] ,
         \mult_22/SUMB[19][20] , \mult_22/SUMB[19][21] ,
         \mult_22/SUMB[19][22] , \mult_22/SUMB[19][23] ,
         \mult_22/SUMB[19][24] , \mult_22/SUMB[19][25] ,
         \mult_22/SUMB[19][26] , \mult_22/SUMB[19][27] ,
         \mult_22/SUMB[19][28] , \mult_22/SUMB[19][29] ,
         \mult_22/SUMB[19][30] , \mult_22/SUMB[19][31] ,
         \mult_22/SUMB[19][32] , \mult_22/SUMB[19][33] ,
         \mult_22/SUMB[19][34] , \mult_22/SUMB[19][35] ,
         \mult_22/SUMB[19][36] , \mult_22/SUMB[19][37] ,
         \mult_22/SUMB[19][38] , \mult_22/SUMB[19][39] ,
         \mult_22/SUMB[19][40] , \mult_22/SUMB[19][41] ,
         \mult_22/SUMB[19][42] , \mult_22/SUMB[19][43] ,
         \mult_22/SUMB[19][44] , \mult_22/SUMB[19][45] ,
         \mult_22/SUMB[19][46] , \mult_22/SUMB[19][47] ,
         \mult_22/SUMB[19][48] , \mult_22/SUMB[19][49] ,
         \mult_22/SUMB[19][50] , \mult_22/SUMB[19][51] ,
         \mult_22/SUMB[19][52] , \mult_22/SUMB[19][53] ,
         \mult_22/SUMB[19][54] , \mult_22/SUMB[19][55] ,
         \mult_22/SUMB[19][56] , \mult_22/SUMB[19][57] ,
         \mult_22/SUMB[19][58] , \mult_22/SUMB[19][59] ,
         \mult_22/SUMB[19][60] , \mult_22/SUMB[19][61] ,
         \mult_22/SUMB[19][62] , \mult_22/SUMB[20][1] , \mult_22/SUMB[20][2] ,
         \mult_22/SUMB[20][3] , \mult_22/SUMB[20][4] , \mult_22/SUMB[20][5] ,
         \mult_22/SUMB[20][6] , \mult_22/SUMB[20][7] , \mult_22/SUMB[20][8] ,
         \mult_22/SUMB[20][9] , \mult_22/SUMB[20][10] , \mult_22/SUMB[20][11] ,
         \mult_22/SUMB[20][12] , \mult_22/SUMB[20][13] ,
         \mult_22/SUMB[20][14] , \mult_22/SUMB[20][15] ,
         \mult_22/SUMB[20][16] , \mult_22/SUMB[20][17] ,
         \mult_22/SUMB[20][18] , \mult_22/SUMB[20][19] ,
         \mult_22/SUMB[20][20] , \mult_22/SUMB[20][21] ,
         \mult_22/SUMB[20][22] , \mult_22/SUMB[20][23] ,
         \mult_22/SUMB[20][24] , \mult_22/SUMB[20][25] ,
         \mult_22/SUMB[20][26] , \mult_22/SUMB[20][27] ,
         \mult_22/SUMB[20][28] , \mult_22/SUMB[20][29] ,
         \mult_22/SUMB[20][30] , \mult_22/SUMB[20][31] ,
         \mult_22/SUMB[20][32] , \mult_22/SUMB[20][33] ,
         \mult_22/SUMB[20][34] , \mult_22/SUMB[20][35] ,
         \mult_22/SUMB[20][36] , \mult_22/SUMB[20][37] ,
         \mult_22/SUMB[20][38] , \mult_22/SUMB[20][39] ,
         \mult_22/SUMB[20][40] , \mult_22/SUMB[20][41] ,
         \mult_22/SUMB[20][42] , \mult_22/SUMB[20][43] ,
         \mult_22/SUMB[20][44] , \mult_22/SUMB[20][45] ,
         \mult_22/SUMB[20][46] , \mult_22/SUMB[20][47] ,
         \mult_22/SUMB[20][48] , \mult_22/SUMB[20][49] ,
         \mult_22/SUMB[20][50] , \mult_22/SUMB[20][51] ,
         \mult_22/SUMB[20][52] , \mult_22/SUMB[20][53] ,
         \mult_22/SUMB[20][54] , \mult_22/SUMB[20][55] ,
         \mult_22/SUMB[20][56] , \mult_22/SUMB[20][57] ,
         \mult_22/SUMB[20][58] , \mult_22/SUMB[20][59] ,
         \mult_22/SUMB[20][60] , \mult_22/SUMB[20][61] ,
         \mult_22/SUMB[20][62] , \mult_22/SUMB[21][1] , \mult_22/SUMB[21][2] ,
         \mult_22/SUMB[21][3] , \mult_22/SUMB[21][4] , \mult_22/SUMB[21][5] ,
         \mult_22/SUMB[21][6] , \mult_22/SUMB[21][7] , \mult_22/SUMB[21][8] ,
         \mult_22/SUMB[21][9] , \mult_22/SUMB[21][10] , \mult_22/SUMB[21][11] ,
         \mult_22/SUMB[21][12] , \mult_22/SUMB[21][13] ,
         \mult_22/SUMB[21][14] , \mult_22/SUMB[21][15] ,
         \mult_22/SUMB[21][16] , \mult_22/SUMB[21][17] ,
         \mult_22/SUMB[21][18] , \mult_22/SUMB[21][19] ,
         \mult_22/SUMB[21][20] , \mult_22/SUMB[21][21] ,
         \mult_22/SUMB[21][22] , \mult_22/SUMB[21][23] ,
         \mult_22/SUMB[21][24] , \mult_22/SUMB[21][25] ,
         \mult_22/SUMB[21][26] , \mult_22/SUMB[21][27] ,
         \mult_22/SUMB[21][28] , \mult_22/SUMB[21][29] ,
         \mult_22/SUMB[21][30] , \mult_22/SUMB[21][31] ,
         \mult_22/SUMB[21][32] , \mult_22/SUMB[21][33] ,
         \mult_22/SUMB[21][34] , \mult_22/SUMB[21][35] ,
         \mult_22/SUMB[21][36] , \mult_22/SUMB[21][37] ,
         \mult_22/SUMB[21][38] , \mult_22/SUMB[21][39] ,
         \mult_22/SUMB[21][40] , \mult_22/SUMB[21][41] ,
         \mult_22/SUMB[21][42] , \mult_22/SUMB[21][43] ,
         \mult_22/SUMB[21][44] , \mult_22/SUMB[21][45] ,
         \mult_22/SUMB[21][46] , \mult_22/SUMB[21][47] ,
         \mult_22/SUMB[21][48] , \mult_22/SUMB[21][49] ,
         \mult_22/SUMB[21][50] , \mult_22/SUMB[21][51] ,
         \mult_22/SUMB[21][52] , \mult_22/SUMB[21][53] ,
         \mult_22/SUMB[21][54] , \mult_22/SUMB[21][55] ,
         \mult_22/SUMB[21][56] , \mult_22/SUMB[21][57] ,
         \mult_22/SUMB[21][58] , \mult_22/SUMB[21][59] ,
         \mult_22/SUMB[21][60] , \mult_22/SUMB[21][61] ,
         \mult_22/SUMB[21][62] , \mult_22/SUMB[22][1] , \mult_22/SUMB[22][2] ,
         \mult_22/SUMB[22][3] , \mult_22/SUMB[22][4] , \mult_22/SUMB[22][5] ,
         \mult_22/SUMB[22][6] , \mult_22/SUMB[22][7] , \mult_22/SUMB[22][8] ,
         \mult_22/SUMB[22][9] , \mult_22/SUMB[22][10] , \mult_22/SUMB[22][11] ,
         \mult_22/SUMB[22][12] , \mult_22/SUMB[22][13] ,
         \mult_22/SUMB[22][14] , \mult_22/SUMB[22][15] ,
         \mult_22/SUMB[22][16] , \mult_22/SUMB[22][17] ,
         \mult_22/SUMB[22][18] , \mult_22/SUMB[22][19] ,
         \mult_22/SUMB[22][20] , \mult_22/SUMB[22][21] ,
         \mult_22/SUMB[22][22] , \mult_22/SUMB[22][23] ,
         \mult_22/SUMB[22][24] , \mult_22/SUMB[22][25] ,
         \mult_22/SUMB[22][26] , \mult_22/SUMB[22][27] ,
         \mult_22/SUMB[22][28] , \mult_22/SUMB[22][29] ,
         \mult_22/SUMB[22][30] , \mult_22/SUMB[22][31] ,
         \mult_22/SUMB[22][32] , \mult_22/SUMB[22][33] ,
         \mult_22/SUMB[22][34] , \mult_22/SUMB[22][35] ,
         \mult_22/SUMB[22][36] , \mult_22/SUMB[22][37] ,
         \mult_22/SUMB[22][39] , \mult_22/SUMB[22][40] ,
         \mult_22/SUMB[22][41] , \mult_22/SUMB[22][42] ,
         \mult_22/SUMB[22][43] , \mult_22/SUMB[22][44] ,
         \mult_22/SUMB[22][45] , \mult_22/SUMB[22][46] ,
         \mult_22/SUMB[22][47] , \mult_22/SUMB[22][48] ,
         \mult_22/SUMB[22][49] , \mult_22/SUMB[22][50] ,
         \mult_22/SUMB[22][51] , \mult_22/SUMB[22][52] ,
         \mult_22/SUMB[22][53] , \mult_22/SUMB[22][54] ,
         \mult_22/SUMB[22][55] , \mult_22/SUMB[22][56] ,
         \mult_22/SUMB[22][57] , \mult_22/SUMB[22][58] ,
         \mult_22/SUMB[22][59] , \mult_22/SUMB[22][60] ,
         \mult_22/SUMB[22][61] , \mult_22/SUMB[22][62] , \mult_22/SUMB[23][1] ,
         \mult_22/SUMB[23][2] , \mult_22/SUMB[23][3] , \mult_22/SUMB[23][4] ,
         \mult_22/SUMB[23][5] , \mult_22/SUMB[23][6] , \mult_22/SUMB[23][7] ,
         \mult_22/SUMB[23][8] , \mult_22/SUMB[23][9] , \mult_22/SUMB[23][10] ,
         \mult_22/SUMB[23][11] , \mult_22/SUMB[23][12] ,
         \mult_22/SUMB[23][13] , \mult_22/SUMB[23][14] ,
         \mult_22/SUMB[23][15] , \mult_22/SUMB[23][16] ,
         \mult_22/SUMB[23][17] , \mult_22/SUMB[23][18] ,
         \mult_22/SUMB[23][19] , \mult_22/SUMB[23][20] ,
         \mult_22/SUMB[23][21] , \mult_22/SUMB[23][22] ,
         \mult_22/SUMB[23][23] , \mult_22/SUMB[23][24] ,
         \mult_22/SUMB[23][25] , \mult_22/SUMB[23][26] ,
         \mult_22/SUMB[23][27] , \mult_22/SUMB[23][28] ,
         \mult_22/SUMB[23][29] , \mult_22/SUMB[23][30] ,
         \mult_22/SUMB[23][31] , \mult_22/SUMB[23][32] ,
         \mult_22/SUMB[23][33] , \mult_22/SUMB[23][34] ,
         \mult_22/SUMB[23][35] , \mult_22/SUMB[23][36] ,
         \mult_22/SUMB[23][37] , \mult_22/SUMB[23][38] ,
         \mult_22/SUMB[23][39] , \mult_22/SUMB[23][40] ,
         \mult_22/SUMB[23][41] , \mult_22/SUMB[23][42] ,
         \mult_22/SUMB[23][43] , \mult_22/SUMB[23][44] ,
         \mult_22/SUMB[23][45] , \mult_22/SUMB[23][46] ,
         \mult_22/SUMB[23][47] , \mult_22/SUMB[23][48] ,
         \mult_22/SUMB[23][49] , \mult_22/SUMB[23][50] ,
         \mult_22/SUMB[23][51] , \mult_22/SUMB[23][52] ,
         \mult_22/SUMB[23][53] , \mult_22/SUMB[23][54] ,
         \mult_22/SUMB[23][55] , \mult_22/SUMB[23][56] ,
         \mult_22/SUMB[23][57] , \mult_22/SUMB[23][58] ,
         \mult_22/SUMB[23][59] , \mult_22/SUMB[23][60] ,
         \mult_22/SUMB[23][61] , \mult_22/SUMB[23][62] ,
         \mult_22/CARRYB[16][0] , \mult_22/CARRYB[16][1] ,
         \mult_22/CARRYB[16][2] , \mult_22/CARRYB[16][3] ,
         \mult_22/CARRYB[16][4] , \mult_22/CARRYB[16][5] ,
         \mult_22/CARRYB[16][6] , \mult_22/CARRYB[16][7] ,
         \mult_22/CARRYB[16][8] , \mult_22/CARRYB[16][9] ,
         \mult_22/CARRYB[16][10] , \mult_22/CARRYB[16][11] ,
         \mult_22/CARRYB[16][12] , \mult_22/CARRYB[16][13] ,
         \mult_22/CARRYB[16][14] , \mult_22/CARRYB[16][15] ,
         \mult_22/CARRYB[16][16] , \mult_22/CARRYB[16][17] ,
         \mult_22/CARRYB[16][18] , \mult_22/CARRYB[16][19] ,
         \mult_22/CARRYB[16][20] , \mult_22/CARRYB[16][21] ,
         \mult_22/CARRYB[16][22] , \mult_22/CARRYB[16][23] ,
         \mult_22/CARRYB[16][24] , \mult_22/CARRYB[16][25] ,
         \mult_22/CARRYB[16][26] , \mult_22/CARRYB[16][27] ,
         \mult_22/CARRYB[16][28] , \mult_22/CARRYB[16][29] ,
         \mult_22/CARRYB[16][30] , \mult_22/CARRYB[16][31] ,
         \mult_22/CARRYB[16][32] , \mult_22/CARRYB[16][33] ,
         \mult_22/CARRYB[16][34] , \mult_22/CARRYB[16][35] ,
         \mult_22/CARRYB[16][36] , \mult_22/CARRYB[16][37] ,
         \mult_22/CARRYB[16][38] , \mult_22/CARRYB[16][39] ,
         \mult_22/CARRYB[16][40] , \mult_22/CARRYB[16][41] ,
         \mult_22/CARRYB[16][42] , \mult_22/CARRYB[16][43] ,
         \mult_22/CARRYB[16][44] , \mult_22/CARRYB[16][45] ,
         \mult_22/CARRYB[16][46] , \mult_22/CARRYB[16][47] ,
         \mult_22/CARRYB[16][48] , \mult_22/CARRYB[16][49] ,
         \mult_22/CARRYB[16][50] , \mult_22/CARRYB[16][51] ,
         \mult_22/CARRYB[16][52] , \mult_22/CARRYB[16][53] ,
         \mult_22/CARRYB[16][54] , \mult_22/CARRYB[16][55] ,
         \mult_22/CARRYB[16][56] , \mult_22/CARRYB[16][57] ,
         \mult_22/CARRYB[16][58] , \mult_22/CARRYB[16][59] ,
         \mult_22/CARRYB[16][60] , \mult_22/CARRYB[16][61] ,
         \mult_22/CARRYB[16][62] , \mult_22/CARRYB[17][0] ,
         \mult_22/CARRYB[17][1] , \mult_22/CARRYB[17][2] ,
         \mult_22/CARRYB[17][3] , \mult_22/CARRYB[17][4] ,
         \mult_22/CARRYB[17][5] , \mult_22/CARRYB[17][6] ,
         \mult_22/CARRYB[17][7] , \mult_22/CARRYB[17][8] ,
         \mult_22/CARRYB[17][9] , \mult_22/CARRYB[17][10] ,
         \mult_22/CARRYB[17][11] , \mult_22/CARRYB[17][12] ,
         \mult_22/CARRYB[17][13] , \mult_22/CARRYB[17][14] ,
         \mult_22/CARRYB[17][15] , \mult_22/CARRYB[17][16] ,
         \mult_22/CARRYB[17][17] , \mult_22/CARRYB[17][18] ,
         \mult_22/CARRYB[17][19] , \mult_22/CARRYB[17][20] ,
         \mult_22/CARRYB[17][21] , \mult_22/CARRYB[17][22] ,
         \mult_22/CARRYB[17][23] , \mult_22/CARRYB[17][24] ,
         \mult_22/CARRYB[17][25] , \mult_22/CARRYB[17][26] ,
         \mult_22/CARRYB[17][27] , \mult_22/CARRYB[17][28] ,
         \mult_22/CARRYB[17][29] , \mult_22/CARRYB[17][30] ,
         \mult_22/CARRYB[17][31] , \mult_22/CARRYB[17][32] ,
         \mult_22/CARRYB[17][33] , \mult_22/CARRYB[17][34] ,
         \mult_22/CARRYB[17][35] , \mult_22/CARRYB[17][36] ,
         \mult_22/CARRYB[17][37] , \mult_22/CARRYB[17][38] ,
         \mult_22/CARRYB[17][39] , \mult_22/CARRYB[17][40] ,
         \mult_22/CARRYB[17][41] , \mult_22/CARRYB[17][42] ,
         \mult_22/CARRYB[17][43] , \mult_22/CARRYB[17][44] ,
         \mult_22/CARRYB[17][45] , \mult_22/CARRYB[17][46] ,
         \mult_22/CARRYB[17][47] , \mult_22/CARRYB[17][48] ,
         \mult_22/CARRYB[17][49] , \mult_22/CARRYB[17][50] ,
         \mult_22/CARRYB[17][51] , \mult_22/CARRYB[17][52] ,
         \mult_22/CARRYB[17][53] , \mult_22/CARRYB[17][54] ,
         \mult_22/CARRYB[17][55] , \mult_22/CARRYB[17][56] ,
         \mult_22/CARRYB[17][57] , \mult_22/CARRYB[17][58] ,
         \mult_22/CARRYB[17][59] , \mult_22/CARRYB[17][60] ,
         \mult_22/CARRYB[17][61] , \mult_22/CARRYB[17][62] ,
         \mult_22/CARRYB[18][0] , \mult_22/CARRYB[18][1] ,
         \mult_22/CARRYB[18][2] , \mult_22/CARRYB[18][3] ,
         \mult_22/CARRYB[18][4] , \mult_22/CARRYB[18][5] ,
         \mult_22/CARRYB[18][6] , \mult_22/CARRYB[18][7] ,
         \mult_22/CARRYB[18][8] , \mult_22/CARRYB[18][9] ,
         \mult_22/CARRYB[18][10] , \mult_22/CARRYB[18][11] ,
         \mult_22/CARRYB[18][12] , \mult_22/CARRYB[18][13] ,
         \mult_22/CARRYB[18][14] , \mult_22/CARRYB[18][15] ,
         \mult_22/CARRYB[18][16] , \mult_22/CARRYB[18][17] ,
         \mult_22/CARRYB[18][18] , \mult_22/CARRYB[18][19] ,
         \mult_22/CARRYB[18][20] , \mult_22/CARRYB[18][21] ,
         \mult_22/CARRYB[18][22] , \mult_22/CARRYB[18][23] ,
         \mult_22/CARRYB[18][24] , \mult_22/CARRYB[18][25] ,
         \mult_22/CARRYB[18][26] , \mult_22/CARRYB[18][27] ,
         \mult_22/CARRYB[18][28] , \mult_22/CARRYB[18][29] ,
         \mult_22/CARRYB[18][30] , \mult_22/CARRYB[18][31] ,
         \mult_22/CARRYB[18][32] , \mult_22/CARRYB[18][33] ,
         \mult_22/CARRYB[18][34] , \mult_22/CARRYB[18][35] ,
         \mult_22/CARRYB[18][36] , \mult_22/CARRYB[18][37] ,
         \mult_22/CARRYB[18][38] , \mult_22/CARRYB[18][39] ,
         \mult_22/CARRYB[18][40] , \mult_22/CARRYB[18][41] ,
         \mult_22/CARRYB[18][42] , \mult_22/CARRYB[18][43] ,
         \mult_22/CARRYB[18][44] , \mult_22/CARRYB[18][45] ,
         \mult_22/CARRYB[18][46] , \mult_22/CARRYB[18][47] ,
         \mult_22/CARRYB[18][48] , \mult_22/CARRYB[18][49] ,
         \mult_22/CARRYB[18][50] , \mult_22/CARRYB[18][51] ,
         \mult_22/CARRYB[18][52] , \mult_22/CARRYB[18][53] ,
         \mult_22/CARRYB[18][54] , \mult_22/CARRYB[18][55] ,
         \mult_22/CARRYB[18][56] , \mult_22/CARRYB[18][57] ,
         \mult_22/CARRYB[18][58] , \mult_22/CARRYB[18][59] ,
         \mult_22/CARRYB[18][60] , \mult_22/CARRYB[18][61] ,
         \mult_22/CARRYB[18][62] , \mult_22/CARRYB[19][0] ,
         \mult_22/CARRYB[19][1] , \mult_22/CARRYB[19][2] ,
         \mult_22/CARRYB[19][3] , \mult_22/CARRYB[19][4] ,
         \mult_22/CARRYB[19][5] , \mult_22/CARRYB[19][6] ,
         \mult_22/CARRYB[19][7] , \mult_22/CARRYB[19][8] ,
         \mult_22/CARRYB[19][9] , \mult_22/CARRYB[19][10] ,
         \mult_22/CARRYB[19][11] , \mult_22/CARRYB[19][12] ,
         \mult_22/CARRYB[19][13] , \mult_22/CARRYB[19][14] ,
         \mult_22/CARRYB[19][15] , \mult_22/CARRYB[19][16] ,
         \mult_22/CARRYB[19][17] , \mult_22/CARRYB[19][18] ,
         \mult_22/CARRYB[19][19] , \mult_22/CARRYB[19][20] ,
         \mult_22/CARRYB[19][21] , \mult_22/CARRYB[19][22] ,
         \mult_22/CARRYB[19][23] , \mult_22/CARRYB[19][24] ,
         \mult_22/CARRYB[19][25] , \mult_22/CARRYB[19][26] ,
         \mult_22/CARRYB[19][27] , \mult_22/CARRYB[19][28] ,
         \mult_22/CARRYB[19][29] , \mult_22/CARRYB[19][30] ,
         \mult_22/CARRYB[19][31] , \mult_22/CARRYB[19][32] ,
         \mult_22/CARRYB[19][33] , \mult_22/CARRYB[19][34] ,
         \mult_22/CARRYB[19][35] , \mult_22/CARRYB[19][36] ,
         \mult_22/CARRYB[19][37] , \mult_22/CARRYB[19][38] ,
         \mult_22/CARRYB[19][39] , \mult_22/CARRYB[19][40] ,
         \mult_22/CARRYB[19][41] , \mult_22/CARRYB[19][42] ,
         \mult_22/CARRYB[19][43] , \mult_22/CARRYB[19][44] ,
         \mult_22/CARRYB[19][45] , \mult_22/CARRYB[19][46] ,
         \mult_22/CARRYB[19][47] , \mult_22/CARRYB[19][48] ,
         \mult_22/CARRYB[19][49] , \mult_22/CARRYB[19][50] ,
         \mult_22/CARRYB[19][51] , \mult_22/CARRYB[19][52] ,
         \mult_22/CARRYB[19][53] , \mult_22/CARRYB[19][54] ,
         \mult_22/CARRYB[19][55] , \mult_22/CARRYB[19][56] ,
         \mult_22/CARRYB[19][57] , \mult_22/CARRYB[19][58] ,
         \mult_22/CARRYB[19][59] , \mult_22/CARRYB[19][60] ,
         \mult_22/CARRYB[19][61] , \mult_22/CARRYB[19][62] ,
         \mult_22/CARRYB[20][0] , \mult_22/CARRYB[20][1] ,
         \mult_22/CARRYB[20][2] , \mult_22/CARRYB[20][3] ,
         \mult_22/CARRYB[20][4] , \mult_22/CARRYB[20][5] ,
         \mult_22/CARRYB[20][6] , \mult_22/CARRYB[20][7] ,
         \mult_22/CARRYB[20][8] , \mult_22/CARRYB[20][9] ,
         \mult_22/CARRYB[20][10] , \mult_22/CARRYB[20][11] ,
         \mult_22/CARRYB[20][12] , \mult_22/CARRYB[20][13] ,
         \mult_22/CARRYB[20][14] , \mult_22/CARRYB[20][15] ,
         \mult_22/CARRYB[20][16] , \mult_22/CARRYB[20][17] ,
         \mult_22/CARRYB[20][18] , \mult_22/CARRYB[20][19] ,
         \mult_22/CARRYB[20][20] , \mult_22/CARRYB[20][21] ,
         \mult_22/CARRYB[20][22] , \mult_22/CARRYB[20][23] ,
         \mult_22/CARRYB[20][24] , \mult_22/CARRYB[20][25] ,
         \mult_22/CARRYB[20][26] , \mult_22/CARRYB[20][27] ,
         \mult_22/CARRYB[20][28] , \mult_22/CARRYB[20][29] ,
         \mult_22/CARRYB[20][30] , \mult_22/CARRYB[20][31] ,
         \mult_22/CARRYB[20][32] , \mult_22/CARRYB[20][33] ,
         \mult_22/CARRYB[20][34] , \mult_22/CARRYB[20][35] ,
         \mult_22/CARRYB[20][36] , \mult_22/CARRYB[20][37] ,
         \mult_22/CARRYB[20][38] , \mult_22/CARRYB[20][39] ,
         \mult_22/CARRYB[20][40] , \mult_22/CARRYB[20][41] ,
         \mult_22/CARRYB[20][42] , \mult_22/CARRYB[20][43] ,
         \mult_22/CARRYB[20][44] , \mult_22/CARRYB[20][45] ,
         \mult_22/CARRYB[20][46] , \mult_22/CARRYB[20][47] ,
         \mult_22/CARRYB[20][48] , \mult_22/CARRYB[20][49] ,
         \mult_22/CARRYB[20][50] , \mult_22/CARRYB[20][51] ,
         \mult_22/CARRYB[20][52] , \mult_22/CARRYB[20][53] ,
         \mult_22/CARRYB[20][54] , \mult_22/CARRYB[20][55] ,
         \mult_22/CARRYB[20][56] , \mult_22/CARRYB[20][57] ,
         \mult_22/CARRYB[20][58] , \mult_22/CARRYB[20][59] ,
         \mult_22/CARRYB[20][60] , \mult_22/CARRYB[20][61] ,
         \mult_22/CARRYB[20][62] , \mult_22/CARRYB[21][0] ,
         \mult_22/CARRYB[21][1] , \mult_22/CARRYB[21][2] ,
         \mult_22/CARRYB[21][3] , \mult_22/CARRYB[21][4] ,
         \mult_22/CARRYB[21][5] , \mult_22/CARRYB[21][6] ,
         \mult_22/CARRYB[21][7] , \mult_22/CARRYB[21][8] ,
         \mult_22/CARRYB[21][9] , \mult_22/CARRYB[21][10] ,
         \mult_22/CARRYB[21][11] , \mult_22/CARRYB[21][12] ,
         \mult_22/CARRYB[21][13] , \mult_22/CARRYB[21][14] ,
         \mult_22/CARRYB[21][15] , \mult_22/CARRYB[21][16] ,
         \mult_22/CARRYB[21][17] , \mult_22/CARRYB[21][18] ,
         \mult_22/CARRYB[21][19] , \mult_22/CARRYB[21][20] ,
         \mult_22/CARRYB[21][21] , \mult_22/CARRYB[21][22] ,
         \mult_22/CARRYB[21][23] , \mult_22/CARRYB[21][24] ,
         \mult_22/CARRYB[21][25] , \mult_22/CARRYB[21][26] ,
         \mult_22/CARRYB[21][27] , \mult_22/CARRYB[21][28] ,
         \mult_22/CARRYB[21][29] , \mult_22/CARRYB[21][30] ,
         \mult_22/CARRYB[21][31] , \mult_22/CARRYB[21][32] ,
         \mult_22/CARRYB[21][33] , \mult_22/CARRYB[21][34] ,
         \mult_22/CARRYB[21][35] , \mult_22/CARRYB[21][36] ,
         \mult_22/CARRYB[21][37] , \mult_22/CARRYB[21][39] ,
         \mult_22/CARRYB[21][40] , \mult_22/CARRYB[21][41] ,
         \mult_22/CARRYB[21][42] , \mult_22/CARRYB[21][43] ,
         \mult_22/CARRYB[21][44] , \mult_22/CARRYB[21][45] ,
         \mult_22/CARRYB[21][46] , \mult_22/CARRYB[21][47] ,
         \mult_22/CARRYB[21][48] , \mult_22/CARRYB[21][49] ,
         \mult_22/CARRYB[21][50] , \mult_22/CARRYB[21][51] ,
         \mult_22/CARRYB[21][52] , \mult_22/CARRYB[21][53] ,
         \mult_22/CARRYB[21][54] , \mult_22/CARRYB[21][55] ,
         \mult_22/CARRYB[21][56] , \mult_22/CARRYB[21][57] ,
         \mult_22/CARRYB[21][58] , \mult_22/CARRYB[21][59] ,
         \mult_22/CARRYB[21][60] , \mult_22/CARRYB[21][61] ,
         \mult_22/CARRYB[21][62] , \mult_22/CARRYB[22][0] ,
         \mult_22/CARRYB[22][1] , \mult_22/CARRYB[22][2] ,
         \mult_22/CARRYB[22][3] , \mult_22/CARRYB[22][4] ,
         \mult_22/CARRYB[22][5] , \mult_22/CARRYB[22][6] ,
         \mult_22/CARRYB[22][7] , \mult_22/CARRYB[22][8] ,
         \mult_22/CARRYB[22][9] , \mult_22/CARRYB[22][10] ,
         \mult_22/CARRYB[22][11] , \mult_22/CARRYB[22][12] ,
         \mult_22/CARRYB[22][13] , \mult_22/CARRYB[22][14] ,
         \mult_22/CARRYB[22][15] , \mult_22/CARRYB[22][16] ,
         \mult_22/CARRYB[22][17] , \mult_22/CARRYB[22][18] ,
         \mult_22/CARRYB[22][19] , \mult_22/CARRYB[22][20] ,
         \mult_22/CARRYB[22][21] , \mult_22/CARRYB[22][22] ,
         \mult_22/CARRYB[22][23] , \mult_22/CARRYB[22][24] ,
         \mult_22/CARRYB[22][25] , \mult_22/CARRYB[22][26] ,
         \mult_22/CARRYB[22][27] , \mult_22/CARRYB[22][28] ,
         \mult_22/CARRYB[22][29] , \mult_22/CARRYB[22][30] ,
         \mult_22/CARRYB[22][31] , \mult_22/CARRYB[22][32] ,
         \mult_22/CARRYB[22][33] , \mult_22/CARRYB[22][34] ,
         \mult_22/CARRYB[22][35] , \mult_22/CARRYB[22][36] ,
         \mult_22/CARRYB[22][37] , \mult_22/CARRYB[22][38] ,
         \mult_22/CARRYB[22][39] , \mult_22/CARRYB[22][40] ,
         \mult_22/CARRYB[22][41] , \mult_22/CARRYB[22][42] ,
         \mult_22/CARRYB[22][43] , \mult_22/CARRYB[22][44] ,
         \mult_22/CARRYB[22][45] , \mult_22/CARRYB[22][46] ,
         \mult_22/CARRYB[22][47] , \mult_22/CARRYB[22][48] ,
         \mult_22/CARRYB[22][49] , \mult_22/CARRYB[22][50] ,
         \mult_22/CARRYB[22][51] , \mult_22/CARRYB[22][52] ,
         \mult_22/CARRYB[22][53] , \mult_22/CARRYB[22][54] ,
         \mult_22/CARRYB[22][55] , \mult_22/CARRYB[22][56] ,
         \mult_22/CARRYB[22][57] , \mult_22/CARRYB[22][58] ,
         \mult_22/CARRYB[22][59] , \mult_22/CARRYB[22][60] ,
         \mult_22/CARRYB[22][61] , \mult_22/CARRYB[22][62] ,
         \mult_22/CARRYB[23][0] , \mult_22/CARRYB[23][1] ,
         \mult_22/CARRYB[23][2] , \mult_22/CARRYB[23][3] ,
         \mult_22/CARRYB[23][4] , \mult_22/CARRYB[23][5] ,
         \mult_22/CARRYB[23][6] , \mult_22/CARRYB[23][7] ,
         \mult_22/CARRYB[23][8] , \mult_22/CARRYB[23][9] ,
         \mult_22/CARRYB[23][10] , \mult_22/CARRYB[23][11] ,
         \mult_22/CARRYB[23][12] , \mult_22/CARRYB[23][13] ,
         \mult_22/CARRYB[23][14] , \mult_22/CARRYB[23][15] ,
         \mult_22/CARRYB[23][16] , \mult_22/CARRYB[23][17] ,
         \mult_22/CARRYB[23][18] , \mult_22/CARRYB[23][19] ,
         \mult_22/CARRYB[23][20] , \mult_22/CARRYB[23][21] ,
         \mult_22/CARRYB[23][22] , \mult_22/CARRYB[23][23] ,
         \mult_22/CARRYB[23][24] , \mult_22/CARRYB[23][25] ,
         \mult_22/CARRYB[23][26] , \mult_22/CARRYB[23][27] ,
         \mult_22/CARRYB[23][28] , \mult_22/CARRYB[23][29] ,
         \mult_22/CARRYB[23][30] , \mult_22/CARRYB[23][31] ,
         \mult_22/CARRYB[23][32] , \mult_22/CARRYB[23][33] ,
         \mult_22/CARRYB[23][34] , \mult_22/CARRYB[23][35] ,
         \mult_22/CARRYB[23][36] , \mult_22/CARRYB[23][37] ,
         \mult_22/CARRYB[23][38] , \mult_22/CARRYB[23][39] ,
         \mult_22/CARRYB[23][40] , \mult_22/CARRYB[23][41] ,
         \mult_22/CARRYB[23][42] , \mult_22/CARRYB[23][43] ,
         \mult_22/CARRYB[23][44] , \mult_22/CARRYB[23][45] ,
         \mult_22/CARRYB[23][46] , \mult_22/CARRYB[23][47] ,
         \mult_22/CARRYB[23][48] , \mult_22/CARRYB[23][49] ,
         \mult_22/CARRYB[23][50] , \mult_22/CARRYB[23][51] ,
         \mult_22/CARRYB[23][52] , \mult_22/CARRYB[23][53] ,
         \mult_22/CARRYB[23][54] , \mult_22/CARRYB[23][55] ,
         \mult_22/CARRYB[23][56] , \mult_22/CARRYB[23][57] ,
         \mult_22/CARRYB[23][58] , \mult_22/CARRYB[23][59] ,
         \mult_22/CARRYB[23][60] , \mult_22/CARRYB[23][61] ,
         \mult_22/CARRYB[23][62] , \mult_22/SUMB[8][1] , \mult_22/SUMB[8][2] ,
         \mult_22/SUMB[8][3] , \mult_22/SUMB[8][4] , \mult_22/SUMB[8][5] ,
         \mult_22/SUMB[8][6] , \mult_22/SUMB[8][7] , \mult_22/SUMB[8][8] ,
         \mult_22/SUMB[8][9] , \mult_22/SUMB[8][10] , \mult_22/SUMB[8][11] ,
         \mult_22/SUMB[8][12] , \mult_22/SUMB[8][13] , \mult_22/SUMB[8][14] ,
         \mult_22/SUMB[8][15] , \mult_22/SUMB[8][16] , \mult_22/SUMB[8][17] ,
         \mult_22/SUMB[8][18] , \mult_22/SUMB[8][19] , \mult_22/SUMB[8][20] ,
         \mult_22/SUMB[8][21] , \mult_22/SUMB[8][22] , \mult_22/SUMB[8][23] ,
         \mult_22/SUMB[8][24] , \mult_22/SUMB[8][25] , \mult_22/SUMB[8][26] ,
         \mult_22/SUMB[8][27] , \mult_22/SUMB[8][28] , \mult_22/SUMB[8][29] ,
         \mult_22/SUMB[8][30] , \mult_22/SUMB[8][31] , \mult_22/SUMB[8][32] ,
         \mult_22/SUMB[8][33] , \mult_22/SUMB[8][34] , \mult_22/SUMB[8][35] ,
         \mult_22/SUMB[8][36] , \mult_22/SUMB[8][37] , \mult_22/SUMB[8][38] ,
         \mult_22/SUMB[8][39] , \mult_22/SUMB[8][40] , \mult_22/SUMB[8][41] ,
         \mult_22/SUMB[8][42] , \mult_22/SUMB[8][43] , \mult_22/SUMB[8][44] ,
         \mult_22/SUMB[8][45] , \mult_22/SUMB[8][46] , \mult_22/SUMB[8][47] ,
         \mult_22/SUMB[8][48] , \mult_22/SUMB[8][49] , \mult_22/SUMB[8][50] ,
         \mult_22/SUMB[8][51] , \mult_22/SUMB[8][52] , \mult_22/SUMB[8][53] ,
         \mult_22/SUMB[8][54] , \mult_22/SUMB[8][55] , \mult_22/SUMB[8][56] ,
         \mult_22/SUMB[8][57] , \mult_22/SUMB[8][58] , \mult_22/SUMB[8][59] ,
         \mult_22/SUMB[8][60] , \mult_22/SUMB[8][61] , \mult_22/SUMB[8][62] ,
         \mult_22/SUMB[9][1] , \mult_22/SUMB[9][2] , \mult_22/SUMB[9][3] ,
         \mult_22/SUMB[9][4] , \mult_22/SUMB[9][5] , \mult_22/SUMB[9][6] ,
         \mult_22/SUMB[9][7] , \mult_22/SUMB[9][8] , \mult_22/SUMB[9][9] ,
         \mult_22/SUMB[9][10] , \mult_22/SUMB[9][11] , \mult_22/SUMB[9][12] ,
         \mult_22/SUMB[9][13] , \mult_22/SUMB[9][14] , \mult_22/SUMB[9][15] ,
         \mult_22/SUMB[9][16] , \mult_22/SUMB[9][17] , \mult_22/SUMB[9][18] ,
         \mult_22/SUMB[9][19] , \mult_22/SUMB[9][20] , \mult_22/SUMB[9][21] ,
         \mult_22/SUMB[9][22] , \mult_22/SUMB[9][23] , \mult_22/SUMB[9][24] ,
         \mult_22/SUMB[9][25] , \mult_22/SUMB[9][26] , \mult_22/SUMB[9][27] ,
         \mult_22/SUMB[9][28] , \mult_22/SUMB[9][29] , \mult_22/SUMB[9][30] ,
         \mult_22/SUMB[9][31] , \mult_22/SUMB[9][32] , \mult_22/SUMB[9][33] ,
         \mult_22/SUMB[9][34] , \mult_22/SUMB[9][35] , \mult_22/SUMB[9][36] ,
         \mult_22/SUMB[9][37] , \mult_22/SUMB[9][38] , \mult_22/SUMB[9][39] ,
         \mult_22/SUMB[9][40] , \mult_22/SUMB[9][41] , \mult_22/SUMB[9][42] ,
         \mult_22/SUMB[9][43] , \mult_22/SUMB[9][44] , \mult_22/SUMB[9][45] ,
         \mult_22/SUMB[9][46] , \mult_22/SUMB[9][47] , \mult_22/SUMB[9][48] ,
         \mult_22/SUMB[9][49] , \mult_22/SUMB[9][50] , \mult_22/SUMB[9][51] ,
         \mult_22/SUMB[9][52] , \mult_22/SUMB[9][53] , \mult_22/SUMB[9][54] ,
         \mult_22/SUMB[9][55] , \mult_22/SUMB[9][56] , \mult_22/SUMB[9][57] ,
         \mult_22/SUMB[9][58] , \mult_22/SUMB[9][59] , \mult_22/SUMB[9][60] ,
         \mult_22/SUMB[9][61] , \mult_22/SUMB[9][62] , \mult_22/SUMB[10][1] ,
         \mult_22/SUMB[10][2] , \mult_22/SUMB[10][3] , \mult_22/SUMB[10][4] ,
         \mult_22/SUMB[10][5] , \mult_22/SUMB[10][6] , \mult_22/SUMB[10][7] ,
         \mult_22/SUMB[10][8] , \mult_22/SUMB[10][9] , \mult_22/SUMB[10][10] ,
         \mult_22/SUMB[10][11] , \mult_22/SUMB[10][12] ,
         \mult_22/SUMB[10][13] , \mult_22/SUMB[10][14] ,
         \mult_22/SUMB[10][15] , \mult_22/SUMB[10][16] ,
         \mult_22/SUMB[10][17] , \mult_22/SUMB[10][18] ,
         \mult_22/SUMB[10][19] , \mult_22/SUMB[10][20] ,
         \mult_22/SUMB[10][21] , \mult_22/SUMB[10][22] ,
         \mult_22/SUMB[10][23] , \mult_22/SUMB[10][24] ,
         \mult_22/SUMB[10][25] , \mult_22/SUMB[10][26] ,
         \mult_22/SUMB[10][27] , \mult_22/SUMB[10][28] ,
         \mult_22/SUMB[10][29] , \mult_22/SUMB[10][30] ,
         \mult_22/SUMB[10][31] , \mult_22/SUMB[10][32] ,
         \mult_22/SUMB[10][33] , \mult_22/SUMB[10][34] ,
         \mult_22/SUMB[10][35] , \mult_22/SUMB[10][36] ,
         \mult_22/SUMB[10][37] , \mult_22/SUMB[10][38] ,
         \mult_22/SUMB[10][39] , \mult_22/SUMB[10][40] ,
         \mult_22/SUMB[10][41] , \mult_22/SUMB[10][42] ,
         \mult_22/SUMB[10][43] , \mult_22/SUMB[10][44] ,
         \mult_22/SUMB[10][45] , \mult_22/SUMB[10][46] ,
         \mult_22/SUMB[10][47] , \mult_22/SUMB[10][48] ,
         \mult_22/SUMB[10][49] , \mult_22/SUMB[10][50] ,
         \mult_22/SUMB[10][51] , \mult_22/SUMB[10][52] ,
         \mult_22/SUMB[10][53] , \mult_22/SUMB[10][54] ,
         \mult_22/SUMB[10][55] , \mult_22/SUMB[10][56] ,
         \mult_22/SUMB[10][57] , \mult_22/SUMB[10][58] ,
         \mult_22/SUMB[10][59] , \mult_22/SUMB[10][60] ,
         \mult_22/SUMB[10][61] , \mult_22/SUMB[10][62] , \mult_22/SUMB[11][1] ,
         \mult_22/SUMB[11][2] , \mult_22/SUMB[11][3] , \mult_22/SUMB[11][4] ,
         \mult_22/SUMB[11][5] , \mult_22/SUMB[11][6] , \mult_22/SUMB[11][7] ,
         \mult_22/SUMB[11][8] , \mult_22/SUMB[11][9] , \mult_22/SUMB[11][10] ,
         \mult_22/SUMB[11][11] , \mult_22/SUMB[11][12] ,
         \mult_22/SUMB[11][13] , \mult_22/SUMB[11][14] ,
         \mult_22/SUMB[11][15] , \mult_22/SUMB[11][16] ,
         \mult_22/SUMB[11][17] , \mult_22/SUMB[11][18] ,
         \mult_22/SUMB[11][19] , \mult_22/SUMB[11][20] ,
         \mult_22/SUMB[11][21] , \mult_22/SUMB[11][22] ,
         \mult_22/SUMB[11][23] , \mult_22/SUMB[11][24] ,
         \mult_22/SUMB[11][25] , \mult_22/SUMB[11][26] ,
         \mult_22/SUMB[11][27] , \mult_22/SUMB[11][28] ,
         \mult_22/SUMB[11][29] , \mult_22/SUMB[11][30] ,
         \mult_22/SUMB[11][31] , \mult_22/SUMB[11][32] ,
         \mult_22/SUMB[11][33] , \mult_22/SUMB[11][34] ,
         \mult_22/SUMB[11][35] , \mult_22/SUMB[11][36] ,
         \mult_22/SUMB[11][37] , \mult_22/SUMB[11][38] ,
         \mult_22/SUMB[11][39] , \mult_22/SUMB[11][40] ,
         \mult_22/SUMB[11][41] , \mult_22/SUMB[11][42] ,
         \mult_22/SUMB[11][43] , \mult_22/SUMB[11][44] ,
         \mult_22/SUMB[11][45] , \mult_22/SUMB[11][46] ,
         \mult_22/SUMB[11][47] , \mult_22/SUMB[11][48] ,
         \mult_22/SUMB[11][49] , \mult_22/SUMB[11][50] ,
         \mult_22/SUMB[11][51] , \mult_22/SUMB[11][52] ,
         \mult_22/SUMB[11][53] , \mult_22/SUMB[11][54] ,
         \mult_22/SUMB[11][55] , \mult_22/SUMB[11][56] ,
         \mult_22/SUMB[11][57] , \mult_22/SUMB[11][58] ,
         \mult_22/SUMB[11][59] , \mult_22/SUMB[11][60] ,
         \mult_22/SUMB[11][61] , \mult_22/SUMB[11][62] , \mult_22/SUMB[12][1] ,
         \mult_22/SUMB[12][2] , \mult_22/SUMB[12][3] , \mult_22/SUMB[12][4] ,
         \mult_22/SUMB[12][5] , \mult_22/SUMB[12][6] , \mult_22/SUMB[12][7] ,
         \mult_22/SUMB[12][8] , \mult_22/SUMB[12][9] , \mult_22/SUMB[12][10] ,
         \mult_22/SUMB[12][11] , \mult_22/SUMB[12][12] ,
         \mult_22/SUMB[12][13] , \mult_22/SUMB[12][14] ,
         \mult_22/SUMB[12][15] , \mult_22/SUMB[12][16] ,
         \mult_22/SUMB[12][17] , \mult_22/SUMB[12][18] ,
         \mult_22/SUMB[12][19] , \mult_22/SUMB[12][20] ,
         \mult_22/SUMB[12][21] , \mult_22/SUMB[12][22] ,
         \mult_22/SUMB[12][23] , \mult_22/SUMB[12][24] ,
         \mult_22/SUMB[12][25] , \mult_22/SUMB[12][26] ,
         \mult_22/SUMB[12][27] , \mult_22/SUMB[12][28] ,
         \mult_22/SUMB[12][29] , \mult_22/SUMB[12][30] ,
         \mult_22/SUMB[12][31] , \mult_22/SUMB[12][32] ,
         \mult_22/SUMB[12][33] , \mult_22/SUMB[12][34] ,
         \mult_22/SUMB[12][35] , \mult_22/SUMB[12][36] ,
         \mult_22/SUMB[12][37] , \mult_22/SUMB[12][38] ,
         \mult_22/SUMB[12][39] , \mult_22/SUMB[12][40] ,
         \mult_22/SUMB[12][41] , \mult_22/SUMB[12][42] ,
         \mult_22/SUMB[12][43] , \mult_22/SUMB[12][44] ,
         \mult_22/SUMB[12][45] , \mult_22/SUMB[12][46] ,
         \mult_22/SUMB[12][47] , \mult_22/SUMB[12][48] ,
         \mult_22/SUMB[12][49] , \mult_22/SUMB[12][50] ,
         \mult_22/SUMB[12][51] , \mult_22/SUMB[12][52] ,
         \mult_22/SUMB[12][53] , \mult_22/SUMB[12][54] ,
         \mult_22/SUMB[12][55] , \mult_22/SUMB[12][56] ,
         \mult_22/SUMB[12][57] , \mult_22/SUMB[12][58] ,
         \mult_22/SUMB[12][59] , \mult_22/SUMB[12][60] ,
         \mult_22/SUMB[12][61] , \mult_22/SUMB[12][62] , \mult_22/SUMB[13][1] ,
         \mult_22/SUMB[13][2] , \mult_22/SUMB[13][3] , \mult_22/SUMB[13][4] ,
         \mult_22/SUMB[13][5] , \mult_22/SUMB[13][6] , \mult_22/SUMB[13][7] ,
         \mult_22/SUMB[13][8] , \mult_22/SUMB[13][9] , \mult_22/SUMB[13][10] ,
         \mult_22/SUMB[13][11] , \mult_22/SUMB[13][12] ,
         \mult_22/SUMB[13][13] , \mult_22/SUMB[13][14] ,
         \mult_22/SUMB[13][15] , \mult_22/SUMB[13][16] ,
         \mult_22/SUMB[13][17] , \mult_22/SUMB[13][18] ,
         \mult_22/SUMB[13][19] , \mult_22/SUMB[13][20] ,
         \mult_22/SUMB[13][21] , \mult_22/SUMB[13][22] ,
         \mult_22/SUMB[13][23] , \mult_22/SUMB[13][24] ,
         \mult_22/SUMB[13][25] , \mult_22/SUMB[13][26] ,
         \mult_22/SUMB[13][27] , \mult_22/SUMB[13][28] ,
         \mult_22/SUMB[13][29] , \mult_22/SUMB[13][30] ,
         \mult_22/SUMB[13][31] , \mult_22/SUMB[13][32] ,
         \mult_22/SUMB[13][33] , \mult_22/SUMB[13][34] ,
         \mult_22/SUMB[13][35] , \mult_22/SUMB[13][36] ,
         \mult_22/SUMB[13][37] , \mult_22/SUMB[13][38] ,
         \mult_22/SUMB[13][39] , \mult_22/SUMB[13][40] ,
         \mult_22/SUMB[13][41] , \mult_22/SUMB[13][42] ,
         \mult_22/SUMB[13][43] , \mult_22/SUMB[13][44] ,
         \mult_22/SUMB[13][45] , \mult_22/SUMB[13][46] ,
         \mult_22/SUMB[13][47] , \mult_22/SUMB[13][48] ,
         \mult_22/SUMB[13][49] , \mult_22/SUMB[13][50] ,
         \mult_22/SUMB[13][51] , \mult_22/SUMB[13][52] ,
         \mult_22/SUMB[13][53] , \mult_22/SUMB[13][54] ,
         \mult_22/SUMB[13][55] , \mult_22/SUMB[13][56] ,
         \mult_22/SUMB[13][57] , \mult_22/SUMB[13][58] ,
         \mult_22/SUMB[13][59] , \mult_22/SUMB[13][60] ,
         \mult_22/SUMB[13][61] , \mult_22/SUMB[13][62] , \mult_22/SUMB[14][1] ,
         \mult_22/SUMB[14][2] , \mult_22/SUMB[14][3] , \mult_22/SUMB[14][4] ,
         \mult_22/SUMB[14][5] , \mult_22/SUMB[14][6] , \mult_22/SUMB[14][7] ,
         \mult_22/SUMB[14][8] , \mult_22/SUMB[14][9] , \mult_22/SUMB[14][10] ,
         \mult_22/SUMB[14][11] , \mult_22/SUMB[14][12] ,
         \mult_22/SUMB[14][13] , \mult_22/SUMB[14][14] ,
         \mult_22/SUMB[14][15] , \mult_22/SUMB[14][16] ,
         \mult_22/SUMB[14][17] , \mult_22/SUMB[14][18] ,
         \mult_22/SUMB[14][19] , \mult_22/SUMB[14][20] ,
         \mult_22/SUMB[14][21] , \mult_22/SUMB[14][22] ,
         \mult_22/SUMB[14][23] , \mult_22/SUMB[14][24] ,
         \mult_22/SUMB[14][25] , \mult_22/SUMB[14][26] ,
         \mult_22/SUMB[14][27] , \mult_22/SUMB[14][28] ,
         \mult_22/SUMB[14][29] , \mult_22/SUMB[14][30] ,
         \mult_22/SUMB[14][31] , \mult_22/SUMB[14][32] ,
         \mult_22/SUMB[14][33] , \mult_22/SUMB[14][34] ,
         \mult_22/SUMB[14][35] , \mult_22/SUMB[14][36] ,
         \mult_22/SUMB[14][37] , \mult_22/SUMB[14][38] ,
         \mult_22/SUMB[14][39] , \mult_22/SUMB[14][40] ,
         \mult_22/SUMB[14][41] , \mult_22/SUMB[14][42] ,
         \mult_22/SUMB[14][43] , \mult_22/SUMB[14][44] ,
         \mult_22/SUMB[14][45] , \mult_22/SUMB[14][46] ,
         \mult_22/SUMB[14][47] , \mult_22/SUMB[14][48] ,
         \mult_22/SUMB[14][49] , \mult_22/SUMB[14][50] ,
         \mult_22/SUMB[14][51] , \mult_22/SUMB[14][52] ,
         \mult_22/SUMB[14][53] , \mult_22/SUMB[14][54] ,
         \mult_22/SUMB[14][55] , \mult_22/SUMB[14][56] ,
         \mult_22/SUMB[14][57] , \mult_22/SUMB[14][58] ,
         \mult_22/SUMB[14][59] , \mult_22/SUMB[14][60] ,
         \mult_22/SUMB[14][61] , \mult_22/SUMB[14][62] , \mult_22/SUMB[15][1] ,
         \mult_22/SUMB[15][2] , \mult_22/SUMB[15][3] , \mult_22/SUMB[15][4] ,
         \mult_22/SUMB[15][5] , \mult_22/SUMB[15][6] , \mult_22/SUMB[15][7] ,
         \mult_22/SUMB[15][8] , \mult_22/SUMB[15][9] , \mult_22/SUMB[15][10] ,
         \mult_22/SUMB[15][11] , \mult_22/SUMB[15][12] ,
         \mult_22/SUMB[15][13] , \mult_22/SUMB[15][14] ,
         \mult_22/SUMB[15][15] , \mult_22/SUMB[15][16] ,
         \mult_22/SUMB[15][17] , \mult_22/SUMB[15][18] ,
         \mult_22/SUMB[15][19] , \mult_22/SUMB[15][20] ,
         \mult_22/SUMB[15][21] , \mult_22/SUMB[15][22] ,
         \mult_22/SUMB[15][23] , \mult_22/SUMB[15][24] ,
         \mult_22/SUMB[15][25] , \mult_22/SUMB[15][26] ,
         \mult_22/SUMB[15][27] , \mult_22/SUMB[15][28] ,
         \mult_22/SUMB[15][29] , \mult_22/SUMB[15][30] ,
         \mult_22/SUMB[15][31] , \mult_22/SUMB[15][32] ,
         \mult_22/SUMB[15][33] , \mult_22/SUMB[15][34] ,
         \mult_22/SUMB[15][35] , \mult_22/SUMB[15][36] ,
         \mult_22/SUMB[15][37] , \mult_22/SUMB[15][38] ,
         \mult_22/SUMB[15][39] , \mult_22/SUMB[15][40] ,
         \mult_22/SUMB[15][41] , \mult_22/SUMB[15][42] ,
         \mult_22/SUMB[15][43] , \mult_22/SUMB[15][44] ,
         \mult_22/SUMB[15][45] , \mult_22/SUMB[15][46] ,
         \mult_22/SUMB[15][47] , \mult_22/SUMB[15][48] ,
         \mult_22/SUMB[15][49] , \mult_22/SUMB[15][50] ,
         \mult_22/SUMB[15][51] , \mult_22/SUMB[15][52] ,
         \mult_22/SUMB[15][53] , \mult_22/SUMB[15][54] ,
         \mult_22/SUMB[15][55] , \mult_22/SUMB[15][56] ,
         \mult_22/SUMB[15][57] , \mult_22/SUMB[15][58] ,
         \mult_22/SUMB[15][59] , \mult_22/SUMB[15][60] ,
         \mult_22/SUMB[15][61] , \mult_22/SUMB[15][62] ,
         \mult_22/CARRYB[8][0] , \mult_22/CARRYB[8][1] ,
         \mult_22/CARRYB[8][2] , \mult_22/CARRYB[8][3] ,
         \mult_22/CARRYB[8][4] , \mult_22/CARRYB[8][5] ,
         \mult_22/CARRYB[8][6] , \mult_22/CARRYB[8][7] ,
         \mult_22/CARRYB[8][8] , \mult_22/CARRYB[8][9] ,
         \mult_22/CARRYB[8][10] , \mult_22/CARRYB[8][11] ,
         \mult_22/CARRYB[8][12] , \mult_22/CARRYB[8][13] ,
         \mult_22/CARRYB[8][14] , \mult_22/CARRYB[8][15] ,
         \mult_22/CARRYB[8][16] , \mult_22/CARRYB[8][17] ,
         \mult_22/CARRYB[8][18] , \mult_22/CARRYB[8][19] ,
         \mult_22/CARRYB[8][20] , \mult_22/CARRYB[8][21] ,
         \mult_22/CARRYB[8][22] , \mult_22/CARRYB[8][23] ,
         \mult_22/CARRYB[8][24] , \mult_22/CARRYB[8][25] ,
         \mult_22/CARRYB[8][26] , \mult_22/CARRYB[8][27] ,
         \mult_22/CARRYB[8][28] , \mult_22/CARRYB[8][29] ,
         \mult_22/CARRYB[8][30] , \mult_22/CARRYB[8][31] ,
         \mult_22/CARRYB[8][32] , \mult_22/CARRYB[8][33] ,
         \mult_22/CARRYB[8][34] , \mult_22/CARRYB[8][35] ,
         \mult_22/CARRYB[8][36] , \mult_22/CARRYB[8][37] ,
         \mult_22/CARRYB[8][38] , \mult_22/CARRYB[8][39] ,
         \mult_22/CARRYB[8][40] , \mult_22/CARRYB[8][41] ,
         \mult_22/CARRYB[8][42] , \mult_22/CARRYB[8][43] ,
         \mult_22/CARRYB[8][44] , \mult_22/CARRYB[8][45] ,
         \mult_22/CARRYB[8][46] , \mult_22/CARRYB[8][47] ,
         \mult_22/CARRYB[8][48] , \mult_22/CARRYB[8][49] ,
         \mult_22/CARRYB[8][50] , \mult_22/CARRYB[8][51] ,
         \mult_22/CARRYB[8][52] , \mult_22/CARRYB[8][53] ,
         \mult_22/CARRYB[8][54] , \mult_22/CARRYB[8][55] ,
         \mult_22/CARRYB[8][56] , \mult_22/CARRYB[8][57] ,
         \mult_22/CARRYB[8][58] , \mult_22/CARRYB[8][59] ,
         \mult_22/CARRYB[8][60] , \mult_22/CARRYB[8][61] ,
         \mult_22/CARRYB[8][62] , \mult_22/CARRYB[9][0] ,
         \mult_22/CARRYB[9][1] , \mult_22/CARRYB[9][2] ,
         \mult_22/CARRYB[9][3] , \mult_22/CARRYB[9][4] ,
         \mult_22/CARRYB[9][5] , \mult_22/CARRYB[9][6] ,
         \mult_22/CARRYB[9][7] , \mult_22/CARRYB[9][8] ,
         \mult_22/CARRYB[9][9] , \mult_22/CARRYB[9][10] ,
         \mult_22/CARRYB[9][11] , \mult_22/CARRYB[9][12] ,
         \mult_22/CARRYB[9][13] , \mult_22/CARRYB[9][14] ,
         \mult_22/CARRYB[9][15] , \mult_22/CARRYB[9][16] ,
         \mult_22/CARRYB[9][17] , \mult_22/CARRYB[9][18] ,
         \mult_22/CARRYB[9][19] , \mult_22/CARRYB[9][20] ,
         \mult_22/CARRYB[9][21] , \mult_22/CARRYB[9][22] ,
         \mult_22/CARRYB[9][23] , \mult_22/CARRYB[9][24] ,
         \mult_22/CARRYB[9][25] , \mult_22/CARRYB[9][26] ,
         \mult_22/CARRYB[9][27] , \mult_22/CARRYB[9][28] ,
         \mult_22/CARRYB[9][29] , \mult_22/CARRYB[9][30] ,
         \mult_22/CARRYB[9][31] , \mult_22/CARRYB[9][32] ,
         \mult_22/CARRYB[9][33] , \mult_22/CARRYB[9][34] ,
         \mult_22/CARRYB[9][35] , \mult_22/CARRYB[9][36] ,
         \mult_22/CARRYB[9][37] , \mult_22/CARRYB[9][38] ,
         \mult_22/CARRYB[9][39] , \mult_22/CARRYB[9][40] ,
         \mult_22/CARRYB[9][41] , \mult_22/CARRYB[9][42] ,
         \mult_22/CARRYB[9][43] , \mult_22/CARRYB[9][44] ,
         \mult_22/CARRYB[9][45] , \mult_22/CARRYB[9][46] ,
         \mult_22/CARRYB[9][47] , \mult_22/CARRYB[9][48] ,
         \mult_22/CARRYB[9][49] , \mult_22/CARRYB[9][50] ,
         \mult_22/CARRYB[9][51] , \mult_22/CARRYB[9][52] ,
         \mult_22/CARRYB[9][53] , \mult_22/CARRYB[9][54] ,
         \mult_22/CARRYB[9][55] , \mult_22/CARRYB[9][56] ,
         \mult_22/CARRYB[9][57] , \mult_22/CARRYB[9][58] ,
         \mult_22/CARRYB[9][59] , \mult_22/CARRYB[9][60] ,
         \mult_22/CARRYB[9][61] , \mult_22/CARRYB[9][62] ,
         \mult_22/CARRYB[10][0] , \mult_22/CARRYB[10][1] ,
         \mult_22/CARRYB[10][2] , \mult_22/CARRYB[10][3] ,
         \mult_22/CARRYB[10][4] , \mult_22/CARRYB[10][5] ,
         \mult_22/CARRYB[10][6] , \mult_22/CARRYB[10][7] ,
         \mult_22/CARRYB[10][8] , \mult_22/CARRYB[10][9] ,
         \mult_22/CARRYB[10][10] , \mult_22/CARRYB[10][11] ,
         \mult_22/CARRYB[10][12] , \mult_22/CARRYB[10][13] ,
         \mult_22/CARRYB[10][14] , \mult_22/CARRYB[10][15] ,
         \mult_22/CARRYB[10][16] , \mult_22/CARRYB[10][17] ,
         \mult_22/CARRYB[10][18] , \mult_22/CARRYB[10][19] ,
         \mult_22/CARRYB[10][20] , \mult_22/CARRYB[10][21] ,
         \mult_22/CARRYB[10][22] , \mult_22/CARRYB[10][23] ,
         \mult_22/CARRYB[10][24] , \mult_22/CARRYB[10][25] ,
         \mult_22/CARRYB[10][26] , \mult_22/CARRYB[10][27] ,
         \mult_22/CARRYB[10][28] , \mult_22/CARRYB[10][29] ,
         \mult_22/CARRYB[10][30] , \mult_22/CARRYB[10][31] ,
         \mult_22/CARRYB[10][32] , \mult_22/CARRYB[10][33] ,
         \mult_22/CARRYB[10][34] , \mult_22/CARRYB[10][35] ,
         \mult_22/CARRYB[10][36] , \mult_22/CARRYB[10][37] ,
         \mult_22/CARRYB[10][38] , \mult_22/CARRYB[10][39] ,
         \mult_22/CARRYB[10][40] , \mult_22/CARRYB[10][41] ,
         \mult_22/CARRYB[10][42] , \mult_22/CARRYB[10][43] ,
         \mult_22/CARRYB[10][44] , \mult_22/CARRYB[10][45] ,
         \mult_22/CARRYB[10][46] , \mult_22/CARRYB[10][47] ,
         \mult_22/CARRYB[10][48] , \mult_22/CARRYB[10][49] ,
         \mult_22/CARRYB[10][50] , \mult_22/CARRYB[10][51] ,
         \mult_22/CARRYB[10][52] , \mult_22/CARRYB[10][53] ,
         \mult_22/CARRYB[10][54] , \mult_22/CARRYB[10][55] ,
         \mult_22/CARRYB[10][56] , \mult_22/CARRYB[10][57] ,
         \mult_22/CARRYB[10][58] , \mult_22/CARRYB[10][59] ,
         \mult_22/CARRYB[10][60] , \mult_22/CARRYB[10][61] ,
         \mult_22/CARRYB[10][62] , \mult_22/CARRYB[11][0] ,
         \mult_22/CARRYB[11][1] , \mult_22/CARRYB[11][2] ,
         \mult_22/CARRYB[11][3] , \mult_22/CARRYB[11][4] ,
         \mult_22/CARRYB[11][5] , \mult_22/CARRYB[11][6] ,
         \mult_22/CARRYB[11][7] , \mult_22/CARRYB[11][8] ,
         \mult_22/CARRYB[11][9] , \mult_22/CARRYB[11][10] ,
         \mult_22/CARRYB[11][11] , \mult_22/CARRYB[11][12] ,
         \mult_22/CARRYB[11][13] , \mult_22/CARRYB[11][14] ,
         \mult_22/CARRYB[11][15] , \mult_22/CARRYB[11][16] ,
         \mult_22/CARRYB[11][17] , \mult_22/CARRYB[11][18] ,
         \mult_22/CARRYB[11][19] , \mult_22/CARRYB[11][20] ,
         \mult_22/CARRYB[11][21] , \mult_22/CARRYB[11][22] ,
         \mult_22/CARRYB[11][23] , \mult_22/CARRYB[11][24] ,
         \mult_22/CARRYB[11][25] , \mult_22/CARRYB[11][26] ,
         \mult_22/CARRYB[11][27] , \mult_22/CARRYB[11][28] ,
         \mult_22/CARRYB[11][29] , \mult_22/CARRYB[11][30] ,
         \mult_22/CARRYB[11][31] , \mult_22/CARRYB[11][32] ,
         \mult_22/CARRYB[11][33] , \mult_22/CARRYB[11][34] ,
         \mult_22/CARRYB[11][35] , \mult_22/CARRYB[11][36] ,
         \mult_22/CARRYB[11][37] , \mult_22/CARRYB[11][38] ,
         \mult_22/CARRYB[11][39] , \mult_22/CARRYB[11][40] ,
         \mult_22/CARRYB[11][41] , \mult_22/CARRYB[11][42] ,
         \mult_22/CARRYB[11][43] , \mult_22/CARRYB[11][44] ,
         \mult_22/CARRYB[11][45] , \mult_22/CARRYB[11][46] ,
         \mult_22/CARRYB[11][47] , \mult_22/CARRYB[11][48] ,
         \mult_22/CARRYB[11][49] , \mult_22/CARRYB[11][50] ,
         \mult_22/CARRYB[11][51] , \mult_22/CARRYB[11][52] ,
         \mult_22/CARRYB[11][53] , \mult_22/CARRYB[11][54] ,
         \mult_22/CARRYB[11][55] , \mult_22/CARRYB[11][56] ,
         \mult_22/CARRYB[11][57] , \mult_22/CARRYB[11][58] ,
         \mult_22/CARRYB[11][59] , \mult_22/CARRYB[11][60] ,
         \mult_22/CARRYB[11][61] , \mult_22/CARRYB[11][62] ,
         \mult_22/CARRYB[12][0] , \mult_22/CARRYB[12][1] ,
         \mult_22/CARRYB[12][2] , \mult_22/CARRYB[12][3] ,
         \mult_22/CARRYB[12][4] , \mult_22/CARRYB[12][5] ,
         \mult_22/CARRYB[12][6] , \mult_22/CARRYB[12][7] ,
         \mult_22/CARRYB[12][8] , \mult_22/CARRYB[12][9] ,
         \mult_22/CARRYB[12][10] , \mult_22/CARRYB[12][11] ,
         \mult_22/CARRYB[12][12] , \mult_22/CARRYB[12][13] ,
         \mult_22/CARRYB[12][14] , \mult_22/CARRYB[12][15] ,
         \mult_22/CARRYB[12][16] , \mult_22/CARRYB[12][17] ,
         \mult_22/CARRYB[12][18] , \mult_22/CARRYB[12][19] ,
         \mult_22/CARRYB[12][20] , \mult_22/CARRYB[12][21] ,
         \mult_22/CARRYB[12][22] , \mult_22/CARRYB[12][23] ,
         \mult_22/CARRYB[12][24] , \mult_22/CARRYB[12][25] ,
         \mult_22/CARRYB[12][26] , \mult_22/CARRYB[12][27] ,
         \mult_22/CARRYB[12][28] , \mult_22/CARRYB[12][29] ,
         \mult_22/CARRYB[12][30] , \mult_22/CARRYB[12][31] ,
         \mult_22/CARRYB[12][32] , \mult_22/CARRYB[12][33] ,
         \mult_22/CARRYB[12][34] , \mult_22/CARRYB[12][35] ,
         \mult_22/CARRYB[12][36] , \mult_22/CARRYB[12][37] ,
         \mult_22/CARRYB[12][38] , \mult_22/CARRYB[12][39] ,
         \mult_22/CARRYB[12][40] , \mult_22/CARRYB[12][41] ,
         \mult_22/CARRYB[12][42] , \mult_22/CARRYB[12][43] ,
         \mult_22/CARRYB[12][44] , \mult_22/CARRYB[12][45] ,
         \mult_22/CARRYB[12][46] , \mult_22/CARRYB[12][47] ,
         \mult_22/CARRYB[12][48] , \mult_22/CARRYB[12][49] ,
         \mult_22/CARRYB[12][50] , \mult_22/CARRYB[12][51] ,
         \mult_22/CARRYB[12][52] , \mult_22/CARRYB[12][53] ,
         \mult_22/CARRYB[12][54] , \mult_22/CARRYB[12][55] ,
         \mult_22/CARRYB[12][56] , \mult_22/CARRYB[12][57] ,
         \mult_22/CARRYB[12][58] , \mult_22/CARRYB[12][59] ,
         \mult_22/CARRYB[12][60] , \mult_22/CARRYB[12][61] ,
         \mult_22/CARRYB[12][62] , \mult_22/CARRYB[13][0] ,
         \mult_22/CARRYB[13][1] , \mult_22/CARRYB[13][2] ,
         \mult_22/CARRYB[13][3] , \mult_22/CARRYB[13][4] ,
         \mult_22/CARRYB[13][5] , \mult_22/CARRYB[13][6] ,
         \mult_22/CARRYB[13][7] , \mult_22/CARRYB[13][8] ,
         \mult_22/CARRYB[13][9] , \mult_22/CARRYB[13][10] ,
         \mult_22/CARRYB[13][11] , \mult_22/CARRYB[13][12] ,
         \mult_22/CARRYB[13][13] , \mult_22/CARRYB[13][14] ,
         \mult_22/CARRYB[13][15] , \mult_22/CARRYB[13][16] ,
         \mult_22/CARRYB[13][17] , \mult_22/CARRYB[13][18] ,
         \mult_22/CARRYB[13][19] , \mult_22/CARRYB[13][20] ,
         \mult_22/CARRYB[13][21] , \mult_22/CARRYB[13][22] ,
         \mult_22/CARRYB[13][23] , \mult_22/CARRYB[13][24] ,
         \mult_22/CARRYB[13][25] , \mult_22/CARRYB[13][26] ,
         \mult_22/CARRYB[13][27] , \mult_22/CARRYB[13][28] ,
         \mult_22/CARRYB[13][29] , \mult_22/CARRYB[13][30] ,
         \mult_22/CARRYB[13][31] , \mult_22/CARRYB[13][32] ,
         \mult_22/CARRYB[13][33] , \mult_22/CARRYB[13][34] ,
         \mult_22/CARRYB[13][35] , \mult_22/CARRYB[13][36] ,
         \mult_22/CARRYB[13][37] , \mult_22/CARRYB[13][38] ,
         \mult_22/CARRYB[13][39] , \mult_22/CARRYB[13][40] ,
         \mult_22/CARRYB[13][41] , \mult_22/CARRYB[13][42] ,
         \mult_22/CARRYB[13][43] , \mult_22/CARRYB[13][44] ,
         \mult_22/CARRYB[13][45] , \mult_22/CARRYB[13][46] ,
         \mult_22/CARRYB[13][47] , \mult_22/CARRYB[13][48] ,
         \mult_22/CARRYB[13][49] , \mult_22/CARRYB[13][50] ,
         \mult_22/CARRYB[13][51] , \mult_22/CARRYB[13][52] ,
         \mult_22/CARRYB[13][53] , \mult_22/CARRYB[13][54] ,
         \mult_22/CARRYB[13][55] , \mult_22/CARRYB[13][56] ,
         \mult_22/CARRYB[13][57] , \mult_22/CARRYB[13][58] ,
         \mult_22/CARRYB[13][59] , \mult_22/CARRYB[13][60] ,
         \mult_22/CARRYB[13][61] , \mult_22/CARRYB[13][62] ,
         \mult_22/CARRYB[14][0] , \mult_22/CARRYB[14][1] ,
         \mult_22/CARRYB[14][2] , \mult_22/CARRYB[14][3] ,
         \mult_22/CARRYB[14][4] , \mult_22/CARRYB[14][5] ,
         \mult_22/CARRYB[14][6] , \mult_22/CARRYB[14][7] ,
         \mult_22/CARRYB[14][8] , \mult_22/CARRYB[14][9] ,
         \mult_22/CARRYB[14][10] , \mult_22/CARRYB[14][11] ,
         \mult_22/CARRYB[14][12] , \mult_22/CARRYB[14][13] ,
         \mult_22/CARRYB[14][14] , \mult_22/CARRYB[14][15] ,
         \mult_22/CARRYB[14][16] , \mult_22/CARRYB[14][17] ,
         \mult_22/CARRYB[14][18] , \mult_22/CARRYB[14][19] ,
         \mult_22/CARRYB[14][20] , \mult_22/CARRYB[14][21] ,
         \mult_22/CARRYB[14][22] , \mult_22/CARRYB[14][23] ,
         \mult_22/CARRYB[14][24] , \mult_22/CARRYB[14][25] ,
         \mult_22/CARRYB[14][26] , \mult_22/CARRYB[14][27] ,
         \mult_22/CARRYB[14][28] , \mult_22/CARRYB[14][29] ,
         \mult_22/CARRYB[14][30] , \mult_22/CARRYB[14][31] ,
         \mult_22/CARRYB[14][32] , \mult_22/CARRYB[14][33] ,
         \mult_22/CARRYB[14][34] , \mult_22/CARRYB[14][35] ,
         \mult_22/CARRYB[14][36] , \mult_22/CARRYB[14][37] ,
         \mult_22/CARRYB[14][38] , \mult_22/CARRYB[14][39] ,
         \mult_22/CARRYB[14][40] , \mult_22/CARRYB[14][41] ,
         \mult_22/CARRYB[14][42] , \mult_22/CARRYB[14][43] ,
         \mult_22/CARRYB[14][44] , \mult_22/CARRYB[14][45] ,
         \mult_22/CARRYB[14][46] , \mult_22/CARRYB[14][47] ,
         \mult_22/CARRYB[14][48] , \mult_22/CARRYB[14][49] ,
         \mult_22/CARRYB[14][50] , \mult_22/CARRYB[14][51] ,
         \mult_22/CARRYB[14][52] , \mult_22/CARRYB[14][53] ,
         \mult_22/CARRYB[14][54] , \mult_22/CARRYB[14][55] ,
         \mult_22/CARRYB[14][56] , \mult_22/CARRYB[14][57] ,
         \mult_22/CARRYB[14][58] , \mult_22/CARRYB[14][59] ,
         \mult_22/CARRYB[14][60] , \mult_22/CARRYB[14][61] ,
         \mult_22/CARRYB[14][62] , \mult_22/CARRYB[15][0] ,
         \mult_22/CARRYB[15][1] , \mult_22/CARRYB[15][2] ,
         \mult_22/CARRYB[15][3] , \mult_22/CARRYB[15][4] ,
         \mult_22/CARRYB[15][5] , \mult_22/CARRYB[15][6] ,
         \mult_22/CARRYB[15][7] , \mult_22/CARRYB[15][8] ,
         \mult_22/CARRYB[15][9] , \mult_22/CARRYB[15][10] ,
         \mult_22/CARRYB[15][11] , \mult_22/CARRYB[15][12] ,
         \mult_22/CARRYB[15][13] , \mult_22/CARRYB[15][14] ,
         \mult_22/CARRYB[15][15] , \mult_22/CARRYB[15][16] ,
         \mult_22/CARRYB[15][17] , \mult_22/CARRYB[15][18] ,
         \mult_22/CARRYB[15][19] , \mult_22/CARRYB[15][20] ,
         \mult_22/CARRYB[15][21] , \mult_22/CARRYB[15][22] ,
         \mult_22/CARRYB[15][23] , \mult_22/CARRYB[15][24] ,
         \mult_22/CARRYB[15][25] , \mult_22/CARRYB[15][26] ,
         \mult_22/CARRYB[15][27] , \mult_22/CARRYB[15][28] ,
         \mult_22/CARRYB[15][29] , \mult_22/CARRYB[15][30] ,
         \mult_22/CARRYB[15][31] , \mult_22/CARRYB[15][32] ,
         \mult_22/CARRYB[15][33] , \mult_22/CARRYB[15][34] ,
         \mult_22/CARRYB[15][35] , \mult_22/CARRYB[15][36] ,
         \mult_22/CARRYB[15][37] , \mult_22/CARRYB[15][38] ,
         \mult_22/CARRYB[15][39] , \mult_22/CARRYB[15][40] ,
         \mult_22/CARRYB[15][41] , \mult_22/CARRYB[15][42] ,
         \mult_22/CARRYB[15][43] , \mult_22/CARRYB[15][44] ,
         \mult_22/CARRYB[15][45] , \mult_22/CARRYB[15][46] ,
         \mult_22/CARRYB[15][47] , \mult_22/CARRYB[15][48] ,
         \mult_22/CARRYB[15][49] , \mult_22/CARRYB[15][50] ,
         \mult_22/CARRYB[15][51] , \mult_22/CARRYB[15][52] ,
         \mult_22/CARRYB[15][53] , \mult_22/CARRYB[15][54] ,
         \mult_22/CARRYB[15][55] , \mult_22/CARRYB[15][56] ,
         \mult_22/CARRYB[15][57] , \mult_22/CARRYB[15][58] ,
         \mult_22/CARRYB[15][59] , \mult_22/CARRYB[15][60] ,
         \mult_22/CARRYB[15][61] , \mult_22/CARRYB[15][62] ,
         \mult_22/SUMB[1][55] , \mult_22/SUMB[1][61] , \mult_22/SUMB[2][1] ,
         \mult_22/SUMB[2][2] , \mult_22/SUMB[2][3] , \mult_22/SUMB[2][4] ,
         \mult_22/SUMB[2][5] , \mult_22/SUMB[2][6] , \mult_22/SUMB[2][7] ,
         \mult_22/SUMB[2][8] , \mult_22/SUMB[2][9] , \mult_22/SUMB[2][10] ,
         \mult_22/SUMB[2][11] , \mult_22/SUMB[2][12] , \mult_22/SUMB[2][13] ,
         \mult_22/SUMB[2][14] , \mult_22/SUMB[2][15] , \mult_22/SUMB[2][16] ,
         \mult_22/SUMB[2][17] , \mult_22/SUMB[2][18] , \mult_22/SUMB[2][19] ,
         \mult_22/SUMB[2][20] , \mult_22/SUMB[2][21] , \mult_22/SUMB[2][22] ,
         \mult_22/SUMB[2][23] , \mult_22/SUMB[2][24] , \mult_22/SUMB[2][25] ,
         \mult_22/SUMB[2][26] , \mult_22/SUMB[2][27] , \mult_22/SUMB[2][28] ,
         \mult_22/SUMB[2][29] , \mult_22/SUMB[2][30] , \mult_22/SUMB[2][31] ,
         \mult_22/SUMB[2][32] , \mult_22/SUMB[2][33] , \mult_22/SUMB[2][34] ,
         \mult_22/SUMB[2][35] , \mult_22/SUMB[2][36] , \mult_22/SUMB[2][37] ,
         \mult_22/SUMB[2][38] , \mult_22/SUMB[2][39] , \mult_22/SUMB[2][40] ,
         \mult_22/SUMB[2][41] , \mult_22/SUMB[2][42] , \mult_22/SUMB[2][43] ,
         \mult_22/SUMB[2][44] , \mult_22/SUMB[2][45] , \mult_22/SUMB[2][46] ,
         \mult_22/SUMB[2][47] , \mult_22/SUMB[2][48] , \mult_22/SUMB[2][49] ,
         \mult_22/SUMB[2][50] , \mult_22/SUMB[2][51] , \mult_22/SUMB[2][52] ,
         \mult_22/SUMB[2][53] , \mult_22/SUMB[2][54] , \mult_22/SUMB[2][55] ,
         \mult_22/SUMB[2][56] , \mult_22/SUMB[2][57] , \mult_22/SUMB[2][58] ,
         \mult_22/SUMB[2][59] , \mult_22/SUMB[2][60] , \mult_22/SUMB[2][61] ,
         \mult_22/SUMB[2][62] , \mult_22/SUMB[3][1] , \mult_22/SUMB[3][2] ,
         \mult_22/SUMB[3][3] , \mult_22/SUMB[3][4] , \mult_22/SUMB[3][5] ,
         \mult_22/SUMB[3][6] , \mult_22/SUMB[3][7] , \mult_22/SUMB[3][8] ,
         \mult_22/SUMB[3][9] , \mult_22/SUMB[3][10] , \mult_22/SUMB[3][11] ,
         \mult_22/SUMB[3][12] , \mult_22/SUMB[3][13] , \mult_22/SUMB[3][14] ,
         \mult_22/SUMB[3][15] , \mult_22/SUMB[3][16] , \mult_22/SUMB[3][17] ,
         \mult_22/SUMB[3][18] , \mult_22/SUMB[3][19] , \mult_22/SUMB[3][20] ,
         \mult_22/SUMB[3][21] , \mult_22/SUMB[3][22] , \mult_22/SUMB[3][23] ,
         \mult_22/SUMB[3][24] , \mult_22/SUMB[3][25] , \mult_22/SUMB[3][26] ,
         \mult_22/SUMB[3][27] , \mult_22/SUMB[3][28] , \mult_22/SUMB[3][29] ,
         \mult_22/SUMB[3][30] , \mult_22/SUMB[3][31] , \mult_22/SUMB[3][32] ,
         \mult_22/SUMB[3][33] , \mult_22/SUMB[3][34] , \mult_22/SUMB[3][35] ,
         \mult_22/SUMB[3][36] , \mult_22/SUMB[3][37] , \mult_22/SUMB[3][38] ,
         \mult_22/SUMB[3][39] , \mult_22/SUMB[3][40] , \mult_22/SUMB[3][41] ,
         \mult_22/SUMB[3][42] , \mult_22/SUMB[3][43] , \mult_22/SUMB[3][44] ,
         \mult_22/SUMB[3][45] , \mult_22/SUMB[3][46] , \mult_22/SUMB[3][47] ,
         \mult_22/SUMB[3][48] , \mult_22/SUMB[3][49] , \mult_22/SUMB[3][50] ,
         \mult_22/SUMB[3][51] , \mult_22/SUMB[3][52] , \mult_22/SUMB[3][53] ,
         \mult_22/SUMB[3][54] , \mult_22/SUMB[3][55] , \mult_22/SUMB[3][56] ,
         \mult_22/SUMB[3][57] , \mult_22/SUMB[3][58] , \mult_22/SUMB[3][59] ,
         \mult_22/SUMB[3][60] , \mult_22/SUMB[3][61] , \mult_22/SUMB[3][62] ,
         \mult_22/SUMB[4][1] , \mult_22/SUMB[4][2] , \mult_22/SUMB[4][3] ,
         \mult_22/SUMB[4][4] , \mult_22/SUMB[4][5] , \mult_22/SUMB[4][6] ,
         \mult_22/SUMB[4][7] , \mult_22/SUMB[4][8] , \mult_22/SUMB[4][9] ,
         \mult_22/SUMB[4][10] , \mult_22/SUMB[4][11] , \mult_22/SUMB[4][12] ,
         \mult_22/SUMB[4][13] , \mult_22/SUMB[4][14] , \mult_22/SUMB[4][15] ,
         \mult_22/SUMB[4][16] , \mult_22/SUMB[4][17] , \mult_22/SUMB[4][18] ,
         \mult_22/SUMB[4][19] , \mult_22/SUMB[4][20] , \mult_22/SUMB[4][21] ,
         \mult_22/SUMB[4][22] , \mult_22/SUMB[4][23] , \mult_22/SUMB[4][24] ,
         \mult_22/SUMB[4][25] , \mult_22/SUMB[4][26] , \mult_22/SUMB[4][27] ,
         \mult_22/SUMB[4][28] , \mult_22/SUMB[4][29] , \mult_22/SUMB[4][30] ,
         \mult_22/SUMB[4][31] , \mult_22/SUMB[4][32] , \mult_22/SUMB[4][33] ,
         \mult_22/SUMB[4][34] , \mult_22/SUMB[4][35] , \mult_22/SUMB[4][36] ,
         \mult_22/SUMB[4][37] , \mult_22/SUMB[4][38] , \mult_22/SUMB[4][39] ,
         \mult_22/SUMB[4][40] , \mult_22/SUMB[4][41] , \mult_22/SUMB[4][42] ,
         \mult_22/SUMB[4][43] , \mult_22/SUMB[4][44] , \mult_22/SUMB[4][45] ,
         \mult_22/SUMB[4][46] , \mult_22/SUMB[4][47] , \mult_22/SUMB[4][48] ,
         \mult_22/SUMB[4][49] , \mult_22/SUMB[4][50] , \mult_22/SUMB[4][51] ,
         \mult_22/SUMB[4][52] , \mult_22/SUMB[4][53] , \mult_22/SUMB[4][54] ,
         \mult_22/SUMB[4][55] , \mult_22/SUMB[4][56] , \mult_22/SUMB[4][57] ,
         \mult_22/SUMB[4][58] , \mult_22/SUMB[4][59] , \mult_22/SUMB[4][60] ,
         \mult_22/SUMB[4][61] , \mult_22/SUMB[4][62] , \mult_22/SUMB[5][1] ,
         \mult_22/SUMB[5][2] , \mult_22/SUMB[5][3] , \mult_22/SUMB[5][4] ,
         \mult_22/SUMB[5][5] , \mult_22/SUMB[5][6] , \mult_22/SUMB[5][7] ,
         \mult_22/SUMB[5][8] , \mult_22/SUMB[5][9] , \mult_22/SUMB[5][10] ,
         \mult_22/SUMB[5][11] , \mult_22/SUMB[5][12] , \mult_22/SUMB[5][13] ,
         \mult_22/SUMB[5][14] , \mult_22/SUMB[5][15] , \mult_22/SUMB[5][16] ,
         \mult_22/SUMB[5][17] , \mult_22/SUMB[5][18] , \mult_22/SUMB[5][19] ,
         \mult_22/SUMB[5][20] , \mult_22/SUMB[5][21] , \mult_22/SUMB[5][22] ,
         \mult_22/SUMB[5][23] , \mult_22/SUMB[5][24] , \mult_22/SUMB[5][25] ,
         \mult_22/SUMB[5][26] , \mult_22/SUMB[5][27] , \mult_22/SUMB[5][28] ,
         \mult_22/SUMB[5][29] , \mult_22/SUMB[5][30] , \mult_22/SUMB[5][31] ,
         \mult_22/SUMB[5][32] , \mult_22/SUMB[5][33] , \mult_22/SUMB[5][34] ,
         \mult_22/SUMB[5][35] , \mult_22/SUMB[5][36] , \mult_22/SUMB[5][37] ,
         \mult_22/SUMB[5][38] , \mult_22/SUMB[5][39] , \mult_22/SUMB[5][40] ,
         \mult_22/SUMB[5][41] , \mult_22/SUMB[5][42] , \mult_22/SUMB[5][43] ,
         \mult_22/SUMB[5][44] , \mult_22/SUMB[5][45] , \mult_22/SUMB[5][46] ,
         \mult_22/SUMB[5][47] , \mult_22/SUMB[5][48] , \mult_22/SUMB[5][49] ,
         \mult_22/SUMB[5][50] , \mult_22/SUMB[5][51] , \mult_22/SUMB[5][52] ,
         \mult_22/SUMB[5][53] , \mult_22/SUMB[5][54] , \mult_22/SUMB[5][55] ,
         \mult_22/SUMB[5][56] , \mult_22/SUMB[5][57] , \mult_22/SUMB[5][58] ,
         \mult_22/SUMB[5][59] , \mult_22/SUMB[5][60] , \mult_22/SUMB[5][61] ,
         \mult_22/SUMB[5][62] , \mult_22/SUMB[6][1] , \mult_22/SUMB[6][2] ,
         \mult_22/SUMB[6][3] , \mult_22/SUMB[6][4] , \mult_22/SUMB[6][5] ,
         \mult_22/SUMB[6][6] , \mult_22/SUMB[6][7] , \mult_22/SUMB[6][8] ,
         \mult_22/SUMB[6][9] , \mult_22/SUMB[6][10] , \mult_22/SUMB[6][11] ,
         \mult_22/SUMB[6][12] , \mult_22/SUMB[6][13] , \mult_22/SUMB[6][14] ,
         \mult_22/SUMB[6][15] , \mult_22/SUMB[6][16] , \mult_22/SUMB[6][17] ,
         \mult_22/SUMB[6][18] , \mult_22/SUMB[6][19] , \mult_22/SUMB[6][20] ,
         \mult_22/SUMB[6][21] , \mult_22/SUMB[6][22] , \mult_22/SUMB[6][23] ,
         \mult_22/SUMB[6][24] , \mult_22/SUMB[6][25] , \mult_22/SUMB[6][26] ,
         \mult_22/SUMB[6][27] , \mult_22/SUMB[6][28] , \mult_22/SUMB[6][29] ,
         \mult_22/SUMB[6][30] , \mult_22/SUMB[6][31] , \mult_22/SUMB[6][32] ,
         \mult_22/SUMB[6][33] , \mult_22/SUMB[6][34] , \mult_22/SUMB[6][35] ,
         \mult_22/SUMB[6][36] , \mult_22/SUMB[6][37] , \mult_22/SUMB[6][38] ,
         \mult_22/SUMB[6][39] , \mult_22/SUMB[6][40] , \mult_22/SUMB[6][41] ,
         \mult_22/SUMB[6][42] , \mult_22/SUMB[6][43] , \mult_22/SUMB[6][44] ,
         \mult_22/SUMB[6][45] , \mult_22/SUMB[6][46] , \mult_22/SUMB[6][47] ,
         \mult_22/SUMB[6][48] , \mult_22/SUMB[6][49] , \mult_22/SUMB[6][50] ,
         \mult_22/SUMB[6][51] , \mult_22/SUMB[6][52] , \mult_22/SUMB[6][53] ,
         \mult_22/SUMB[6][54] , \mult_22/SUMB[6][55] , \mult_22/SUMB[6][56] ,
         \mult_22/SUMB[6][57] , \mult_22/SUMB[6][58] , \mult_22/SUMB[6][59] ,
         \mult_22/SUMB[6][60] , \mult_22/SUMB[6][61] , \mult_22/SUMB[6][62] ,
         \mult_22/SUMB[7][1] , \mult_22/SUMB[7][2] , \mult_22/SUMB[7][3] ,
         \mult_22/SUMB[7][4] , \mult_22/SUMB[7][5] , \mult_22/SUMB[7][6] ,
         \mult_22/SUMB[7][7] , \mult_22/SUMB[7][8] , \mult_22/SUMB[7][9] ,
         \mult_22/SUMB[7][10] , \mult_22/SUMB[7][11] , \mult_22/SUMB[7][12] ,
         \mult_22/SUMB[7][13] , \mult_22/SUMB[7][14] , \mult_22/SUMB[7][15] ,
         \mult_22/SUMB[7][16] , \mult_22/SUMB[7][17] , \mult_22/SUMB[7][18] ,
         \mult_22/SUMB[7][19] , \mult_22/SUMB[7][20] , \mult_22/SUMB[7][21] ,
         \mult_22/SUMB[7][22] , \mult_22/SUMB[7][23] , \mult_22/SUMB[7][24] ,
         \mult_22/SUMB[7][25] , \mult_22/SUMB[7][26] , \mult_22/SUMB[7][27] ,
         \mult_22/SUMB[7][28] , \mult_22/SUMB[7][29] , \mult_22/SUMB[7][30] ,
         \mult_22/SUMB[7][31] , \mult_22/SUMB[7][32] , \mult_22/SUMB[7][33] ,
         \mult_22/SUMB[7][34] , \mult_22/SUMB[7][35] , \mult_22/SUMB[7][36] ,
         \mult_22/SUMB[7][37] , \mult_22/SUMB[7][38] , \mult_22/SUMB[7][39] ,
         \mult_22/SUMB[7][40] , \mult_22/SUMB[7][41] , \mult_22/SUMB[7][42] ,
         \mult_22/SUMB[7][43] , \mult_22/SUMB[7][44] , \mult_22/SUMB[7][45] ,
         \mult_22/SUMB[7][46] , \mult_22/SUMB[7][47] , \mult_22/SUMB[7][48] ,
         \mult_22/SUMB[7][49] , \mult_22/SUMB[7][50] , \mult_22/SUMB[7][51] ,
         \mult_22/SUMB[7][52] , \mult_22/SUMB[7][53] , \mult_22/SUMB[7][54] ,
         \mult_22/SUMB[7][55] , \mult_22/SUMB[7][56] , \mult_22/SUMB[7][57] ,
         \mult_22/SUMB[7][58] , \mult_22/SUMB[7][59] , \mult_22/SUMB[7][60] ,
         \mult_22/SUMB[7][61] , \mult_22/SUMB[7][62] , \mult_22/CARRYB[1][55] ,
         \mult_22/CARRYB[1][58] , \mult_22/CARRYB[2][0] ,
         \mult_22/CARRYB[2][1] , \mult_22/CARRYB[2][2] ,
         \mult_22/CARRYB[2][3] , \mult_22/CARRYB[2][4] ,
         \mult_22/CARRYB[2][5] , \mult_22/CARRYB[2][6] ,
         \mult_22/CARRYB[2][7] , \mult_22/CARRYB[2][8] ,
         \mult_22/CARRYB[2][9] , \mult_22/CARRYB[2][10] ,
         \mult_22/CARRYB[2][11] , \mult_22/CARRYB[2][12] ,
         \mult_22/CARRYB[2][13] , \mult_22/CARRYB[2][14] ,
         \mult_22/CARRYB[2][15] , \mult_22/CARRYB[2][16] ,
         \mult_22/CARRYB[2][17] , \mult_22/CARRYB[2][18] ,
         \mult_22/CARRYB[2][19] , \mult_22/CARRYB[2][20] ,
         \mult_22/CARRYB[2][21] , \mult_22/CARRYB[2][22] ,
         \mult_22/CARRYB[2][23] , \mult_22/CARRYB[2][24] ,
         \mult_22/CARRYB[2][25] , \mult_22/CARRYB[2][26] ,
         \mult_22/CARRYB[2][27] , \mult_22/CARRYB[2][28] ,
         \mult_22/CARRYB[2][29] , \mult_22/CARRYB[2][30] ,
         \mult_22/CARRYB[2][31] , \mult_22/CARRYB[2][32] ,
         \mult_22/CARRYB[2][33] , \mult_22/CARRYB[2][34] ,
         \mult_22/CARRYB[2][35] , \mult_22/CARRYB[2][36] ,
         \mult_22/CARRYB[2][37] , \mult_22/CARRYB[2][38] ,
         \mult_22/CARRYB[2][39] , \mult_22/CARRYB[2][40] ,
         \mult_22/CARRYB[2][41] , \mult_22/CARRYB[2][42] ,
         \mult_22/CARRYB[2][43] , \mult_22/CARRYB[2][44] ,
         \mult_22/CARRYB[2][45] , \mult_22/CARRYB[2][46] ,
         \mult_22/CARRYB[2][47] , \mult_22/CARRYB[2][48] ,
         \mult_22/CARRYB[2][49] , \mult_22/CARRYB[2][50] ,
         \mult_22/CARRYB[2][51] , \mult_22/CARRYB[2][52] ,
         \mult_22/CARRYB[2][53] , \mult_22/CARRYB[2][54] ,
         \mult_22/CARRYB[2][55] , \mult_22/CARRYB[2][56] ,
         \mult_22/CARRYB[2][57] , \mult_22/CARRYB[2][58] ,
         \mult_22/CARRYB[2][59] , \mult_22/CARRYB[2][60] ,
         \mult_22/CARRYB[2][61] , \mult_22/CARRYB[2][62] ,
         \mult_22/CARRYB[3][0] , \mult_22/CARRYB[3][1] ,
         \mult_22/CARRYB[3][2] , \mult_22/CARRYB[3][3] ,
         \mult_22/CARRYB[3][4] , \mult_22/CARRYB[3][5] ,
         \mult_22/CARRYB[3][6] , \mult_22/CARRYB[3][7] ,
         \mult_22/CARRYB[3][8] , \mult_22/CARRYB[3][9] ,
         \mult_22/CARRYB[3][10] , \mult_22/CARRYB[3][11] ,
         \mult_22/CARRYB[3][12] , \mult_22/CARRYB[3][13] ,
         \mult_22/CARRYB[3][14] , \mult_22/CARRYB[3][15] ,
         \mult_22/CARRYB[3][16] , \mult_22/CARRYB[3][17] ,
         \mult_22/CARRYB[3][18] , \mult_22/CARRYB[3][19] ,
         \mult_22/CARRYB[3][20] , \mult_22/CARRYB[3][21] ,
         \mult_22/CARRYB[3][22] , \mult_22/CARRYB[3][23] ,
         \mult_22/CARRYB[3][24] , \mult_22/CARRYB[3][25] ,
         \mult_22/CARRYB[3][26] , \mult_22/CARRYB[3][27] ,
         \mult_22/CARRYB[3][28] , \mult_22/CARRYB[3][29] ,
         \mult_22/CARRYB[3][30] , \mult_22/CARRYB[3][31] ,
         \mult_22/CARRYB[3][32] , \mult_22/CARRYB[3][33] ,
         \mult_22/CARRYB[3][34] , \mult_22/CARRYB[3][35] ,
         \mult_22/CARRYB[3][36] , \mult_22/CARRYB[3][37] ,
         \mult_22/CARRYB[3][38] , \mult_22/CARRYB[3][39] ,
         \mult_22/CARRYB[3][40] , \mult_22/CARRYB[3][41] ,
         \mult_22/CARRYB[3][42] , \mult_22/CARRYB[3][43] ,
         \mult_22/CARRYB[3][44] , \mult_22/CARRYB[3][45] ,
         \mult_22/CARRYB[3][46] , \mult_22/CARRYB[3][47] ,
         \mult_22/CARRYB[3][48] , \mult_22/CARRYB[3][49] ,
         \mult_22/CARRYB[3][50] , \mult_22/CARRYB[3][51] ,
         \mult_22/CARRYB[3][52] , \mult_22/CARRYB[3][53] ,
         \mult_22/CARRYB[3][54] , \mult_22/CARRYB[3][55] ,
         \mult_22/CARRYB[3][56] , \mult_22/CARRYB[3][57] ,
         \mult_22/CARRYB[3][58] , \mult_22/CARRYB[3][59] ,
         \mult_22/CARRYB[3][60] , \mult_22/CARRYB[3][61] ,
         \mult_22/CARRYB[3][62] , \mult_22/CARRYB[4][0] ,
         \mult_22/CARRYB[4][1] , \mult_22/CARRYB[4][2] ,
         \mult_22/CARRYB[4][3] , \mult_22/CARRYB[4][4] ,
         \mult_22/CARRYB[4][5] , \mult_22/CARRYB[4][6] ,
         \mult_22/CARRYB[4][7] , \mult_22/CARRYB[4][8] ,
         \mult_22/CARRYB[4][9] , \mult_22/CARRYB[4][10] ,
         \mult_22/CARRYB[4][11] , \mult_22/CARRYB[4][12] ,
         \mult_22/CARRYB[4][13] , \mult_22/CARRYB[4][14] ,
         \mult_22/CARRYB[4][15] , \mult_22/CARRYB[4][16] ,
         \mult_22/CARRYB[4][17] , \mult_22/CARRYB[4][18] ,
         \mult_22/CARRYB[4][19] , \mult_22/CARRYB[4][20] ,
         \mult_22/CARRYB[4][21] , \mult_22/CARRYB[4][22] ,
         \mult_22/CARRYB[4][23] , \mult_22/CARRYB[4][24] ,
         \mult_22/CARRYB[4][25] , \mult_22/CARRYB[4][26] ,
         \mult_22/CARRYB[4][27] , \mult_22/CARRYB[4][28] ,
         \mult_22/CARRYB[4][29] , \mult_22/CARRYB[4][30] ,
         \mult_22/CARRYB[4][31] , \mult_22/CARRYB[4][32] ,
         \mult_22/CARRYB[4][33] , \mult_22/CARRYB[4][34] ,
         \mult_22/CARRYB[4][35] , \mult_22/CARRYB[4][36] ,
         \mult_22/CARRYB[4][37] , \mult_22/CARRYB[4][38] ,
         \mult_22/CARRYB[4][39] , \mult_22/CARRYB[4][40] ,
         \mult_22/CARRYB[4][41] , \mult_22/CARRYB[4][42] ,
         \mult_22/CARRYB[4][43] , \mult_22/CARRYB[4][44] ,
         \mult_22/CARRYB[4][45] , \mult_22/CARRYB[4][46] ,
         \mult_22/CARRYB[4][47] , \mult_22/CARRYB[4][48] ,
         \mult_22/CARRYB[4][49] , \mult_22/CARRYB[4][50] ,
         \mult_22/CARRYB[4][51] , \mult_22/CARRYB[4][52] ,
         \mult_22/CARRYB[4][53] , \mult_22/CARRYB[4][54] ,
         \mult_22/CARRYB[4][55] , \mult_22/CARRYB[4][56] ,
         \mult_22/CARRYB[4][57] , \mult_22/CARRYB[4][58] ,
         \mult_22/CARRYB[4][59] , \mult_22/CARRYB[4][60] ,
         \mult_22/CARRYB[4][61] , \mult_22/CARRYB[4][62] ,
         \mult_22/CARRYB[5][0] , \mult_22/CARRYB[5][1] ,
         \mult_22/CARRYB[5][2] , \mult_22/CARRYB[5][3] ,
         \mult_22/CARRYB[5][4] , \mult_22/CARRYB[5][5] ,
         \mult_22/CARRYB[5][6] , \mult_22/CARRYB[5][7] ,
         \mult_22/CARRYB[5][8] , \mult_22/CARRYB[5][9] ,
         \mult_22/CARRYB[5][10] , \mult_22/CARRYB[5][11] ,
         \mult_22/CARRYB[5][12] , \mult_22/CARRYB[5][13] ,
         \mult_22/CARRYB[5][14] , \mult_22/CARRYB[5][15] ,
         \mult_22/CARRYB[5][16] , \mult_22/CARRYB[5][17] ,
         \mult_22/CARRYB[5][18] , \mult_22/CARRYB[5][19] ,
         \mult_22/CARRYB[5][20] , \mult_22/CARRYB[5][21] ,
         \mult_22/CARRYB[5][22] , \mult_22/CARRYB[5][23] ,
         \mult_22/CARRYB[5][24] , \mult_22/CARRYB[5][25] ,
         \mult_22/CARRYB[5][26] , \mult_22/CARRYB[5][27] ,
         \mult_22/CARRYB[5][28] , \mult_22/CARRYB[5][29] ,
         \mult_22/CARRYB[5][30] , \mult_22/CARRYB[5][31] ,
         \mult_22/CARRYB[5][32] , \mult_22/CARRYB[5][33] ,
         \mult_22/CARRYB[5][34] , \mult_22/CARRYB[5][35] ,
         \mult_22/CARRYB[5][36] , \mult_22/CARRYB[5][37] ,
         \mult_22/CARRYB[5][38] , \mult_22/CARRYB[5][39] ,
         \mult_22/CARRYB[5][40] , \mult_22/CARRYB[5][41] ,
         \mult_22/CARRYB[5][42] , \mult_22/CARRYB[5][43] ,
         \mult_22/CARRYB[5][44] , \mult_22/CARRYB[5][45] ,
         \mult_22/CARRYB[5][46] , \mult_22/CARRYB[5][47] ,
         \mult_22/CARRYB[5][48] , \mult_22/CARRYB[5][49] ,
         \mult_22/CARRYB[5][50] , \mult_22/CARRYB[5][51] ,
         \mult_22/CARRYB[5][52] , \mult_22/CARRYB[5][53] ,
         \mult_22/CARRYB[5][54] , \mult_22/CARRYB[5][55] ,
         \mult_22/CARRYB[5][56] , \mult_22/CARRYB[5][57] ,
         \mult_22/CARRYB[5][58] , \mult_22/CARRYB[5][59] ,
         \mult_22/CARRYB[5][60] , \mult_22/CARRYB[5][61] ,
         \mult_22/CARRYB[5][62] , \mult_22/CARRYB[6][0] ,
         \mult_22/CARRYB[6][1] , \mult_22/CARRYB[6][2] ,
         \mult_22/CARRYB[6][3] , \mult_22/CARRYB[6][4] ,
         \mult_22/CARRYB[6][5] , \mult_22/CARRYB[6][6] ,
         \mult_22/CARRYB[6][7] , \mult_22/CARRYB[6][8] ,
         \mult_22/CARRYB[6][9] , \mult_22/CARRYB[6][10] ,
         \mult_22/CARRYB[6][11] , \mult_22/CARRYB[6][12] ,
         \mult_22/CARRYB[6][13] , \mult_22/CARRYB[6][14] ,
         \mult_22/CARRYB[6][15] , \mult_22/CARRYB[6][16] ,
         \mult_22/CARRYB[6][17] , \mult_22/CARRYB[6][18] ,
         \mult_22/CARRYB[6][19] , \mult_22/CARRYB[6][20] ,
         \mult_22/CARRYB[6][21] , \mult_22/CARRYB[6][22] ,
         \mult_22/CARRYB[6][23] , \mult_22/CARRYB[6][24] ,
         \mult_22/CARRYB[6][25] , \mult_22/CARRYB[6][26] ,
         \mult_22/CARRYB[6][27] , \mult_22/CARRYB[6][28] ,
         \mult_22/CARRYB[6][29] , \mult_22/CARRYB[6][30] ,
         \mult_22/CARRYB[6][31] , \mult_22/CARRYB[6][32] ,
         \mult_22/CARRYB[6][33] , \mult_22/CARRYB[6][34] ,
         \mult_22/CARRYB[6][35] , \mult_22/CARRYB[6][36] ,
         \mult_22/CARRYB[6][37] , \mult_22/CARRYB[6][38] ,
         \mult_22/CARRYB[6][39] , \mult_22/CARRYB[6][40] ,
         \mult_22/CARRYB[6][41] , \mult_22/CARRYB[6][42] ,
         \mult_22/CARRYB[6][43] , \mult_22/CARRYB[6][44] ,
         \mult_22/CARRYB[6][45] , \mult_22/CARRYB[6][46] ,
         \mult_22/CARRYB[6][47] , \mult_22/CARRYB[6][48] ,
         \mult_22/CARRYB[6][49] , \mult_22/CARRYB[6][50] ,
         \mult_22/CARRYB[6][51] , \mult_22/CARRYB[6][52] ,
         \mult_22/CARRYB[6][53] , \mult_22/CARRYB[6][54] ,
         \mult_22/CARRYB[6][55] , \mult_22/CARRYB[6][56] ,
         \mult_22/CARRYB[6][57] , \mult_22/CARRYB[6][58] ,
         \mult_22/CARRYB[6][59] , \mult_22/CARRYB[6][60] ,
         \mult_22/CARRYB[6][61] , \mult_22/CARRYB[6][62] ,
         \mult_22/CARRYB[7][0] , \mult_22/CARRYB[7][1] ,
         \mult_22/CARRYB[7][2] , \mult_22/CARRYB[7][3] ,
         \mult_22/CARRYB[7][4] , \mult_22/CARRYB[7][5] ,
         \mult_22/CARRYB[7][6] , \mult_22/CARRYB[7][7] ,
         \mult_22/CARRYB[7][8] , \mult_22/CARRYB[7][9] ,
         \mult_22/CARRYB[7][10] , \mult_22/CARRYB[7][11] ,
         \mult_22/CARRYB[7][12] , \mult_22/CARRYB[7][13] ,
         \mult_22/CARRYB[7][14] , \mult_22/CARRYB[7][15] ,
         \mult_22/CARRYB[7][16] , \mult_22/CARRYB[7][17] ,
         \mult_22/CARRYB[7][18] , \mult_22/CARRYB[7][19] ,
         \mult_22/CARRYB[7][20] , \mult_22/CARRYB[7][21] ,
         \mult_22/CARRYB[7][22] , \mult_22/CARRYB[7][23] ,
         \mult_22/CARRYB[7][24] , \mult_22/CARRYB[7][25] ,
         \mult_22/CARRYB[7][26] , \mult_22/CARRYB[7][27] ,
         \mult_22/CARRYB[7][28] , \mult_22/CARRYB[7][29] ,
         \mult_22/CARRYB[7][30] , \mult_22/CARRYB[7][31] ,
         \mult_22/CARRYB[7][32] , \mult_22/CARRYB[7][33] ,
         \mult_22/CARRYB[7][34] , \mult_22/CARRYB[7][35] ,
         \mult_22/CARRYB[7][36] , \mult_22/CARRYB[7][37] ,
         \mult_22/CARRYB[7][38] , \mult_22/CARRYB[7][39] ,
         \mult_22/CARRYB[7][40] , \mult_22/CARRYB[7][41] ,
         \mult_22/CARRYB[7][42] , \mult_22/CARRYB[7][43] ,
         \mult_22/CARRYB[7][44] , \mult_22/CARRYB[7][45] ,
         \mult_22/CARRYB[7][46] , \mult_22/CARRYB[7][47] ,
         \mult_22/CARRYB[7][48] , \mult_22/CARRYB[7][49] ,
         \mult_22/CARRYB[7][50] , \mult_22/CARRYB[7][51] ,
         \mult_22/CARRYB[7][52] , \mult_22/CARRYB[7][53] ,
         \mult_22/CARRYB[7][54] , \mult_22/CARRYB[7][55] ,
         \mult_22/CARRYB[7][56] , \mult_22/CARRYB[7][57] ,
         \mult_22/CARRYB[7][58] , \mult_22/CARRYB[7][59] ,
         \mult_22/CARRYB[7][60] , \mult_22/CARRYB[7][61] ,
         \mult_22/CARRYB[7][62] , \mult_22/ab[0][56] , \mult_22/ab[1][55] ,
         \mult_22/ab[1][63] , \mult_22/ab[2][0] , \mult_22/ab[2][1] ,
         \mult_22/ab[2][2] , \mult_22/ab[2][3] , \mult_22/ab[2][4] ,
         \mult_22/ab[2][5] , \mult_22/ab[2][6] , \mult_22/ab[2][7] ,
         \mult_22/ab[2][8] , \mult_22/ab[2][9] , \mult_22/ab[2][10] ,
         \mult_22/ab[2][11] , \mult_22/ab[2][12] , \mult_22/ab[2][13] ,
         \mult_22/ab[2][14] , \mult_22/ab[2][15] , \mult_22/ab[2][16] ,
         \mult_22/ab[2][17] , \mult_22/ab[2][18] , \mult_22/ab[2][19] ,
         \mult_22/ab[2][20] , \mult_22/ab[2][21] , \mult_22/ab[2][22] ,
         \mult_22/ab[2][23] , \mult_22/ab[2][24] , \mult_22/ab[2][25] ,
         \mult_22/ab[2][26] , \mult_22/ab[2][27] , \mult_22/ab[2][28] ,
         \mult_22/ab[2][29] , \mult_22/ab[2][30] , \mult_22/ab[2][31] ,
         \mult_22/ab[2][32] , \mult_22/ab[2][33] , \mult_22/ab[2][34] ,
         \mult_22/ab[2][35] , \mult_22/ab[2][36] , \mult_22/ab[2][37] ,
         \mult_22/ab[2][38] , \mult_22/ab[2][39] , \mult_22/ab[2][40] ,
         \mult_22/ab[2][41] , \mult_22/ab[2][42] , \mult_22/ab[2][43] ,
         \mult_22/ab[2][44] , \mult_22/ab[2][45] , \mult_22/ab[2][46] ,
         \mult_22/ab[2][47] , \mult_22/ab[2][48] , \mult_22/ab[2][49] ,
         \mult_22/ab[2][50] , \mult_22/ab[2][51] , \mult_22/ab[2][52] ,
         \mult_22/ab[2][53] , \mult_22/ab[2][54] , \mult_22/ab[2][55] ,
         \mult_22/ab[2][56] , \mult_22/ab[2][57] , \mult_22/ab[2][58] ,
         \mult_22/ab[2][59] , \mult_22/ab[2][60] , \mult_22/ab[2][61] ,
         \mult_22/ab[2][62] , \mult_22/ab[2][63] , \mult_22/ab[3][0] ,
         \mult_22/ab[3][1] , \mult_22/ab[3][2] , \mult_22/ab[3][3] ,
         \mult_22/ab[3][4] , \mult_22/ab[3][5] , \mult_22/ab[3][6] ,
         \mult_22/ab[3][7] , \mult_22/ab[3][8] , \mult_22/ab[3][9] ,
         \mult_22/ab[3][10] , \mult_22/ab[3][11] , \mult_22/ab[3][12] ,
         \mult_22/ab[3][13] , \mult_22/ab[3][14] , \mult_22/ab[3][15] ,
         \mult_22/ab[3][16] , \mult_22/ab[3][17] , \mult_22/ab[3][18] ,
         \mult_22/ab[3][19] , \mult_22/ab[3][20] , \mult_22/ab[3][21] ,
         \mult_22/ab[3][22] , \mult_22/ab[3][23] , \mult_22/ab[3][24] ,
         \mult_22/ab[3][25] , \mult_22/ab[3][26] , \mult_22/ab[3][27] ,
         \mult_22/ab[3][28] , \mult_22/ab[3][29] , \mult_22/ab[3][30] ,
         \mult_22/ab[3][31] , \mult_22/ab[3][32] , \mult_22/ab[3][33] ,
         \mult_22/ab[3][34] , \mult_22/ab[3][35] , \mult_22/ab[3][36] ,
         \mult_22/ab[3][37] , \mult_22/ab[3][38] , \mult_22/ab[3][39] ,
         \mult_22/ab[3][40] , \mult_22/ab[3][41] , \mult_22/ab[3][42] ,
         \mult_22/ab[3][43] , \mult_22/ab[3][44] , \mult_22/ab[3][45] ,
         \mult_22/ab[3][46] , \mult_22/ab[3][47] , \mult_22/ab[3][48] ,
         \mult_22/ab[3][49] , \mult_22/ab[3][50] , \mult_22/ab[3][51] ,
         \mult_22/ab[3][52] , \mult_22/ab[3][53] , \mult_22/ab[3][54] ,
         \mult_22/ab[3][55] , \mult_22/ab[3][57] , \mult_22/ab[3][58] ,
         \mult_22/ab[3][59] , \mult_22/ab[3][60] , \mult_22/ab[3][61] ,
         \mult_22/ab[3][62] , \mult_22/ab[3][63] , \mult_22/ab[4][0] ,
         \mult_22/ab[4][1] , \mult_22/ab[4][2] , \mult_22/ab[4][3] ,
         \mult_22/ab[4][4] , \mult_22/ab[4][5] , \mult_22/ab[4][6] ,
         \mult_22/ab[4][7] , \mult_22/ab[4][8] , \mult_22/ab[4][9] ,
         \mult_22/ab[4][10] , \mult_22/ab[4][11] , \mult_22/ab[4][12] ,
         \mult_22/ab[4][13] , \mult_22/ab[4][14] , \mult_22/ab[4][15] ,
         \mult_22/ab[4][16] , \mult_22/ab[4][17] , \mult_22/ab[4][18] ,
         \mult_22/ab[4][19] , \mult_22/ab[4][20] , \mult_22/ab[4][21] ,
         \mult_22/ab[4][22] , \mult_22/ab[4][23] , \mult_22/ab[4][24] ,
         \mult_22/ab[4][25] , \mult_22/ab[4][26] , \mult_22/ab[4][27] ,
         \mult_22/ab[4][28] , \mult_22/ab[4][29] , \mult_22/ab[4][30] ,
         \mult_22/ab[4][31] , \mult_22/ab[4][32] , \mult_22/ab[4][33] ,
         \mult_22/ab[4][34] , \mult_22/ab[4][35] , \mult_22/ab[4][36] ,
         \mult_22/ab[4][37] , \mult_22/ab[4][38] , \mult_22/ab[4][39] ,
         \mult_22/ab[4][40] , \mult_22/ab[4][41] , \mult_22/ab[4][42] ,
         \mult_22/ab[4][43] , \mult_22/ab[4][44] , \mult_22/ab[4][45] ,
         \mult_22/ab[4][46] , \mult_22/ab[4][47] , \mult_22/ab[4][48] ,
         \mult_22/ab[4][49] , \mult_22/ab[4][50] , \mult_22/ab[4][51] ,
         \mult_22/ab[4][53] , \mult_22/ab[4][54] , \mult_22/ab[4][55] ,
         \mult_22/ab[4][56] , \mult_22/ab[4][57] , \mult_22/ab[4][58] ,
         \mult_22/ab[4][59] , \mult_22/ab[4][60] , \mult_22/ab[4][61] ,
         \mult_22/ab[4][62] , \mult_22/ab[4][63] , \mult_22/ab[5][0] ,
         \mult_22/ab[5][1] , \mult_22/ab[5][2] , \mult_22/ab[5][3] ,
         \mult_22/ab[5][4] , \mult_22/ab[5][5] , \mult_22/ab[5][6] ,
         \mult_22/ab[5][7] , \mult_22/ab[5][8] , \mult_22/ab[5][9] ,
         \mult_22/ab[5][10] , \mult_22/ab[5][11] , \mult_22/ab[5][12] ,
         \mult_22/ab[5][13] , \mult_22/ab[5][14] , \mult_22/ab[5][15] ,
         \mult_22/ab[5][16] , \mult_22/ab[5][17] , \mult_22/ab[5][18] ,
         \mult_22/ab[5][19] , \mult_22/ab[5][20] , \mult_22/ab[5][21] ,
         \mult_22/ab[5][22] , \mult_22/ab[5][23] , \mult_22/ab[5][24] ,
         \mult_22/ab[5][25] , \mult_22/ab[5][26] , \mult_22/ab[5][27] ,
         \mult_22/ab[5][28] , \mult_22/ab[5][29] , \mult_22/ab[5][30] ,
         \mult_22/ab[5][31] , \mult_22/ab[5][32] , \mult_22/ab[5][33] ,
         \mult_22/ab[5][34] , \mult_22/ab[5][35] , \mult_22/ab[5][36] ,
         \mult_22/ab[5][37] , \mult_22/ab[5][38] , \mult_22/ab[5][39] ,
         \mult_22/ab[5][40] , \mult_22/ab[5][41] , \mult_22/ab[5][42] ,
         \mult_22/ab[5][43] , \mult_22/ab[5][44] , \mult_22/ab[5][45] ,
         \mult_22/ab[5][46] , \mult_22/ab[5][47] , \mult_22/ab[5][48] ,
         \mult_22/ab[5][49] , \mult_22/ab[5][50] , \mult_22/ab[5][51] ,
         \mult_22/ab[5][52] , \mult_22/ab[5][53] , \mult_22/ab[5][54] ,
         \mult_22/ab[5][55] , \mult_22/ab[5][56] , \mult_22/ab[5][57] ,
         \mult_22/ab[5][58] , \mult_22/ab[5][59] , \mult_22/ab[5][60] ,
         \mult_22/ab[5][61] , \mult_22/ab[5][62] , \mult_22/ab[5][63] ,
         \mult_22/ab[6][0] , \mult_22/ab[6][1] , \mult_22/ab[6][2] ,
         \mult_22/ab[6][3] , \mult_22/ab[6][4] , \mult_22/ab[6][5] ,
         \mult_22/ab[6][6] , \mult_22/ab[6][7] , \mult_22/ab[6][8] ,
         \mult_22/ab[6][9] , \mult_22/ab[6][10] , \mult_22/ab[6][11] ,
         \mult_22/ab[6][12] , \mult_22/ab[6][13] , \mult_22/ab[6][14] ,
         \mult_22/ab[6][15] , \mult_22/ab[6][16] , \mult_22/ab[6][17] ,
         \mult_22/ab[6][18] , \mult_22/ab[6][19] , \mult_22/ab[6][20] ,
         \mult_22/ab[6][21] , \mult_22/ab[6][22] , \mult_22/ab[6][23] ,
         \mult_22/ab[6][24] , \mult_22/ab[6][25] , \mult_22/ab[6][26] ,
         \mult_22/ab[6][27] , \mult_22/ab[6][28] , \mult_22/ab[6][29] ,
         \mult_22/ab[6][30] , \mult_22/ab[6][31] , \mult_22/ab[6][32] ,
         \mult_22/ab[6][33] , \mult_22/ab[6][34] , \mult_22/ab[6][35] ,
         \mult_22/ab[6][36] , \mult_22/ab[6][37] , \mult_22/ab[6][38] ,
         \mult_22/ab[6][39] , \mult_22/ab[6][40] , \mult_22/ab[6][41] ,
         \mult_22/ab[6][42] , \mult_22/ab[6][43] , \mult_22/ab[6][44] ,
         \mult_22/ab[6][45] , \mult_22/ab[6][46] , \mult_22/ab[6][47] ,
         \mult_22/ab[6][48] , \mult_22/ab[6][49] , \mult_22/ab[6][50] ,
         \mult_22/ab[6][51] , \mult_22/ab[6][52] , \mult_22/ab[6][53] ,
         \mult_22/ab[6][54] , \mult_22/ab[6][55] , \mult_22/ab[6][56] ,
         \mult_22/ab[6][57] , \mult_22/ab[6][58] , \mult_22/ab[6][59] ,
         \mult_22/ab[6][60] , \mult_22/ab[6][61] , \mult_22/ab[6][62] ,
         \mult_22/ab[6][63] , \mult_22/ab[7][0] , \mult_22/ab[7][1] ,
         \mult_22/ab[7][2] , \mult_22/ab[7][3] , \mult_22/ab[7][4] ,
         \mult_22/ab[7][5] , \mult_22/ab[7][6] , \mult_22/ab[7][7] ,
         \mult_22/ab[7][8] , \mult_22/ab[7][9] , \mult_22/ab[7][10] ,
         \mult_22/ab[7][11] , \mult_22/ab[7][12] , \mult_22/ab[7][13] ,
         \mult_22/ab[7][14] , \mult_22/ab[7][15] , \mult_22/ab[7][16] ,
         \mult_22/ab[7][17] , \mult_22/ab[7][18] , \mult_22/ab[7][19] ,
         \mult_22/ab[7][20] , \mult_22/ab[7][21] , \mult_22/ab[7][22] ,
         \mult_22/ab[7][23] , \mult_22/ab[7][24] , \mult_22/ab[7][25] ,
         \mult_22/ab[7][26] , \mult_22/ab[7][27] , \mult_22/ab[7][28] ,
         \mult_22/ab[7][29] , \mult_22/ab[7][30] , \mult_22/ab[7][31] ,
         \mult_22/ab[7][32] , \mult_22/ab[7][33] , \mult_22/ab[7][34] ,
         \mult_22/ab[7][35] , \mult_22/ab[7][36] , \mult_22/ab[7][37] ,
         \mult_22/ab[7][38] , \mult_22/ab[7][39] , \mult_22/ab[7][40] ,
         \mult_22/ab[7][41] , \mult_22/ab[7][42] , \mult_22/ab[7][43] ,
         \mult_22/ab[7][44] , \mult_22/ab[7][45] , \mult_22/ab[7][46] ,
         \mult_22/ab[7][47] , \mult_22/ab[7][48] , \mult_22/ab[7][49] ,
         \mult_22/ab[7][50] , \mult_22/ab[7][51] , \mult_22/ab[7][52] ,
         \mult_22/ab[7][53] , \mult_22/ab[7][54] , \mult_22/ab[7][55] ,
         \mult_22/ab[7][56] , \mult_22/ab[7][57] , \mult_22/ab[7][58] ,
         \mult_22/ab[7][59] , \mult_22/ab[7][60] , \mult_22/ab[7][61] ,
         \mult_22/ab[7][62] , \mult_22/ab[7][63] , \mult_22/ab[8][0] ,
         \mult_22/ab[8][1] , \mult_22/ab[8][2] , \mult_22/ab[8][3] ,
         \mult_22/ab[8][4] , \mult_22/ab[8][5] , \mult_22/ab[8][6] ,
         \mult_22/ab[8][7] , \mult_22/ab[8][8] , \mult_22/ab[8][9] ,
         \mult_22/ab[8][10] , \mult_22/ab[8][11] , \mult_22/ab[8][12] ,
         \mult_22/ab[8][13] , \mult_22/ab[8][14] , \mult_22/ab[8][15] ,
         \mult_22/ab[8][16] , \mult_22/ab[8][17] , \mult_22/ab[8][18] ,
         \mult_22/ab[8][19] , \mult_22/ab[8][20] , \mult_22/ab[8][21] ,
         \mult_22/ab[8][22] , \mult_22/ab[8][23] , \mult_22/ab[8][24] ,
         \mult_22/ab[8][25] , \mult_22/ab[8][26] , \mult_22/ab[8][27] ,
         \mult_22/ab[8][28] , \mult_22/ab[8][29] , \mult_22/ab[8][30] ,
         \mult_22/ab[8][31] , \mult_22/ab[8][32] , \mult_22/ab[8][33] ,
         \mult_22/ab[8][34] , \mult_22/ab[8][35] , \mult_22/ab[8][36] ,
         \mult_22/ab[8][37] , \mult_22/ab[8][38] , \mult_22/ab[8][39] ,
         \mult_22/ab[8][40] , \mult_22/ab[8][41] , \mult_22/ab[8][42] ,
         \mult_22/ab[8][43] , \mult_22/ab[8][44] , \mult_22/ab[8][45] ,
         \mult_22/ab[8][46] , \mult_22/ab[8][47] , \mult_22/ab[8][48] ,
         \mult_22/ab[8][49] , \mult_22/ab[8][51] , \mult_22/ab[8][52] ,
         \mult_22/ab[8][53] , \mult_22/ab[8][54] , \mult_22/ab[8][55] ,
         \mult_22/ab[8][56] , \mult_22/ab[8][57] , \mult_22/ab[8][58] ,
         \mult_22/ab[8][59] , \mult_22/ab[8][60] , \mult_22/ab[8][61] ,
         \mult_22/ab[8][62] , \mult_22/ab[8][63] , \mult_22/ab[9][0] ,
         \mult_22/ab[9][1] , \mult_22/ab[9][2] , \mult_22/ab[9][3] ,
         \mult_22/ab[9][4] , \mult_22/ab[9][5] , \mult_22/ab[9][6] ,
         \mult_22/ab[9][7] , \mult_22/ab[9][8] , \mult_22/ab[9][9] ,
         \mult_22/ab[9][10] , \mult_22/ab[9][11] , \mult_22/ab[9][12] ,
         \mult_22/ab[9][13] , \mult_22/ab[9][14] , \mult_22/ab[9][15] ,
         \mult_22/ab[9][16] , \mult_22/ab[9][17] , \mult_22/ab[9][18] ,
         \mult_22/ab[9][19] , \mult_22/ab[9][20] , \mult_22/ab[9][21] ,
         \mult_22/ab[9][22] , \mult_22/ab[9][23] , \mult_22/ab[9][24] ,
         \mult_22/ab[9][25] , \mult_22/ab[9][26] , \mult_22/ab[9][27] ,
         \mult_22/ab[9][28] , \mult_22/ab[9][29] , \mult_22/ab[9][30] ,
         \mult_22/ab[9][31] , \mult_22/ab[9][32] , \mult_22/ab[9][33] ,
         \mult_22/ab[9][34] , \mult_22/ab[9][35] , \mult_22/ab[9][36] ,
         \mult_22/ab[9][37] , \mult_22/ab[9][38] , \mult_22/ab[9][39] ,
         \mult_22/ab[9][40] , \mult_22/ab[9][41] , \mult_22/ab[9][42] ,
         \mult_22/ab[9][43] , \mult_22/ab[9][44] , \mult_22/ab[9][45] ,
         \mult_22/ab[9][46] , \mult_22/ab[9][47] , \mult_22/ab[9][48] ,
         \mult_22/ab[9][49] , \mult_22/ab[9][50] , \mult_22/ab[9][51] ,
         \mult_22/ab[9][52] , \mult_22/ab[9][53] , \mult_22/ab[9][54] ,
         \mult_22/ab[9][55] , \mult_22/ab[9][56] , \mult_22/ab[9][57] ,
         \mult_22/ab[9][58] , \mult_22/ab[9][59] , \mult_22/ab[9][60] ,
         \mult_22/ab[9][61] , \mult_22/ab[9][62] , \mult_22/ab[9][63] ,
         \mult_22/ab[10][0] , \mult_22/ab[10][1] , \mult_22/ab[10][2] ,
         \mult_22/ab[10][3] , \mult_22/ab[10][4] , \mult_22/ab[10][5] ,
         \mult_22/ab[10][6] , \mult_22/ab[10][7] , \mult_22/ab[10][8] ,
         \mult_22/ab[10][9] , \mult_22/ab[10][10] , \mult_22/ab[10][11] ,
         \mult_22/ab[10][12] , \mult_22/ab[10][13] , \mult_22/ab[10][14] ,
         \mult_22/ab[10][15] , \mult_22/ab[10][16] , \mult_22/ab[10][17] ,
         \mult_22/ab[10][18] , \mult_22/ab[10][19] , \mult_22/ab[10][20] ,
         \mult_22/ab[10][21] , \mult_22/ab[10][22] , \mult_22/ab[10][23] ,
         \mult_22/ab[10][24] , \mult_22/ab[10][25] , \mult_22/ab[10][26] ,
         \mult_22/ab[10][27] , \mult_22/ab[10][28] , \mult_22/ab[10][29] ,
         \mult_22/ab[10][30] , \mult_22/ab[10][31] , \mult_22/ab[10][32] ,
         \mult_22/ab[10][33] , \mult_22/ab[10][34] , \mult_22/ab[10][35] ,
         \mult_22/ab[10][36] , \mult_22/ab[10][37] , \mult_22/ab[10][38] ,
         \mult_22/ab[10][39] , \mult_22/ab[10][40] , \mult_22/ab[10][41] ,
         \mult_22/ab[10][42] , \mult_22/ab[10][43] , \mult_22/ab[10][44] ,
         \mult_22/ab[10][45] , \mult_22/ab[10][46] , \mult_22/ab[10][47] ,
         \mult_22/ab[10][48] , \mult_22/ab[10][49] , \mult_22/ab[10][50] ,
         \mult_22/ab[10][51] , \mult_22/ab[10][52] , \mult_22/ab[10][53] ,
         \mult_22/ab[10][54] , \mult_22/ab[10][55] , \mult_22/ab[10][56] ,
         \mult_22/ab[10][57] , \mult_22/ab[10][58] , \mult_22/ab[10][59] ,
         \mult_22/ab[10][60] , \mult_22/ab[10][61] , \mult_22/ab[10][62] ,
         \mult_22/ab[10][63] , \mult_22/ab[11][0] , \mult_22/ab[11][1] ,
         \mult_22/ab[11][2] , \mult_22/ab[11][3] , \mult_22/ab[11][4] ,
         \mult_22/ab[11][5] , \mult_22/ab[11][6] , \mult_22/ab[11][7] ,
         \mult_22/ab[11][8] , \mult_22/ab[11][9] , \mult_22/ab[11][10] ,
         \mult_22/ab[11][11] , \mult_22/ab[11][12] , \mult_22/ab[11][13] ,
         \mult_22/ab[11][14] , \mult_22/ab[11][15] , \mult_22/ab[11][16] ,
         \mult_22/ab[11][17] , \mult_22/ab[11][18] , \mult_22/ab[11][19] ,
         \mult_22/ab[11][20] , \mult_22/ab[11][21] , \mult_22/ab[11][22] ,
         \mult_22/ab[11][23] , \mult_22/ab[11][24] , \mult_22/ab[11][25] ,
         \mult_22/ab[11][26] , \mult_22/ab[11][27] , \mult_22/ab[11][28] ,
         \mult_22/ab[11][29] , \mult_22/ab[11][30] , \mult_22/ab[11][31] ,
         \mult_22/ab[11][32] , \mult_22/ab[11][33] , \mult_22/ab[11][34] ,
         \mult_22/ab[11][35] , \mult_22/ab[11][36] , \mult_22/ab[11][37] ,
         \mult_22/ab[11][38] , \mult_22/ab[11][39] , \mult_22/ab[11][40] ,
         \mult_22/ab[11][41] , \mult_22/ab[11][42] , \mult_22/ab[11][43] ,
         \mult_22/ab[11][44] , \mult_22/ab[11][45] , \mult_22/ab[11][47] ,
         \mult_22/ab[11][48] , \mult_22/ab[11][49] , \mult_22/ab[11][50] ,
         \mult_22/ab[11][51] , \mult_22/ab[11][52] , \mult_22/ab[11][53] ,
         \mult_22/ab[11][54] , \mult_22/ab[11][55] , \mult_22/ab[11][56] ,
         \mult_22/ab[11][57] , \mult_22/ab[11][58] , \mult_22/ab[11][59] ,
         \mult_22/ab[11][60] , \mult_22/ab[11][61] , \mult_22/ab[11][62] ,
         \mult_22/ab[11][63] , \mult_22/ab[12][0] , \mult_22/ab[12][1] ,
         \mult_22/ab[12][2] , \mult_22/ab[12][3] , \mult_22/ab[12][4] ,
         \mult_22/ab[12][5] , \mult_22/ab[12][6] , \mult_22/ab[12][7] ,
         \mult_22/ab[12][8] , \mult_22/ab[12][9] , \mult_22/ab[12][10] ,
         \mult_22/ab[12][11] , \mult_22/ab[12][12] , \mult_22/ab[12][13] ,
         \mult_22/ab[12][14] , \mult_22/ab[12][15] , \mult_22/ab[12][16] ,
         \mult_22/ab[12][17] , \mult_22/ab[12][18] , \mult_22/ab[12][19] ,
         \mult_22/ab[12][20] , \mult_22/ab[12][21] , \mult_22/ab[12][22] ,
         \mult_22/ab[12][23] , \mult_22/ab[12][24] , \mult_22/ab[12][25] ,
         \mult_22/ab[12][26] , \mult_22/ab[12][27] , \mult_22/ab[12][28] ,
         \mult_22/ab[12][29] , \mult_22/ab[12][30] , \mult_22/ab[12][31] ,
         \mult_22/ab[12][32] , \mult_22/ab[12][33] , \mult_22/ab[12][34] ,
         \mult_22/ab[12][35] , \mult_22/ab[12][36] , \mult_22/ab[12][37] ,
         \mult_22/ab[12][38] , \mult_22/ab[12][39] , \mult_22/ab[12][40] ,
         \mult_22/ab[12][41] , \mult_22/ab[12][42] , \mult_22/ab[12][43] ,
         \mult_22/ab[12][44] , \mult_22/ab[12][45] , \mult_22/ab[12][46] ,
         \mult_22/ab[12][47] , \mult_22/ab[12][48] , \mult_22/ab[12][49] ,
         \mult_22/ab[12][50] , \mult_22/ab[12][51] , \mult_22/ab[12][52] ,
         \mult_22/ab[12][53] , \mult_22/ab[12][54] , \mult_22/ab[12][55] ,
         \mult_22/ab[12][56] , \mult_22/ab[12][57] , \mult_22/ab[12][58] ,
         \mult_22/ab[12][59] , \mult_22/ab[12][60] , \mult_22/ab[12][61] ,
         \mult_22/ab[12][62] , \mult_22/ab[12][63] , \mult_22/ab[13][0] ,
         \mult_22/ab[13][1] , \mult_22/ab[13][2] , \mult_22/ab[13][3] ,
         \mult_22/ab[13][4] , \mult_22/ab[13][5] , \mult_22/ab[13][6] ,
         \mult_22/ab[13][7] , \mult_22/ab[13][8] , \mult_22/ab[13][9] ,
         \mult_22/ab[13][10] , \mult_22/ab[13][11] , \mult_22/ab[13][12] ,
         \mult_22/ab[13][13] , \mult_22/ab[13][14] , \mult_22/ab[13][15] ,
         \mult_22/ab[13][16] , \mult_22/ab[13][17] , \mult_22/ab[13][18] ,
         \mult_22/ab[13][19] , \mult_22/ab[13][20] , \mult_22/ab[13][21] ,
         \mult_22/ab[13][22] , \mult_22/ab[13][23] , \mult_22/ab[13][24] ,
         \mult_22/ab[13][25] , \mult_22/ab[13][26] , \mult_22/ab[13][27] ,
         \mult_22/ab[13][28] , \mult_22/ab[13][29] , \mult_22/ab[13][30] ,
         \mult_22/ab[13][31] , \mult_22/ab[13][32] , \mult_22/ab[13][33] ,
         \mult_22/ab[13][34] , \mult_22/ab[13][35] , \mult_22/ab[13][36] ,
         \mult_22/ab[13][37] , \mult_22/ab[13][38] , \mult_22/ab[13][39] ,
         \mult_22/ab[13][40] , \mult_22/ab[13][41] , \mult_22/ab[13][42] ,
         \mult_22/ab[13][43] , \mult_22/ab[13][44] , \mult_22/ab[13][45] ,
         \mult_22/ab[13][46] , \mult_22/ab[13][47] , \mult_22/ab[13][48] ,
         \mult_22/ab[13][49] , \mult_22/ab[13][50] , \mult_22/ab[13][51] ,
         \mult_22/ab[13][52] , \mult_22/ab[13][53] , \mult_22/ab[13][54] ,
         \mult_22/ab[13][55] , \mult_22/ab[13][56] , \mult_22/ab[13][57] ,
         \mult_22/ab[13][58] , \mult_22/ab[13][59] , \mult_22/ab[13][60] ,
         \mult_22/ab[13][61] , \mult_22/ab[13][62] , \mult_22/ab[13][63] ,
         \mult_22/ab[14][0] , \mult_22/ab[14][1] , \mult_22/ab[14][2] ,
         \mult_22/ab[14][3] , \mult_22/ab[14][4] , \mult_22/ab[14][5] ,
         \mult_22/ab[14][6] , \mult_22/ab[14][7] , \mult_22/ab[14][8] ,
         \mult_22/ab[14][9] , \mult_22/ab[14][10] , \mult_22/ab[14][11] ,
         \mult_22/ab[14][12] , \mult_22/ab[14][13] , \mult_22/ab[14][14] ,
         \mult_22/ab[14][15] , \mult_22/ab[14][16] , \mult_22/ab[14][17] ,
         \mult_22/ab[14][18] , \mult_22/ab[14][19] , \mult_22/ab[14][20] ,
         \mult_22/ab[14][21] , \mult_22/ab[14][22] , \mult_22/ab[14][23] ,
         \mult_22/ab[14][24] , \mult_22/ab[14][25] , \mult_22/ab[14][26] ,
         \mult_22/ab[14][27] , \mult_22/ab[14][28] , \mult_22/ab[14][29] ,
         \mult_22/ab[14][30] , \mult_22/ab[14][31] , \mult_22/ab[14][32] ,
         \mult_22/ab[14][33] , \mult_22/ab[14][34] , \mult_22/ab[14][35] ,
         \mult_22/ab[14][36] , \mult_22/ab[14][37] , \mult_22/ab[14][38] ,
         \mult_22/ab[14][39] , \mult_22/ab[14][40] , \mult_22/ab[14][41] ,
         \mult_22/ab[14][42] , \mult_22/ab[14][43] , \mult_22/ab[14][44] ,
         \mult_22/ab[14][45] , \mult_22/ab[14][46] , \mult_22/ab[14][47] ,
         \mult_22/ab[14][48] , \mult_22/ab[14][49] , \mult_22/ab[14][50] ,
         \mult_22/ab[14][51] , \mult_22/ab[14][52] , \mult_22/ab[14][53] ,
         \mult_22/ab[14][54] , \mult_22/ab[14][55] , \mult_22/ab[14][56] ,
         \mult_22/ab[14][57] , \mult_22/ab[14][58] , \mult_22/ab[14][59] ,
         \mult_22/ab[14][60] , \mult_22/ab[14][61] , \mult_22/ab[14][62] ,
         \mult_22/ab[14][63] , \mult_22/ab[15][0] , \mult_22/ab[15][1] ,
         \mult_22/ab[15][2] , \mult_22/ab[15][3] , \mult_22/ab[15][4] ,
         \mult_22/ab[15][5] , \mult_22/ab[15][6] , \mult_22/ab[15][7] ,
         \mult_22/ab[15][8] , \mult_22/ab[15][9] , \mult_22/ab[15][10] ,
         \mult_22/ab[15][11] , \mult_22/ab[15][12] , \mult_22/ab[15][13] ,
         \mult_22/ab[15][14] , \mult_22/ab[15][15] , \mult_22/ab[15][16] ,
         \mult_22/ab[15][17] , \mult_22/ab[15][18] , \mult_22/ab[15][19] ,
         \mult_22/ab[15][20] , \mult_22/ab[15][21] , \mult_22/ab[15][22] ,
         \mult_22/ab[15][23] , \mult_22/ab[15][24] , \mult_22/ab[15][25] ,
         \mult_22/ab[15][26] , \mult_22/ab[15][27] , \mult_22/ab[15][28] ,
         \mult_22/ab[15][29] , \mult_22/ab[15][30] , \mult_22/ab[15][31] ,
         \mult_22/ab[15][32] , \mult_22/ab[15][33] , \mult_22/ab[15][34] ,
         \mult_22/ab[15][35] , \mult_22/ab[15][36] , \mult_22/ab[15][37] ,
         \mult_22/ab[15][38] , \mult_22/ab[15][39] , \mult_22/ab[15][40] ,
         \mult_22/ab[15][41] , \mult_22/ab[15][42] , \mult_22/ab[15][43] ,
         \mult_22/ab[15][44] , \mult_22/ab[15][45] , \mult_22/ab[15][46] ,
         \mult_22/ab[15][47] , \mult_22/ab[15][48] , \mult_22/ab[15][49] ,
         \mult_22/ab[15][50] , \mult_22/ab[15][51] , \mult_22/ab[15][52] ,
         \mult_22/ab[15][53] , \mult_22/ab[15][54] , \mult_22/ab[15][55] ,
         \mult_22/ab[15][56] , \mult_22/ab[15][57] , \mult_22/ab[15][58] ,
         \mult_22/ab[15][59] , \mult_22/ab[15][60] , \mult_22/ab[15][61] ,
         \mult_22/ab[15][62] , \mult_22/ab[15][63] , \mult_22/ab[16][0] ,
         \mult_22/ab[16][1] , \mult_22/ab[16][2] , \mult_22/ab[16][3] ,
         \mult_22/ab[16][4] , \mult_22/ab[16][5] , \mult_22/ab[16][6] ,
         \mult_22/ab[16][7] , \mult_22/ab[16][8] , \mult_22/ab[16][9] ,
         \mult_22/ab[16][10] , \mult_22/ab[16][11] , \mult_22/ab[16][12] ,
         \mult_22/ab[16][13] , \mult_22/ab[16][14] , \mult_22/ab[16][15] ,
         \mult_22/ab[16][16] , \mult_22/ab[16][17] , \mult_22/ab[16][18] ,
         \mult_22/ab[16][19] , \mult_22/ab[16][20] , \mult_22/ab[16][21] ,
         \mult_22/ab[16][22] , \mult_22/ab[16][23] , \mult_22/ab[16][24] ,
         \mult_22/ab[16][25] , \mult_22/ab[16][26] , \mult_22/ab[16][27] ,
         \mult_22/ab[16][28] , \mult_22/ab[16][29] , \mult_22/ab[16][30] ,
         \mult_22/ab[16][31] , \mult_22/ab[16][32] , \mult_22/ab[16][33] ,
         \mult_22/ab[16][34] , \mult_22/ab[16][35] , \mult_22/ab[16][36] ,
         \mult_22/ab[16][37] , \mult_22/ab[16][38] , \mult_22/ab[16][39] ,
         \mult_22/ab[16][40] , \mult_22/ab[16][41] , \mult_22/ab[16][42] ,
         \mult_22/ab[16][43] , \mult_22/ab[16][44] , \mult_22/ab[16][45] ,
         \mult_22/ab[16][46] , \mult_22/ab[16][47] , \mult_22/ab[16][48] ,
         \mult_22/ab[16][49] , \mult_22/ab[16][50] , \mult_22/ab[16][51] ,
         \mult_22/ab[16][52] , \mult_22/ab[16][53] , \mult_22/ab[16][54] ,
         \mult_22/ab[16][55] , \mult_22/ab[16][56] , \mult_22/ab[16][57] ,
         \mult_22/ab[16][58] , \mult_22/ab[16][59] , \mult_22/ab[16][60] ,
         \mult_22/ab[16][61] , \mult_22/ab[16][62] , \mult_22/ab[16][63] ,
         \mult_22/ab[17][0] , \mult_22/ab[17][1] , \mult_22/ab[17][2] ,
         \mult_22/ab[17][3] , \mult_22/ab[17][4] , \mult_22/ab[17][5] ,
         \mult_22/ab[17][6] , \mult_22/ab[17][7] , \mult_22/ab[17][8] ,
         \mult_22/ab[17][9] , \mult_22/ab[17][10] , \mult_22/ab[17][11] ,
         \mult_22/ab[17][12] , \mult_22/ab[17][13] , \mult_22/ab[17][14] ,
         \mult_22/ab[17][15] , \mult_22/ab[17][16] , \mult_22/ab[17][17] ,
         \mult_22/ab[17][18] , \mult_22/ab[17][19] , \mult_22/ab[17][20] ,
         \mult_22/ab[17][21] , \mult_22/ab[17][22] , \mult_22/ab[17][23] ,
         \mult_22/ab[17][24] , \mult_22/ab[17][25] , \mult_22/ab[17][26] ,
         \mult_22/ab[17][27] , \mult_22/ab[17][28] , \mult_22/ab[17][29] ,
         \mult_22/ab[17][30] , \mult_22/ab[17][31] , \mult_22/ab[17][32] ,
         \mult_22/ab[17][33] , \mult_22/ab[17][34] , \mult_22/ab[17][35] ,
         \mult_22/ab[17][36] , \mult_22/ab[17][37] , \mult_22/ab[17][38] ,
         \mult_22/ab[17][39] , \mult_22/ab[17][40] , \mult_22/ab[17][41] ,
         \mult_22/ab[17][42] , \mult_22/ab[17][43] , \mult_22/ab[17][44] ,
         \mult_22/ab[17][45] , \mult_22/ab[17][46] , \mult_22/ab[17][47] ,
         \mult_22/ab[17][48] , \mult_22/ab[17][49] , \mult_22/ab[17][50] ,
         \mult_22/ab[17][51] , \mult_22/ab[17][52] , \mult_22/ab[17][53] ,
         \mult_22/ab[17][54] , \mult_22/ab[17][55] , \mult_22/ab[17][56] ,
         \mult_22/ab[17][57] , \mult_22/ab[17][58] , \mult_22/ab[17][59] ,
         \mult_22/ab[17][60] , \mult_22/ab[17][61] , \mult_22/ab[17][62] ,
         \mult_22/ab[17][63] , \mult_22/ab[18][0] , \mult_22/ab[18][1] ,
         \mult_22/ab[18][2] , \mult_22/ab[18][3] , \mult_22/ab[18][4] ,
         \mult_22/ab[18][5] , \mult_22/ab[18][6] , \mult_22/ab[18][7] ,
         \mult_22/ab[18][8] , \mult_22/ab[18][9] , \mult_22/ab[18][10] ,
         \mult_22/ab[18][11] , \mult_22/ab[18][12] , \mult_22/ab[18][13] ,
         \mult_22/ab[18][14] , \mult_22/ab[18][15] , \mult_22/ab[18][16] ,
         \mult_22/ab[18][17] , \mult_22/ab[18][18] , \mult_22/ab[18][19] ,
         \mult_22/ab[18][20] , \mult_22/ab[18][21] , \mult_22/ab[18][22] ,
         \mult_22/ab[18][23] , \mult_22/ab[18][24] , \mult_22/ab[18][25] ,
         \mult_22/ab[18][26] , \mult_22/ab[18][27] , \mult_22/ab[18][28] ,
         \mult_22/ab[18][29] , \mult_22/ab[18][30] , \mult_22/ab[18][31] ,
         \mult_22/ab[18][32] , \mult_22/ab[18][33] , \mult_22/ab[18][34] ,
         \mult_22/ab[18][35] , \mult_22/ab[18][36] , \mult_22/ab[18][37] ,
         \mult_22/ab[18][38] , \mult_22/ab[18][39] , \mult_22/ab[18][41] ,
         \mult_22/ab[18][42] , \mult_22/ab[18][43] , \mult_22/ab[18][44] ,
         \mult_22/ab[18][45] , \mult_22/ab[18][46] , \mult_22/ab[18][47] ,
         \mult_22/ab[18][48] , \mult_22/ab[18][49] , \mult_22/ab[18][50] ,
         \mult_22/ab[18][51] , \mult_22/ab[18][52] , \mult_22/ab[18][53] ,
         \mult_22/ab[18][54] , \mult_22/ab[18][55] , \mult_22/ab[18][56] ,
         \mult_22/ab[18][57] , \mult_22/ab[18][58] , \mult_22/ab[18][59] ,
         \mult_22/ab[18][60] , \mult_22/ab[18][61] , \mult_22/ab[18][62] ,
         \mult_22/ab[18][63] , \mult_22/ab[19][0] , \mult_22/ab[19][1] ,
         \mult_22/ab[19][2] , \mult_22/ab[19][3] , \mult_22/ab[19][4] ,
         \mult_22/ab[19][5] , \mult_22/ab[19][6] , \mult_22/ab[19][7] ,
         \mult_22/ab[19][8] , \mult_22/ab[19][9] , \mult_22/ab[19][10] ,
         \mult_22/ab[19][11] , \mult_22/ab[19][12] , \mult_22/ab[19][13] ,
         \mult_22/ab[19][14] , \mult_22/ab[19][15] , \mult_22/ab[19][16] ,
         \mult_22/ab[19][17] , \mult_22/ab[19][18] , \mult_22/ab[19][19] ,
         \mult_22/ab[19][20] , \mult_22/ab[19][21] , \mult_22/ab[19][22] ,
         \mult_22/ab[19][23] , \mult_22/ab[19][24] , \mult_22/ab[19][25] ,
         \mult_22/ab[19][26] , \mult_22/ab[19][27] , \mult_22/ab[19][28] ,
         \mult_22/ab[19][29] , \mult_22/ab[19][30] , \mult_22/ab[19][31] ,
         \mult_22/ab[19][32] , \mult_22/ab[19][33] , \mult_22/ab[19][34] ,
         \mult_22/ab[19][35] , \mult_22/ab[19][36] , \mult_22/ab[19][37] ,
         \mult_22/ab[19][38] , \mult_22/ab[19][39] , \mult_22/ab[19][40] ,
         \mult_22/ab[19][41] , \mult_22/ab[19][42] , \mult_22/ab[19][43] ,
         \mult_22/ab[19][44] , \mult_22/ab[19][45] , \mult_22/ab[19][46] ,
         \mult_22/ab[19][47] , \mult_22/ab[19][48] , \mult_22/ab[19][49] ,
         \mult_22/ab[19][50] , \mult_22/ab[19][51] , \mult_22/ab[19][52] ,
         \mult_22/ab[19][53] , \mult_22/ab[19][54] , \mult_22/ab[19][55] ,
         \mult_22/ab[19][56] , \mult_22/ab[19][57] , \mult_22/ab[19][58] ,
         \mult_22/ab[19][59] , \mult_22/ab[19][60] , \mult_22/ab[19][61] ,
         \mult_22/ab[19][62] , \mult_22/ab[19][63] , \mult_22/ab[20][0] ,
         \mult_22/ab[20][1] , \mult_22/ab[20][2] , \mult_22/ab[20][3] ,
         \mult_22/ab[20][4] , \mult_22/ab[20][5] , \mult_22/ab[20][6] ,
         \mult_22/ab[20][7] , \mult_22/ab[20][8] , \mult_22/ab[20][9] ,
         \mult_22/ab[20][10] , \mult_22/ab[20][11] , \mult_22/ab[20][12] ,
         \mult_22/ab[20][13] , \mult_22/ab[20][14] , \mult_22/ab[20][15] ,
         \mult_22/ab[20][16] , \mult_22/ab[20][17] , \mult_22/ab[20][18] ,
         \mult_22/ab[20][19] , \mult_22/ab[20][20] , \mult_22/ab[20][21] ,
         \mult_22/ab[20][22] , \mult_22/ab[20][23] , \mult_22/ab[20][24] ,
         \mult_22/ab[20][25] , \mult_22/ab[20][26] , \mult_22/ab[20][27] ,
         \mult_22/ab[20][28] , \mult_22/ab[20][29] , \mult_22/ab[20][30] ,
         \mult_22/ab[20][31] , \mult_22/ab[20][32] , \mult_22/ab[20][33] ,
         \mult_22/ab[20][34] , \mult_22/ab[20][35] , \mult_22/ab[20][36] ,
         \mult_22/ab[20][37] , \mult_22/ab[20][38] , \mult_22/ab[20][39] ,
         \mult_22/ab[20][40] , \mult_22/ab[20][41] , \mult_22/ab[20][42] ,
         \mult_22/ab[20][43] , \mult_22/ab[20][44] , \mult_22/ab[20][45] ,
         \mult_22/ab[20][46] , \mult_22/ab[20][47] , \mult_22/ab[20][48] ,
         \mult_22/ab[20][49] , \mult_22/ab[20][50] , \mult_22/ab[20][51] ,
         \mult_22/ab[20][52] , \mult_22/ab[20][53] , \mult_22/ab[20][54] ,
         \mult_22/ab[20][55] , \mult_22/ab[20][56] , \mult_22/ab[20][57] ,
         \mult_22/ab[20][58] , \mult_22/ab[20][59] , \mult_22/ab[20][60] ,
         \mult_22/ab[20][61] , \mult_22/ab[20][62] , \mult_22/ab[20][63] ,
         \mult_22/ab[21][0] , \mult_22/ab[21][1] , \mult_22/ab[21][2] ,
         \mult_22/ab[21][3] , \mult_22/ab[21][4] , \mult_22/ab[21][5] ,
         \mult_22/ab[21][6] , \mult_22/ab[21][7] , \mult_22/ab[21][8] ,
         \mult_22/ab[21][9] , \mult_22/ab[21][10] , \mult_22/ab[21][11] ,
         \mult_22/ab[21][12] , \mult_22/ab[21][13] , \mult_22/ab[21][14] ,
         \mult_22/ab[21][15] , \mult_22/ab[21][16] , \mult_22/ab[21][17] ,
         \mult_22/ab[21][18] , \mult_22/ab[21][19] , \mult_22/ab[21][20] ,
         \mult_22/ab[21][21] , \mult_22/ab[21][22] , \mult_22/ab[21][23] ,
         \mult_22/ab[21][24] , \mult_22/ab[21][25] , \mult_22/ab[21][26] ,
         \mult_22/ab[21][27] , \mult_22/ab[21][28] , \mult_22/ab[21][29] ,
         \mult_22/ab[21][30] , \mult_22/ab[21][31] , \mult_22/ab[21][32] ,
         \mult_22/ab[21][33] , \mult_22/ab[21][34] , \mult_22/ab[21][35] ,
         \mult_22/ab[21][37] , \mult_22/ab[21][39] , \mult_22/ab[21][40] ,
         \mult_22/ab[21][41] , \mult_22/ab[21][42] , \mult_22/ab[21][43] ,
         \mult_22/ab[21][44] , \mult_22/ab[21][45] , \mult_22/ab[21][46] ,
         \mult_22/ab[21][47] , \mult_22/ab[21][48] , \mult_22/ab[21][49] ,
         \mult_22/ab[21][50] , \mult_22/ab[21][51] , \mult_22/ab[21][52] ,
         \mult_22/ab[21][53] , \mult_22/ab[21][54] , \mult_22/ab[21][55] ,
         \mult_22/ab[21][56] , \mult_22/ab[21][57] , \mult_22/ab[21][58] ,
         \mult_22/ab[21][59] , \mult_22/ab[21][60] , \mult_22/ab[21][61] ,
         \mult_22/ab[21][62] , \mult_22/ab[21][63] , \mult_22/ab[22][0] ,
         \mult_22/ab[22][1] , \mult_22/ab[22][2] , \mult_22/ab[22][3] ,
         \mult_22/ab[22][4] , \mult_22/ab[22][5] , \mult_22/ab[22][6] ,
         \mult_22/ab[22][7] , \mult_22/ab[22][8] , \mult_22/ab[22][9] ,
         \mult_22/ab[22][10] , \mult_22/ab[22][11] , \mult_22/ab[22][12] ,
         \mult_22/ab[22][13] , \mult_22/ab[22][14] , \mult_22/ab[22][15] ,
         \mult_22/ab[22][16] , \mult_22/ab[22][17] , \mult_22/ab[22][18] ,
         \mult_22/ab[22][19] , \mult_22/ab[22][20] , \mult_22/ab[22][21] ,
         \mult_22/ab[22][22] , \mult_22/ab[22][23] , \mult_22/ab[22][24] ,
         \mult_22/ab[22][25] , \mult_22/ab[22][26] , \mult_22/ab[22][27] ,
         \mult_22/ab[22][28] , \mult_22/ab[22][29] , \mult_22/ab[22][30] ,
         \mult_22/ab[22][31] , \mult_22/ab[22][32] , \mult_22/ab[22][33] ,
         \mult_22/ab[22][34] , \mult_22/ab[22][35] , \mult_22/ab[22][36] ,
         \mult_22/ab[22][37] , \mult_22/ab[22][39] , \mult_22/ab[22][40] ,
         \mult_22/ab[22][41] , \mult_22/ab[22][42] , \mult_22/ab[22][43] ,
         \mult_22/ab[22][44] , \mult_22/ab[22][45] , \mult_22/ab[22][46] ,
         \mult_22/ab[22][47] , \mult_22/ab[22][48] , \mult_22/ab[22][49] ,
         \mult_22/ab[22][50] , \mult_22/ab[22][51] , \mult_22/ab[22][52] ,
         \mult_22/ab[22][53] , \mult_22/ab[22][54] , \mult_22/ab[22][55] ,
         \mult_22/ab[22][56] , \mult_22/ab[22][57] , \mult_22/ab[22][58] ,
         \mult_22/ab[22][59] , \mult_22/ab[22][60] , \mult_22/ab[22][61] ,
         \mult_22/ab[22][62] , \mult_22/ab[22][63] , \mult_22/ab[23][0] ,
         \mult_22/ab[23][1] , \mult_22/ab[23][2] , \mult_22/ab[23][3] ,
         \mult_22/ab[23][4] , \mult_22/ab[23][5] , \mult_22/ab[23][6] ,
         \mult_22/ab[23][7] , \mult_22/ab[23][8] , \mult_22/ab[23][9] ,
         \mult_22/ab[23][10] , \mult_22/ab[23][11] , \mult_22/ab[23][12] ,
         \mult_22/ab[23][13] , \mult_22/ab[23][14] , \mult_22/ab[23][15] ,
         \mult_22/ab[23][16] , \mult_22/ab[23][17] , \mult_22/ab[23][18] ,
         \mult_22/ab[23][19] , \mult_22/ab[23][20] , \mult_22/ab[23][21] ,
         \mult_22/ab[23][22] , \mult_22/ab[23][23] , \mult_22/ab[23][24] ,
         \mult_22/ab[23][25] , \mult_22/ab[23][26] , \mult_22/ab[23][27] ,
         \mult_22/ab[23][28] , \mult_22/ab[23][29] , \mult_22/ab[23][30] ,
         \mult_22/ab[23][31] , \mult_22/ab[23][32] , \mult_22/ab[23][33] ,
         \mult_22/ab[23][34] , \mult_22/ab[23][35] , \mult_22/ab[23][36] ,
         \mult_22/ab[23][38] , \mult_22/ab[23][39] , \mult_22/ab[23][40] ,
         \mult_22/ab[23][41] , \mult_22/ab[23][42] , \mult_22/ab[23][43] ,
         \mult_22/ab[23][44] , \mult_22/ab[23][45] , \mult_22/ab[23][46] ,
         \mult_22/ab[23][47] , \mult_22/ab[23][48] , \mult_22/ab[23][49] ,
         \mult_22/ab[23][50] , \mult_22/ab[23][51] , \mult_22/ab[23][52] ,
         \mult_22/ab[23][53] , \mult_22/ab[23][54] , \mult_22/ab[23][55] ,
         \mult_22/ab[23][56] , \mult_22/ab[23][57] , \mult_22/ab[23][58] ,
         \mult_22/ab[23][59] , \mult_22/ab[23][60] , \mult_22/ab[23][61] ,
         \mult_22/ab[23][62] , \mult_22/ab[23][63] , \mult_22/ab[24][0] ,
         \mult_22/ab[24][1] , \mult_22/ab[24][2] , \mult_22/ab[24][3] ,
         \mult_22/ab[24][4] , \mult_22/ab[24][5] , \mult_22/ab[24][6] ,
         \mult_22/ab[24][7] , \mult_22/ab[24][8] , \mult_22/ab[24][9] ,
         \mult_22/ab[24][10] , \mult_22/ab[24][11] , \mult_22/ab[24][12] ,
         \mult_22/ab[24][13] , \mult_22/ab[24][14] , \mult_22/ab[24][15] ,
         \mult_22/ab[24][16] , \mult_22/ab[24][17] , \mult_22/ab[24][18] ,
         \mult_22/ab[24][19] , \mult_22/ab[24][20] , \mult_22/ab[24][21] ,
         \mult_22/ab[24][22] , \mult_22/ab[24][23] , \mult_22/ab[24][24] ,
         \mult_22/ab[24][25] , \mult_22/ab[24][26] , \mult_22/ab[24][27] ,
         \mult_22/ab[24][28] , \mult_22/ab[24][29] , \mult_22/ab[24][30] ,
         \mult_22/ab[24][31] , \mult_22/ab[24][33] , \mult_22/ab[24][34] ,
         \mult_22/ab[24][35] , \mult_22/ab[24][36] , \mult_22/ab[24][37] ,
         \mult_22/ab[24][38] , \mult_22/ab[24][39] , \mult_22/ab[24][40] ,
         \mult_22/ab[24][41] , \mult_22/ab[24][42] , \mult_22/ab[24][43] ,
         \mult_22/ab[24][44] , \mult_22/ab[24][45] , \mult_22/ab[24][46] ,
         \mult_22/ab[24][47] , \mult_22/ab[24][48] , \mult_22/ab[24][49] ,
         \mult_22/ab[24][50] , \mult_22/ab[24][51] , \mult_22/ab[24][52] ,
         \mult_22/ab[24][53] , \mult_22/ab[24][54] , \mult_22/ab[24][55] ,
         \mult_22/ab[24][56] , \mult_22/ab[24][57] , \mult_22/ab[24][58] ,
         \mult_22/ab[24][59] , \mult_22/ab[24][60] , \mult_22/ab[24][61] ,
         \mult_22/ab[24][62] , \mult_22/ab[24][63] , \mult_22/ab[25][0] ,
         \mult_22/ab[25][1] , \mult_22/ab[25][2] , \mult_22/ab[25][3] ,
         \mult_22/ab[25][4] , \mult_22/ab[25][5] , \mult_22/ab[25][6] ,
         \mult_22/ab[25][7] , \mult_22/ab[25][8] , \mult_22/ab[25][9] ,
         \mult_22/ab[25][10] , \mult_22/ab[25][11] , \mult_22/ab[25][12] ,
         \mult_22/ab[25][13] , \mult_22/ab[25][14] , \mult_22/ab[25][15] ,
         \mult_22/ab[25][16] , \mult_22/ab[25][17] , \mult_22/ab[25][18] ,
         \mult_22/ab[25][19] , \mult_22/ab[25][20] , \mult_22/ab[25][21] ,
         \mult_22/ab[25][22] , \mult_22/ab[25][23] , \mult_22/ab[25][24] ,
         \mult_22/ab[25][25] , \mult_22/ab[25][26] , \mult_22/ab[25][27] ,
         \mult_22/ab[25][28] , \mult_22/ab[25][29] , \mult_22/ab[25][30] ,
         \mult_22/ab[25][31] , \mult_22/ab[25][32] , \mult_22/ab[25][33] ,
         \mult_22/ab[25][34] , \mult_22/ab[25][36] , \mult_22/ab[25][37] ,
         \mult_22/ab[25][38] , \mult_22/ab[25][39] , \mult_22/ab[25][40] ,
         \mult_22/ab[25][41] , \mult_22/ab[25][42] , \mult_22/ab[25][43] ,
         \mult_22/ab[25][44] , \mult_22/ab[25][45] , \mult_22/ab[25][46] ,
         \mult_22/ab[25][47] , \mult_22/ab[25][48] , \mult_22/ab[25][49] ,
         \mult_22/ab[25][50] , \mult_22/ab[25][51] , \mult_22/ab[25][52] ,
         \mult_22/ab[25][53] , \mult_22/ab[25][54] , \mult_22/ab[25][55] ,
         \mult_22/ab[25][56] , \mult_22/ab[25][57] , \mult_22/ab[25][58] ,
         \mult_22/ab[25][59] , \mult_22/ab[25][60] , \mult_22/ab[25][61] ,
         \mult_22/ab[25][62] , \mult_22/ab[25][63] , \mult_22/ab[26][0] ,
         \mult_22/ab[26][1] , \mult_22/ab[26][2] , \mult_22/ab[26][3] ,
         \mult_22/ab[26][4] , \mult_22/ab[26][5] , \mult_22/ab[26][6] ,
         \mult_22/ab[26][7] , \mult_22/ab[26][8] , \mult_22/ab[26][9] ,
         \mult_22/ab[26][10] , \mult_22/ab[26][11] , \mult_22/ab[26][12] ,
         \mult_22/ab[26][13] , \mult_22/ab[26][14] , \mult_22/ab[26][15] ,
         \mult_22/ab[26][16] , \mult_22/ab[26][17] , \mult_22/ab[26][18] ,
         \mult_22/ab[26][19] , \mult_22/ab[26][20] , \mult_22/ab[26][21] ,
         \mult_22/ab[26][22] , \mult_22/ab[26][23] , \mult_22/ab[26][24] ,
         \mult_22/ab[26][25] , \mult_22/ab[26][26] , \mult_22/ab[26][27] ,
         \mult_22/ab[26][28] , \mult_22/ab[26][29] , \mult_22/ab[26][30] ,
         \mult_22/ab[26][31] , \mult_22/ab[26][32] , \mult_22/ab[26][33] ,
         \mult_22/ab[26][36] , \mult_22/ab[26][37] , \mult_22/ab[26][38] ,
         \mult_22/ab[26][39] , \mult_22/ab[26][40] , \mult_22/ab[26][41] ,
         \mult_22/ab[26][42] , \mult_22/ab[26][43] , \mult_22/ab[26][44] ,
         \mult_22/ab[26][45] , \mult_22/ab[26][46] , \mult_22/ab[26][47] ,
         \mult_22/ab[26][48] , \mult_22/ab[26][49] , \mult_22/ab[26][50] ,
         \mult_22/ab[26][51] , \mult_22/ab[26][52] , \mult_22/ab[26][53] ,
         \mult_22/ab[26][54] , \mult_22/ab[26][55] , \mult_22/ab[26][56] ,
         \mult_22/ab[26][57] , \mult_22/ab[26][58] , \mult_22/ab[26][59] ,
         \mult_22/ab[26][60] , \mult_22/ab[26][61] , \mult_22/ab[26][62] ,
         \mult_22/ab[26][63] , \mult_22/ab[27][0] , \mult_22/ab[27][1] ,
         \mult_22/ab[27][2] , \mult_22/ab[27][3] , \mult_22/ab[27][4] ,
         \mult_22/ab[27][5] , \mult_22/ab[27][6] , \mult_22/ab[27][7] ,
         \mult_22/ab[27][8] , \mult_22/ab[27][9] , \mult_22/ab[27][10] ,
         \mult_22/ab[27][11] , \mult_22/ab[27][12] , \mult_22/ab[27][13] ,
         \mult_22/ab[27][14] , \mult_22/ab[27][15] , \mult_22/ab[27][16] ,
         \mult_22/ab[27][17] , \mult_22/ab[27][18] , \mult_22/ab[27][19] ,
         \mult_22/ab[27][20] , \mult_22/ab[27][21] , \mult_22/ab[27][22] ,
         \mult_22/ab[27][23] , \mult_22/ab[27][24] , \mult_22/ab[27][25] ,
         \mult_22/ab[27][26] , \mult_22/ab[27][27] , \mult_22/ab[27][28] ,
         \mult_22/ab[27][29] , \mult_22/ab[27][30] , \mult_22/ab[27][31] ,
         \mult_22/ab[27][32] , \mult_22/ab[27][33] , \mult_22/ab[27][34] ,
         \mult_22/ab[27][35] , \mult_22/ab[27][36] , \mult_22/ab[27][37] ,
         \mult_22/ab[27][38] , \mult_22/ab[27][39] , \mult_22/ab[27][40] ,
         \mult_22/ab[27][41] , \mult_22/ab[27][42] , \mult_22/ab[27][43] ,
         \mult_22/ab[27][44] , \mult_22/ab[27][45] , \mult_22/ab[27][46] ,
         \mult_22/ab[27][47] , \mult_22/ab[27][48] , \mult_22/ab[27][49] ,
         \mult_22/ab[27][50] , \mult_22/ab[27][51] , \mult_22/ab[27][52] ,
         \mult_22/ab[27][53] , \mult_22/ab[27][54] , \mult_22/ab[27][55] ,
         \mult_22/ab[27][56] , \mult_22/ab[27][57] , \mult_22/ab[27][58] ,
         \mult_22/ab[27][59] , \mult_22/ab[27][60] , \mult_22/ab[27][61] ,
         \mult_22/ab[27][62] , \mult_22/ab[27][63] , \mult_22/ab[28][0] ,
         \mult_22/ab[28][1] , \mult_22/ab[28][2] , \mult_22/ab[28][3] ,
         \mult_22/ab[28][4] , \mult_22/ab[28][5] , \mult_22/ab[28][6] ,
         \mult_22/ab[28][7] , \mult_22/ab[28][8] , \mult_22/ab[28][9] ,
         \mult_22/ab[28][10] , \mult_22/ab[28][11] , \mult_22/ab[28][12] ,
         \mult_22/ab[28][13] , \mult_22/ab[28][14] , \mult_22/ab[28][15] ,
         \mult_22/ab[28][16] , \mult_22/ab[28][17] , \mult_22/ab[28][18] ,
         \mult_22/ab[28][19] , \mult_22/ab[28][20] , \mult_22/ab[28][21] ,
         \mult_22/ab[28][22] , \mult_22/ab[28][23] , \mult_22/ab[28][24] ,
         \mult_22/ab[28][25] , \mult_22/ab[28][26] , \mult_22/ab[28][27] ,
         \mult_22/ab[28][28] , \mult_22/ab[28][29] , \mult_22/ab[28][31] ,
         \mult_22/ab[28][32] , \mult_22/ab[28][33] , \mult_22/ab[28][34] ,
         \mult_22/ab[28][35] , \mult_22/ab[28][36] , \mult_22/ab[28][37] ,
         \mult_22/ab[28][38] , \mult_22/ab[28][39] , \mult_22/ab[28][40] ,
         \mult_22/ab[28][41] , \mult_22/ab[28][42] , \mult_22/ab[28][43] ,
         \mult_22/ab[28][44] , \mult_22/ab[28][45] , \mult_22/ab[28][46] ,
         \mult_22/ab[28][47] , \mult_22/ab[28][48] , \mult_22/ab[28][49] ,
         \mult_22/ab[28][50] , \mult_22/ab[28][51] , \mult_22/ab[28][52] ,
         \mult_22/ab[28][53] , \mult_22/ab[28][54] , \mult_22/ab[28][55] ,
         \mult_22/ab[28][56] , \mult_22/ab[28][57] , \mult_22/ab[28][58] ,
         \mult_22/ab[28][59] , \mult_22/ab[28][60] , \mult_22/ab[28][61] ,
         \mult_22/ab[28][62] , \mult_22/ab[28][63] , \mult_22/ab[29][0] ,
         \mult_22/ab[29][1] , \mult_22/ab[29][2] , \mult_22/ab[29][3] ,
         \mult_22/ab[29][4] , \mult_22/ab[29][5] , \mult_22/ab[29][6] ,
         \mult_22/ab[29][7] , \mult_22/ab[29][8] , \mult_22/ab[29][9] ,
         \mult_22/ab[29][10] , \mult_22/ab[29][11] , \mult_22/ab[29][12] ,
         \mult_22/ab[29][13] , \mult_22/ab[29][14] , \mult_22/ab[29][15] ,
         \mult_22/ab[29][16] , \mult_22/ab[29][17] , \mult_22/ab[29][18] ,
         \mult_22/ab[29][19] , \mult_22/ab[29][20] , \mult_22/ab[29][21] ,
         \mult_22/ab[29][22] , \mult_22/ab[29][23] , \mult_22/ab[29][24] ,
         \mult_22/ab[29][25] , \mult_22/ab[29][26] , \mult_22/ab[29][27] ,
         \mult_22/ab[29][28] , \mult_22/ab[29][29] , \mult_22/ab[29][30] ,
         \mult_22/ab[29][31] , \mult_22/ab[29][32] , \mult_22/ab[29][33] ,
         \mult_22/ab[29][34] , \mult_22/ab[29][35] , \mult_22/ab[29][36] ,
         \mult_22/ab[29][37] , \mult_22/ab[29][38] , \mult_22/ab[29][39] ,
         \mult_22/ab[29][40] , \mult_22/ab[29][41] , \mult_22/ab[29][42] ,
         \mult_22/ab[29][43] , \mult_22/ab[29][44] , \mult_22/ab[29][45] ,
         \mult_22/ab[29][46] , \mult_22/ab[29][47] , \mult_22/ab[29][48] ,
         \mult_22/ab[29][49] , \mult_22/ab[29][50] , \mult_22/ab[29][51] ,
         \mult_22/ab[29][52] , \mult_22/ab[29][53] , \mult_22/ab[29][54] ,
         \mult_22/ab[29][55] , \mult_22/ab[29][56] , \mult_22/ab[29][57] ,
         \mult_22/ab[29][58] , \mult_22/ab[29][59] , \mult_22/ab[29][60] ,
         \mult_22/ab[29][61] , \mult_22/ab[29][62] , \mult_22/ab[29][63] ,
         \mult_22/ab[30][0] , \mult_22/ab[30][1] , \mult_22/ab[30][2] ,
         \mult_22/ab[30][3] , \mult_22/ab[30][4] , \mult_22/ab[30][5] ,
         \mult_22/ab[30][6] , \mult_22/ab[30][7] , \mult_22/ab[30][8] ,
         \mult_22/ab[30][9] , \mult_22/ab[30][10] , \mult_22/ab[30][11] ,
         \mult_22/ab[30][12] , \mult_22/ab[30][13] , \mult_22/ab[30][14] ,
         \mult_22/ab[30][15] , \mult_22/ab[30][16] , \mult_22/ab[30][17] ,
         \mult_22/ab[30][18] , \mult_22/ab[30][19] , \mult_22/ab[30][20] ,
         \mult_22/ab[30][21] , \mult_22/ab[30][22] , \mult_22/ab[30][23] ,
         \mult_22/ab[30][24] , \mult_22/ab[30][25] , \mult_22/ab[30][26] ,
         \mult_22/ab[30][27] , \mult_22/ab[30][28] , \mult_22/ab[30][29] ,
         \mult_22/ab[30][30] , \mult_22/ab[30][31] , \mult_22/ab[30][32] ,
         \mult_22/ab[30][33] , \mult_22/ab[30][34] , \mult_22/ab[30][35] ,
         \mult_22/ab[30][36] , \mult_22/ab[30][37] , \mult_22/ab[30][38] ,
         \mult_22/ab[30][39] , \mult_22/ab[30][40] , \mult_22/ab[30][41] ,
         \mult_22/ab[30][42] , \mult_22/ab[30][43] , \mult_22/ab[30][44] ,
         \mult_22/ab[30][45] , \mult_22/ab[30][46] , \mult_22/ab[30][47] ,
         \mult_22/ab[30][48] , \mult_22/ab[30][49] , \mult_22/ab[30][50] ,
         \mult_22/ab[30][51] , \mult_22/ab[30][52] , \mult_22/ab[30][53] ,
         \mult_22/ab[30][54] , \mult_22/ab[30][55] , \mult_22/ab[30][56] ,
         \mult_22/ab[30][57] , \mult_22/ab[30][58] , \mult_22/ab[30][59] ,
         \mult_22/ab[30][60] , \mult_22/ab[30][61] , \mult_22/ab[30][62] ,
         \mult_22/ab[30][63] , \mult_22/ab[31][0] , \mult_22/ab[31][1] ,
         \mult_22/ab[31][2] , \mult_22/ab[31][3] , \mult_22/ab[31][4] ,
         \mult_22/ab[31][5] , \mult_22/ab[31][6] , \mult_22/ab[31][7] ,
         \mult_22/ab[31][8] , \mult_22/ab[31][9] , \mult_22/ab[31][10] ,
         \mult_22/ab[31][11] , \mult_22/ab[31][12] , \mult_22/ab[31][13] ,
         \mult_22/ab[31][14] , \mult_22/ab[31][15] , \mult_22/ab[31][16] ,
         \mult_22/ab[31][17] , \mult_22/ab[31][18] , \mult_22/ab[31][19] ,
         \mult_22/ab[31][20] , \mult_22/ab[31][21] , \mult_22/ab[31][22] ,
         \mult_22/ab[31][23] , \mult_22/ab[31][24] , \mult_22/ab[31][25] ,
         \mult_22/ab[31][26] , \mult_22/ab[31][27] , \mult_22/ab[31][28] ,
         \mult_22/ab[31][29] , \mult_22/ab[31][30] , \mult_22/ab[31][31] ,
         \mult_22/ab[31][32] , \mult_22/ab[31][33] , \mult_22/ab[31][34] ,
         \mult_22/ab[31][35] , \mult_22/ab[31][36] , \mult_22/ab[31][37] ,
         \mult_22/ab[31][38] , \mult_22/ab[31][39] , \mult_22/ab[31][40] ,
         \mult_22/ab[31][41] , \mult_22/ab[31][42] , \mult_22/ab[31][43] ,
         \mult_22/ab[31][44] , \mult_22/ab[31][45] , \mult_22/ab[31][46] ,
         \mult_22/ab[31][47] , \mult_22/ab[31][48] , \mult_22/ab[31][49] ,
         \mult_22/ab[31][50] , \mult_22/ab[31][51] , \mult_22/ab[31][52] ,
         \mult_22/ab[31][53] , \mult_22/ab[31][54] , \mult_22/ab[31][55] ,
         \mult_22/ab[31][56] , \mult_22/ab[31][57] , \mult_22/ab[31][58] ,
         \mult_22/ab[31][59] , \mult_22/ab[31][60] , \mult_22/ab[31][61] ,
         \mult_22/ab[31][62] , \mult_22/ab[31][63] , \mult_22/ab[32][0] ,
         \mult_22/ab[32][1] , \mult_22/ab[32][2] , \mult_22/ab[32][3] ,
         \mult_22/ab[32][4] , \mult_22/ab[32][5] , \mult_22/ab[32][6] ,
         \mult_22/ab[32][7] , \mult_22/ab[32][8] , \mult_22/ab[32][9] ,
         \mult_22/ab[32][10] , \mult_22/ab[32][11] , \mult_22/ab[32][12] ,
         \mult_22/ab[32][13] , \mult_22/ab[32][14] , \mult_22/ab[32][15] ,
         \mult_22/ab[32][16] , \mult_22/ab[32][17] , \mult_22/ab[32][18] ,
         \mult_22/ab[32][19] , \mult_22/ab[32][20] , \mult_22/ab[32][21] ,
         \mult_22/ab[32][22] , \mult_22/ab[32][23] , \mult_22/ab[32][24] ,
         \mult_22/ab[32][25] , \mult_22/ab[32][26] , \mult_22/ab[32][27] ,
         \mult_22/ab[32][28] , \mult_22/ab[32][29] , \mult_22/ab[32][30] ,
         \mult_22/ab[32][31] , \mult_22/ab[32][32] , \mult_22/ab[32][33] ,
         \mult_22/ab[32][34] , \mult_22/ab[32][35] , \mult_22/ab[32][36] ,
         \mult_22/ab[32][37] , \mult_22/ab[32][38] , \mult_22/ab[32][39] ,
         \mult_22/ab[32][40] , \mult_22/ab[32][41] , \mult_22/ab[32][42] ,
         \mult_22/ab[32][43] , \mult_22/ab[32][44] , \mult_22/ab[32][45] ,
         \mult_22/ab[32][46] , \mult_22/ab[32][47] , \mult_22/ab[32][48] ,
         \mult_22/ab[32][49] , \mult_22/ab[32][50] , \mult_22/ab[32][51] ,
         \mult_22/ab[32][52] , \mult_22/ab[32][53] , \mult_22/ab[32][54] ,
         \mult_22/ab[32][55] , \mult_22/ab[32][56] , \mult_22/ab[32][57] ,
         \mult_22/ab[32][58] , \mult_22/ab[32][59] , \mult_22/ab[32][60] ,
         \mult_22/ab[32][61] , \mult_22/ab[32][62] , \mult_22/ab[32][63] ,
         \mult_22/ab[33][0] , \mult_22/ab[33][1] , \mult_22/ab[33][2] ,
         \mult_22/ab[33][3] , \mult_22/ab[33][4] , \mult_22/ab[33][5] ,
         \mult_22/ab[33][6] , \mult_22/ab[33][7] , \mult_22/ab[33][8] ,
         \mult_22/ab[33][9] , \mult_22/ab[33][10] , \mult_22/ab[33][11] ,
         \mult_22/ab[33][12] , \mult_22/ab[33][13] , \mult_22/ab[33][14] ,
         \mult_22/ab[33][15] , \mult_22/ab[33][16] , \mult_22/ab[33][17] ,
         \mult_22/ab[33][18] , \mult_22/ab[33][19] , \mult_22/ab[33][20] ,
         \mult_22/ab[33][21] , \mult_22/ab[33][22] , \mult_22/ab[33][23] ,
         \mult_22/ab[33][24] , \mult_22/ab[33][25] , \mult_22/ab[33][26] ,
         \mult_22/ab[33][27] , \mult_22/ab[33][29] , \mult_22/ab[33][30] ,
         \mult_22/ab[33][31] , \mult_22/ab[33][32] , \mult_22/ab[33][33] ,
         \mult_22/ab[33][34] , \mult_22/ab[33][35] , \mult_22/ab[33][36] ,
         \mult_22/ab[33][37] , \mult_22/ab[33][38] , \mult_22/ab[33][39] ,
         \mult_22/ab[33][40] , \mult_22/ab[33][41] , \mult_22/ab[33][42] ,
         \mult_22/ab[33][43] , \mult_22/ab[33][44] , \mult_22/ab[33][45] ,
         \mult_22/ab[33][46] , \mult_22/ab[33][47] , \mult_22/ab[33][48] ,
         \mult_22/ab[33][49] , \mult_22/ab[33][50] , \mult_22/ab[33][51] ,
         \mult_22/ab[33][52] , \mult_22/ab[33][53] , \mult_22/ab[33][54] ,
         \mult_22/ab[33][55] , \mult_22/ab[33][56] , \mult_22/ab[33][57] ,
         \mult_22/ab[33][58] , \mult_22/ab[33][59] , \mult_22/ab[33][60] ,
         \mult_22/ab[33][61] , \mult_22/ab[33][62] , \mult_22/ab[33][63] ,
         \mult_22/ab[34][0] , \mult_22/ab[34][1] , \mult_22/ab[34][2] ,
         \mult_22/ab[34][3] , \mult_22/ab[34][4] , \mult_22/ab[34][5] ,
         \mult_22/ab[34][6] , \mult_22/ab[34][7] , \mult_22/ab[34][8] ,
         \mult_22/ab[34][9] , \mult_22/ab[34][10] , \mult_22/ab[34][11] ,
         \mult_22/ab[34][12] , \mult_22/ab[34][13] , \mult_22/ab[34][14] ,
         \mult_22/ab[34][15] , \mult_22/ab[34][16] , \mult_22/ab[34][17] ,
         \mult_22/ab[34][18] , \mult_22/ab[34][19] , \mult_22/ab[34][20] ,
         \mult_22/ab[34][21] , \mult_22/ab[34][22] , \mult_22/ab[34][23] ,
         \mult_22/ab[34][24] , \mult_22/ab[34][25] , \mult_22/ab[34][26] ,
         \mult_22/ab[34][27] , \mult_22/ab[34][28] , \mult_22/ab[34][29] ,
         \mult_22/ab[34][30] , \mult_22/ab[34][31] , \mult_22/ab[34][32] ,
         \mult_22/ab[34][33] , \mult_22/ab[34][34] , \mult_22/ab[34][35] ,
         \mult_22/ab[34][36] , \mult_22/ab[34][37] , \mult_22/ab[34][38] ,
         \mult_22/ab[34][39] , \mult_22/ab[34][40] , \mult_22/ab[34][41] ,
         \mult_22/ab[34][42] , \mult_22/ab[34][43] , \mult_22/ab[34][44] ,
         \mult_22/ab[34][45] , \mult_22/ab[34][46] , \mult_22/ab[34][47] ,
         \mult_22/ab[34][48] , \mult_22/ab[34][49] , \mult_22/ab[34][50] ,
         \mult_22/ab[34][51] , \mult_22/ab[34][52] , \mult_22/ab[34][53] ,
         \mult_22/ab[34][54] , \mult_22/ab[34][55] , \mult_22/ab[34][56] ,
         \mult_22/ab[34][57] , \mult_22/ab[34][58] , \mult_22/ab[34][59] ,
         \mult_22/ab[34][60] , \mult_22/ab[34][61] , \mult_22/ab[34][62] ,
         \mult_22/ab[34][63] , \mult_22/ab[35][0] , \mult_22/ab[35][1] ,
         \mult_22/ab[35][2] , \mult_22/ab[35][3] , \mult_22/ab[35][4] ,
         \mult_22/ab[35][5] , \mult_22/ab[35][6] , \mult_22/ab[35][7] ,
         \mult_22/ab[35][8] , \mult_22/ab[35][9] , \mult_22/ab[35][10] ,
         \mult_22/ab[35][11] , \mult_22/ab[35][12] , \mult_22/ab[35][13] ,
         \mult_22/ab[35][14] , \mult_22/ab[35][15] , \mult_22/ab[35][16] ,
         \mult_22/ab[35][17] , \mult_22/ab[35][18] , \mult_22/ab[35][19] ,
         \mult_22/ab[35][20] , \mult_22/ab[35][21] , \mult_22/ab[35][22] ,
         \mult_22/ab[35][23] , \mult_22/ab[35][24] , \mult_22/ab[35][25] ,
         \mult_22/ab[35][26] , \mult_22/ab[35][27] , \mult_22/ab[35][28] ,
         \mult_22/ab[35][29] , \mult_22/ab[35][30] , \mult_22/ab[35][31] ,
         \mult_22/ab[35][32] , \mult_22/ab[35][33] , \mult_22/ab[35][34] ,
         \mult_22/ab[35][35] , \mult_22/ab[35][36] , \mult_22/ab[35][37] ,
         \mult_22/ab[35][38] , \mult_22/ab[35][39] , \mult_22/ab[35][40] ,
         \mult_22/ab[35][41] , \mult_22/ab[35][42] , \mult_22/ab[35][43] ,
         \mult_22/ab[35][44] , \mult_22/ab[35][45] , \mult_22/ab[35][46] ,
         \mult_22/ab[35][47] , \mult_22/ab[35][48] , \mult_22/ab[35][49] ,
         \mult_22/ab[35][50] , \mult_22/ab[35][51] , \mult_22/ab[35][52] ,
         \mult_22/ab[35][53] , \mult_22/ab[35][54] , \mult_22/ab[35][55] ,
         \mult_22/ab[35][56] , \mult_22/ab[35][57] , \mult_22/ab[35][58] ,
         \mult_22/ab[35][59] , \mult_22/ab[35][60] , \mult_22/ab[35][61] ,
         \mult_22/ab[35][62] , \mult_22/ab[35][63] , \mult_22/ab[36][0] ,
         \mult_22/ab[36][1] , \mult_22/ab[36][2] , \mult_22/ab[36][3] ,
         \mult_22/ab[36][4] , \mult_22/ab[36][5] , \mult_22/ab[36][6] ,
         \mult_22/ab[36][7] , \mult_22/ab[36][8] , \mult_22/ab[36][9] ,
         \mult_22/ab[36][10] , \mult_22/ab[36][11] , \mult_22/ab[36][12] ,
         \mult_22/ab[36][13] , \mult_22/ab[36][14] , \mult_22/ab[36][15] ,
         \mult_22/ab[36][16] , \mult_22/ab[36][17] , \mult_22/ab[36][18] ,
         \mult_22/ab[36][19] , \mult_22/ab[36][20] , \mult_22/ab[36][21] ,
         \mult_22/ab[36][22] , \mult_22/ab[36][23] , \mult_22/ab[36][24] ,
         \mult_22/ab[36][25] , \mult_22/ab[36][26] , \mult_22/ab[36][27] ,
         \mult_22/ab[36][28] , \mult_22/ab[36][29] , \mult_22/ab[36][30] ,
         \mult_22/ab[36][31] , \mult_22/ab[36][32] , \mult_22/ab[36][33] ,
         \mult_22/ab[36][34] , \mult_22/ab[36][35] , \mult_22/ab[36][36] ,
         \mult_22/ab[36][37] , \mult_22/ab[36][38] , \mult_22/ab[36][39] ,
         \mult_22/ab[36][40] , \mult_22/ab[36][41] , \mult_22/ab[36][42] ,
         \mult_22/ab[36][43] , \mult_22/ab[36][44] , \mult_22/ab[36][45] ,
         \mult_22/ab[36][46] , \mult_22/ab[36][47] , \mult_22/ab[36][48] ,
         \mult_22/ab[36][49] , \mult_22/ab[36][50] , \mult_22/ab[36][51] ,
         \mult_22/ab[36][52] , \mult_22/ab[36][53] , \mult_22/ab[36][54] ,
         \mult_22/ab[36][55] , \mult_22/ab[36][56] , \mult_22/ab[36][57] ,
         \mult_22/ab[36][58] , \mult_22/ab[36][59] , \mult_22/ab[36][60] ,
         \mult_22/ab[36][61] , \mult_22/ab[36][62] , \mult_22/ab[36][63] ,
         \mult_22/ab[37][0] , \mult_22/ab[37][1] , \mult_22/ab[37][2] ,
         \mult_22/ab[37][3] , \mult_22/ab[37][4] , \mult_22/ab[37][5] ,
         \mult_22/ab[37][6] , \mult_22/ab[37][7] , \mult_22/ab[37][8] ,
         \mult_22/ab[37][9] , \mult_22/ab[37][10] , \mult_22/ab[37][11] ,
         \mult_22/ab[37][12] , \mult_22/ab[37][13] , \mult_22/ab[37][14] ,
         \mult_22/ab[37][15] , \mult_22/ab[37][16] , \mult_22/ab[37][17] ,
         \mult_22/ab[37][18] , \mult_22/ab[37][19] , \mult_22/ab[37][20] ,
         \mult_22/ab[37][21] , \mult_22/ab[37][22] , \mult_22/ab[37][23] ,
         \mult_22/ab[37][24] , \mult_22/ab[37][25] , \mult_22/ab[37][26] ,
         \mult_22/ab[37][27] , \mult_22/ab[37][28] , \mult_22/ab[37][29] ,
         \mult_22/ab[37][30] , \mult_22/ab[37][31] , \mult_22/ab[37][32] ,
         \mult_22/ab[37][33] , \mult_22/ab[37][34] , \mult_22/ab[37][35] ,
         \mult_22/ab[37][36] , \mult_22/ab[37][37] , \mult_22/ab[37][38] ,
         \mult_22/ab[37][39] , \mult_22/ab[37][40] , \mult_22/ab[37][41] ,
         \mult_22/ab[37][42] , \mult_22/ab[37][43] , \mult_22/ab[37][44] ,
         \mult_22/ab[37][45] , \mult_22/ab[37][46] , \mult_22/ab[37][47] ,
         \mult_22/ab[37][48] , \mult_22/ab[37][49] , \mult_22/ab[37][50] ,
         \mult_22/ab[37][51] , \mult_22/ab[37][52] , \mult_22/ab[37][53] ,
         \mult_22/ab[37][54] , \mult_22/ab[37][55] , \mult_22/ab[37][56] ,
         \mult_22/ab[37][57] , \mult_22/ab[37][58] , \mult_22/ab[37][59] ,
         \mult_22/ab[37][60] , \mult_22/ab[37][61] , \mult_22/ab[37][62] ,
         \mult_22/ab[37][63] , \mult_22/ab[38][0] , \mult_22/ab[38][1] ,
         \mult_22/ab[38][2] , \mult_22/ab[38][3] , \mult_22/ab[38][4] ,
         \mult_22/ab[38][5] , \mult_22/ab[38][6] , \mult_22/ab[38][7] ,
         \mult_22/ab[38][8] , \mult_22/ab[38][9] , \mult_22/ab[38][10] ,
         \mult_22/ab[38][11] , \mult_22/ab[38][12] , \mult_22/ab[38][13] ,
         \mult_22/ab[38][14] , \mult_22/ab[38][15] , \mult_22/ab[38][16] ,
         \mult_22/ab[38][17] , \mult_22/ab[38][18] , \mult_22/ab[38][19] ,
         \mult_22/ab[38][20] , \mult_22/ab[38][21] , \mult_22/ab[38][22] ,
         \mult_22/ab[38][23] , \mult_22/ab[38][24] , \mult_22/ab[38][25] ,
         \mult_22/ab[38][26] , \mult_22/ab[38][27] , \mult_22/ab[38][28] ,
         \mult_22/ab[38][29] , \mult_22/ab[38][30] , \mult_22/ab[38][31] ,
         \mult_22/ab[38][32] , \mult_22/ab[38][33] , \mult_22/ab[38][34] ,
         \mult_22/ab[38][35] , \mult_22/ab[38][36] , \mult_22/ab[38][37] ,
         \mult_22/ab[38][38] , \mult_22/ab[38][39] , \mult_22/ab[38][40] ,
         \mult_22/ab[38][41] , \mult_22/ab[38][42] , \mult_22/ab[38][43] ,
         \mult_22/ab[38][44] , \mult_22/ab[38][45] , \mult_22/ab[38][46] ,
         \mult_22/ab[38][47] , \mult_22/ab[38][48] , \mult_22/ab[38][49] ,
         \mult_22/ab[38][50] , \mult_22/ab[38][51] , \mult_22/ab[38][52] ,
         \mult_22/ab[38][53] , \mult_22/ab[38][54] , \mult_22/ab[38][55] ,
         \mult_22/ab[38][56] , \mult_22/ab[38][57] , \mult_22/ab[38][58] ,
         \mult_22/ab[38][59] , \mult_22/ab[38][60] , \mult_22/ab[38][61] ,
         \mult_22/ab[38][62] , \mult_22/ab[38][63] , \mult_22/ab[39][0] ,
         \mult_22/ab[39][1] , \mult_22/ab[39][2] , \mult_22/ab[39][3] ,
         \mult_22/ab[39][4] , \mult_22/ab[39][5] , \mult_22/ab[39][6] ,
         \mult_22/ab[39][7] , \mult_22/ab[39][8] , \mult_22/ab[39][9] ,
         \mult_22/ab[39][10] , \mult_22/ab[39][11] , \mult_22/ab[39][12] ,
         \mult_22/ab[39][13] , \mult_22/ab[39][14] , \mult_22/ab[39][15] ,
         \mult_22/ab[39][16] , \mult_22/ab[39][17] , \mult_22/ab[39][18] ,
         \mult_22/ab[39][19] , \mult_22/ab[39][20] , \mult_22/ab[39][21] ,
         \mult_22/ab[39][22] , \mult_22/ab[39][23] , \mult_22/ab[39][24] ,
         \mult_22/ab[39][25] , \mult_22/ab[39][26] , \mult_22/ab[39][27] ,
         \mult_22/ab[39][28] , \mult_22/ab[39][29] , \mult_22/ab[39][30] ,
         \mult_22/ab[39][31] , \mult_22/ab[39][32] , \mult_22/ab[39][33] ,
         \mult_22/ab[39][34] , \mult_22/ab[39][35] , \mult_22/ab[39][36] ,
         \mult_22/ab[39][37] , \mult_22/ab[39][38] , \mult_22/ab[39][39] ,
         \mult_22/ab[39][40] , \mult_22/ab[39][41] , \mult_22/ab[39][42] ,
         \mult_22/ab[39][43] , \mult_22/ab[39][44] , \mult_22/ab[39][45] ,
         \mult_22/ab[39][46] , \mult_22/ab[39][47] , \mult_22/ab[39][48] ,
         \mult_22/ab[39][49] , \mult_22/ab[39][50] , \mult_22/ab[39][51] ,
         \mult_22/ab[39][52] , \mult_22/ab[39][53] , \mult_22/ab[39][54] ,
         \mult_22/ab[39][55] , \mult_22/ab[39][56] , \mult_22/ab[39][57] ,
         \mult_22/ab[39][58] , \mult_22/ab[39][59] , \mult_22/ab[39][60] ,
         \mult_22/ab[39][61] , \mult_22/ab[39][62] , \mult_22/ab[39][63] ,
         \mult_22/ab[40][0] , \mult_22/ab[40][1] , \mult_22/ab[40][2] ,
         \mult_22/ab[40][3] , \mult_22/ab[40][4] , \mult_22/ab[40][5] ,
         \mult_22/ab[40][6] , \mult_22/ab[40][7] , \mult_22/ab[40][8] ,
         \mult_22/ab[40][9] , \mult_22/ab[40][10] , \mult_22/ab[40][11] ,
         \mult_22/ab[40][12] , \mult_22/ab[40][13] , \mult_22/ab[40][14] ,
         \mult_22/ab[40][15] , \mult_22/ab[40][16] , \mult_22/ab[40][17] ,
         \mult_22/ab[40][18] , \mult_22/ab[40][19] , \mult_22/ab[40][20] ,
         \mult_22/ab[40][21] , \mult_22/ab[40][22] , \mult_22/ab[40][23] ,
         \mult_22/ab[40][24] , \mult_22/ab[40][25] , \mult_22/ab[40][26] ,
         \mult_22/ab[40][27] , \mult_22/ab[40][28] , \mult_22/ab[40][29] ,
         \mult_22/ab[40][30] , \mult_22/ab[40][31] , \mult_22/ab[40][32] ,
         \mult_22/ab[40][33] , \mult_22/ab[40][34] , \mult_22/ab[40][35] ,
         \mult_22/ab[40][36] , \mult_22/ab[40][37] , \mult_22/ab[40][38] ,
         \mult_22/ab[40][39] , \mult_22/ab[40][40] , \mult_22/ab[40][41] ,
         \mult_22/ab[40][42] , \mult_22/ab[40][43] , \mult_22/ab[40][44] ,
         \mult_22/ab[40][45] , \mult_22/ab[40][46] , \mult_22/ab[40][47] ,
         \mult_22/ab[40][48] , \mult_22/ab[40][49] , \mult_22/ab[40][50] ,
         \mult_22/ab[40][51] , \mult_22/ab[40][52] , \mult_22/ab[40][53] ,
         \mult_22/ab[40][54] , \mult_22/ab[40][55] , \mult_22/ab[40][56] ,
         \mult_22/ab[40][57] , \mult_22/ab[40][58] , \mult_22/ab[40][59] ,
         \mult_22/ab[40][60] , \mult_22/ab[40][61] , \mult_22/ab[40][62] ,
         \mult_22/ab[40][63] , \mult_22/ab[41][0] , \mult_22/ab[41][1] ,
         \mult_22/ab[41][2] , \mult_22/ab[41][3] , \mult_22/ab[41][4] ,
         \mult_22/ab[41][5] , \mult_22/ab[41][6] , \mult_22/ab[41][7] ,
         \mult_22/ab[41][8] , \mult_22/ab[41][9] , \mult_22/ab[41][10] ,
         \mult_22/ab[41][11] , \mult_22/ab[41][12] , \mult_22/ab[41][13] ,
         \mult_22/ab[41][14] , \mult_22/ab[41][15] , \mult_22/ab[41][16] ,
         \mult_22/ab[41][17] , \mult_22/ab[41][18] , \mult_22/ab[41][19] ,
         \mult_22/ab[41][20] , \mult_22/ab[41][21] , \mult_22/ab[41][22] ,
         \mult_22/ab[41][23] , \mult_22/ab[41][24] , \mult_22/ab[41][25] ,
         \mult_22/ab[41][26] , \mult_22/ab[41][27] , \mult_22/ab[41][28] ,
         \mult_22/ab[41][29] , \mult_22/ab[41][30] , \mult_22/ab[41][31] ,
         \mult_22/ab[41][32] , \mult_22/ab[41][33] , \mult_22/ab[41][34] ,
         \mult_22/ab[41][35] , \mult_22/ab[41][36] , \mult_22/ab[41][37] ,
         \mult_22/ab[41][38] , \mult_22/ab[41][39] , \mult_22/ab[41][40] ,
         \mult_22/ab[41][41] , \mult_22/ab[41][42] , \mult_22/ab[41][43] ,
         \mult_22/ab[41][44] , \mult_22/ab[41][45] , \mult_22/ab[41][46] ,
         \mult_22/ab[41][47] , \mult_22/ab[41][48] , \mult_22/ab[41][49] ,
         \mult_22/ab[41][50] , \mult_22/ab[41][51] , \mult_22/ab[41][52] ,
         \mult_22/ab[41][53] , \mult_22/ab[41][54] , \mult_22/ab[41][55] ,
         \mult_22/ab[41][56] , \mult_22/ab[41][57] , \mult_22/ab[41][58] ,
         \mult_22/ab[41][59] , \mult_22/ab[41][60] , \mult_22/ab[41][61] ,
         \mult_22/ab[41][62] , \mult_22/ab[41][63] , \mult_22/ab[42][0] ,
         \mult_22/ab[42][1] , \mult_22/ab[42][2] , \mult_22/ab[42][3] ,
         \mult_22/ab[42][4] , \mult_22/ab[42][5] , \mult_22/ab[42][6] ,
         \mult_22/ab[42][7] , \mult_22/ab[42][8] , \mult_22/ab[42][9] ,
         \mult_22/ab[42][10] , \mult_22/ab[42][11] , \mult_22/ab[42][12] ,
         \mult_22/ab[42][13] , \mult_22/ab[42][14] , \mult_22/ab[42][15] ,
         \mult_22/ab[42][16] , \mult_22/ab[42][17] , \mult_22/ab[42][18] ,
         \mult_22/ab[42][19] , \mult_22/ab[42][20] , \mult_22/ab[42][21] ,
         \mult_22/ab[42][22] , \mult_22/ab[42][23] , \mult_22/ab[42][24] ,
         \mult_22/ab[42][25] , \mult_22/ab[42][26] , \mult_22/ab[42][27] ,
         \mult_22/ab[42][28] , \mult_22/ab[42][29] , \mult_22/ab[42][30] ,
         \mult_22/ab[42][31] , \mult_22/ab[42][32] , \mult_22/ab[42][33] ,
         \mult_22/ab[42][34] , \mult_22/ab[42][35] , \mult_22/ab[42][36] ,
         \mult_22/ab[42][37] , \mult_22/ab[42][38] , \mult_22/ab[42][39] ,
         \mult_22/ab[42][40] , \mult_22/ab[42][41] , \mult_22/ab[42][42] ,
         \mult_22/ab[42][43] , \mult_22/ab[42][44] , \mult_22/ab[42][45] ,
         \mult_22/ab[42][46] , \mult_22/ab[42][47] , \mult_22/ab[42][48] ,
         \mult_22/ab[42][49] , \mult_22/ab[42][50] , \mult_22/ab[42][51] ,
         \mult_22/ab[42][52] , \mult_22/ab[42][53] , \mult_22/ab[42][54] ,
         \mult_22/ab[42][55] , \mult_22/ab[42][56] , \mult_22/ab[42][57] ,
         \mult_22/ab[42][58] , \mult_22/ab[42][59] , \mult_22/ab[42][60] ,
         \mult_22/ab[42][61] , \mult_22/ab[42][62] , \mult_22/ab[42][63] ,
         \mult_22/ab[43][0] , \mult_22/ab[43][1] , \mult_22/ab[43][2] ,
         \mult_22/ab[43][3] , \mult_22/ab[43][4] , \mult_22/ab[43][5] ,
         \mult_22/ab[43][6] , \mult_22/ab[43][7] , \mult_22/ab[43][8] ,
         \mult_22/ab[43][9] , \mult_22/ab[43][10] , \mult_22/ab[43][11] ,
         \mult_22/ab[43][12] , \mult_22/ab[43][13] , \mult_22/ab[43][14] ,
         \mult_22/ab[43][15] , \mult_22/ab[43][16] , \mult_22/ab[43][17] ,
         \mult_22/ab[43][18] , \mult_22/ab[43][19] , \mult_22/ab[43][20] ,
         \mult_22/ab[43][21] , \mult_22/ab[43][22] , \mult_22/ab[43][23] ,
         \mult_22/ab[43][24] , \mult_22/ab[43][25] , \mult_22/ab[43][26] ,
         \mult_22/ab[43][27] , \mult_22/ab[43][28] , \mult_22/ab[43][29] ,
         \mult_22/ab[43][30] , \mult_22/ab[43][31] , \mult_22/ab[43][32] ,
         \mult_22/ab[43][33] , \mult_22/ab[43][34] , \mult_22/ab[43][35] ,
         \mult_22/ab[43][36] , \mult_22/ab[43][37] , \mult_22/ab[43][38] ,
         \mult_22/ab[43][39] , \mult_22/ab[43][40] , \mult_22/ab[43][41] ,
         \mult_22/ab[43][42] , \mult_22/ab[43][43] , \mult_22/ab[43][44] ,
         \mult_22/ab[43][45] , \mult_22/ab[43][46] , \mult_22/ab[43][47] ,
         \mult_22/ab[43][48] , \mult_22/ab[43][49] , \mult_22/ab[43][50] ,
         \mult_22/ab[43][51] , \mult_22/ab[43][52] , \mult_22/ab[43][53] ,
         \mult_22/ab[43][54] , \mult_22/ab[43][55] , \mult_22/ab[43][56] ,
         \mult_22/ab[43][57] , \mult_22/ab[43][58] , \mult_22/ab[43][59] ,
         \mult_22/ab[43][60] , \mult_22/ab[43][61] , \mult_22/ab[43][62] ,
         \mult_22/ab[43][63] , \mult_22/ab[44][0] , \mult_22/ab[44][1] ,
         \mult_22/ab[44][2] , \mult_22/ab[44][3] , \mult_22/ab[44][4] ,
         \mult_22/ab[44][5] , \mult_22/ab[44][6] , \mult_22/ab[44][7] ,
         \mult_22/ab[44][8] , \mult_22/ab[44][9] , \mult_22/ab[44][10] ,
         \mult_22/ab[44][11] , \mult_22/ab[44][12] , \mult_22/ab[44][13] ,
         \mult_22/ab[44][14] , \mult_22/ab[44][15] , \mult_22/ab[44][16] ,
         \mult_22/ab[44][17] , \mult_22/ab[44][18] , \mult_22/ab[44][19] ,
         \mult_22/ab[44][20] , \mult_22/ab[44][21] , \mult_22/ab[44][22] ,
         \mult_22/ab[44][23] , \mult_22/ab[44][24] , \mult_22/ab[44][25] ,
         \mult_22/ab[44][26] , \mult_22/ab[44][27] , \mult_22/ab[44][28] ,
         \mult_22/ab[44][29] , \mult_22/ab[44][30] , \mult_22/ab[44][31] ,
         \mult_22/ab[44][32] , \mult_22/ab[44][33] , \mult_22/ab[44][34] ,
         \mult_22/ab[44][35] , \mult_22/ab[44][36] , \mult_22/ab[44][37] ,
         \mult_22/ab[44][38] , \mult_22/ab[44][39] , \mult_22/ab[44][40] ,
         \mult_22/ab[44][41] , \mult_22/ab[44][42] , \mult_22/ab[44][43] ,
         \mult_22/ab[44][44] , \mult_22/ab[44][45] , \mult_22/ab[44][46] ,
         \mult_22/ab[44][47] , \mult_22/ab[44][48] , \mult_22/ab[44][49] ,
         \mult_22/ab[44][50] , \mult_22/ab[44][51] , \mult_22/ab[44][52] ,
         \mult_22/ab[44][53] , \mult_22/ab[44][54] , \mult_22/ab[44][55] ,
         \mult_22/ab[44][56] , \mult_22/ab[44][57] , \mult_22/ab[44][58] ,
         \mult_22/ab[44][59] , \mult_22/ab[44][60] , \mult_22/ab[44][61] ,
         \mult_22/ab[44][62] , \mult_22/ab[44][63] , \mult_22/ab[45][0] ,
         \mult_22/ab[45][1] , \mult_22/ab[45][2] , \mult_22/ab[45][3] ,
         \mult_22/ab[45][4] , \mult_22/ab[45][5] , \mult_22/ab[45][6] ,
         \mult_22/ab[45][7] , \mult_22/ab[45][8] , \mult_22/ab[45][9] ,
         \mult_22/ab[45][10] , \mult_22/ab[45][11] , \mult_22/ab[45][12] ,
         \mult_22/ab[45][13] , \mult_22/ab[45][14] , \mult_22/ab[45][15] ,
         \mult_22/ab[45][16] , \mult_22/ab[45][17] , \mult_22/ab[45][18] ,
         \mult_22/ab[45][19] , \mult_22/ab[45][20] , \mult_22/ab[45][21] ,
         \mult_22/ab[45][22] , \mult_22/ab[45][23] , \mult_22/ab[45][24] ,
         \mult_22/ab[45][25] , \mult_22/ab[45][26] , \mult_22/ab[45][27] ,
         \mult_22/ab[45][28] , \mult_22/ab[45][29] , \mult_22/ab[45][30] ,
         \mult_22/ab[45][31] , \mult_22/ab[45][32] , \mult_22/ab[45][33] ,
         \mult_22/ab[45][34] , \mult_22/ab[45][35] , \mult_22/ab[45][36] ,
         \mult_22/ab[45][37] , \mult_22/ab[45][38] , \mult_22/ab[45][39] ,
         \mult_22/ab[45][40] , \mult_22/ab[45][41] , \mult_22/ab[45][42] ,
         \mult_22/ab[45][43] , \mult_22/ab[45][44] , \mult_22/ab[45][45] ,
         \mult_22/ab[45][46] , \mult_22/ab[45][47] , \mult_22/ab[45][48] ,
         \mult_22/ab[45][49] , \mult_22/ab[45][50] , \mult_22/ab[45][51] ,
         \mult_22/ab[45][52] , \mult_22/ab[45][53] , \mult_22/ab[45][54] ,
         \mult_22/ab[45][55] , \mult_22/ab[45][56] , \mult_22/ab[45][57] ,
         \mult_22/ab[45][58] , \mult_22/ab[45][59] , \mult_22/ab[45][60] ,
         \mult_22/ab[45][61] , \mult_22/ab[45][62] , \mult_22/ab[45][63] ,
         \mult_22/ab[46][0] , \mult_22/ab[46][1] , \mult_22/ab[46][2] ,
         \mult_22/ab[46][3] , \mult_22/ab[46][4] , \mult_22/ab[46][5] ,
         \mult_22/ab[46][6] , \mult_22/ab[46][7] , \mult_22/ab[46][8] ,
         \mult_22/ab[46][9] , \mult_22/ab[46][10] , \mult_22/ab[46][11] ,
         \mult_22/ab[46][12] , \mult_22/ab[46][13] , \mult_22/ab[46][14] ,
         \mult_22/ab[46][15] , \mult_22/ab[46][16] , \mult_22/ab[46][17] ,
         \mult_22/ab[46][18] , \mult_22/ab[46][19] , \mult_22/ab[46][20] ,
         \mult_22/ab[46][21] , \mult_22/ab[46][22] , \mult_22/ab[46][23] ,
         \mult_22/ab[46][24] , \mult_22/ab[46][25] , \mult_22/ab[46][26] ,
         \mult_22/ab[46][27] , \mult_22/ab[46][28] , \mult_22/ab[46][29] ,
         \mult_22/ab[46][30] , \mult_22/ab[46][31] , \mult_22/ab[46][32] ,
         \mult_22/ab[46][33] , \mult_22/ab[46][34] , \mult_22/ab[46][35] ,
         \mult_22/ab[46][36] , \mult_22/ab[46][37] , \mult_22/ab[46][38] ,
         \mult_22/ab[46][39] , \mult_22/ab[46][40] , \mult_22/ab[46][41] ,
         \mult_22/ab[46][42] , \mult_22/ab[46][43] , \mult_22/ab[46][44] ,
         \mult_22/ab[46][45] , \mult_22/ab[46][46] , \mult_22/ab[46][47] ,
         \mult_22/ab[46][48] , \mult_22/ab[46][49] , \mult_22/ab[46][50] ,
         \mult_22/ab[46][51] , \mult_22/ab[46][52] , \mult_22/ab[46][53] ,
         \mult_22/ab[46][54] , \mult_22/ab[46][55] , \mult_22/ab[46][56] ,
         \mult_22/ab[46][57] , \mult_22/ab[46][58] , \mult_22/ab[46][59] ,
         \mult_22/ab[46][60] , \mult_22/ab[46][61] , \mult_22/ab[46][62] ,
         \mult_22/ab[46][63] , \mult_22/ab[47][0] , \mult_22/ab[47][1] ,
         \mult_22/ab[47][2] , \mult_22/ab[47][3] , \mult_22/ab[47][4] ,
         \mult_22/ab[47][5] , \mult_22/ab[47][6] , \mult_22/ab[47][7] ,
         \mult_22/ab[47][8] , \mult_22/ab[47][9] , \mult_22/ab[47][10] ,
         \mult_22/ab[47][11] , \mult_22/ab[47][12] , \mult_22/ab[47][13] ,
         \mult_22/ab[47][14] , \mult_22/ab[47][15] , \mult_22/ab[47][16] ,
         \mult_22/ab[47][17] , \mult_22/ab[47][18] , \mult_22/ab[47][19] ,
         \mult_22/ab[47][20] , \mult_22/ab[47][21] , \mult_22/ab[47][22] ,
         \mult_22/ab[47][23] , \mult_22/ab[47][24] , \mult_22/ab[47][25] ,
         \mult_22/ab[47][26] , \mult_22/ab[47][27] , \mult_22/ab[47][28] ,
         \mult_22/ab[47][29] , \mult_22/ab[47][30] , \mult_22/ab[47][31] ,
         \mult_22/ab[47][32] , \mult_22/ab[47][33] , \mult_22/ab[47][34] ,
         \mult_22/ab[47][35] , \mult_22/ab[47][36] , \mult_22/ab[47][37] ,
         \mult_22/ab[47][38] , \mult_22/ab[47][39] , \mult_22/ab[47][40] ,
         \mult_22/ab[47][41] , \mult_22/ab[47][42] , \mult_22/ab[47][43] ,
         \mult_22/ab[47][44] , \mult_22/ab[47][45] , \mult_22/ab[47][46] ,
         \mult_22/ab[47][47] , \mult_22/ab[47][48] , \mult_22/ab[47][49] ,
         \mult_22/ab[47][50] , \mult_22/ab[47][51] , \mult_22/ab[47][52] ,
         \mult_22/ab[47][53] , \mult_22/ab[47][54] , \mult_22/ab[47][55] ,
         \mult_22/ab[47][56] , \mult_22/ab[47][57] , \mult_22/ab[47][58] ,
         \mult_22/ab[47][59] , \mult_22/ab[47][60] , \mult_22/ab[47][61] ,
         \mult_22/ab[47][62] , \mult_22/ab[47][63] , \mult_22/ab[48][0] ,
         \mult_22/ab[48][1] , \mult_22/ab[48][2] , \mult_22/ab[48][3] ,
         \mult_22/ab[48][4] , \mult_22/ab[48][5] , \mult_22/ab[48][6] ,
         \mult_22/ab[48][7] , \mult_22/ab[48][8] , \mult_22/ab[48][9] ,
         \mult_22/ab[48][10] , \mult_22/ab[48][11] , \mult_22/ab[48][12] ,
         \mult_22/ab[48][13] , \mult_22/ab[48][14] , \mult_22/ab[48][15] ,
         \mult_22/ab[48][16] , \mult_22/ab[48][17] , \mult_22/ab[48][18] ,
         \mult_22/ab[48][19] , \mult_22/ab[48][20] , \mult_22/ab[48][21] ,
         \mult_22/ab[48][22] , \mult_22/ab[48][23] , \mult_22/ab[48][24] ,
         \mult_22/ab[48][25] , \mult_22/ab[48][26] , \mult_22/ab[48][27] ,
         \mult_22/ab[48][28] , \mult_22/ab[48][29] , \mult_22/ab[48][30] ,
         \mult_22/ab[48][31] , \mult_22/ab[48][32] , \mult_22/ab[48][33] ,
         \mult_22/ab[48][34] , \mult_22/ab[48][35] , \mult_22/ab[48][36] ,
         \mult_22/ab[48][37] , \mult_22/ab[48][38] , \mult_22/ab[48][39] ,
         \mult_22/ab[48][40] , \mult_22/ab[48][41] , \mult_22/ab[48][42] ,
         \mult_22/ab[48][43] , \mult_22/ab[48][44] , \mult_22/ab[48][45] ,
         \mult_22/ab[48][46] , \mult_22/ab[48][47] , \mult_22/ab[48][48] ,
         \mult_22/ab[48][49] , \mult_22/ab[48][50] , \mult_22/ab[48][51] ,
         \mult_22/ab[48][52] , \mult_22/ab[48][53] , \mult_22/ab[48][54] ,
         \mult_22/ab[48][55] , \mult_22/ab[48][56] , \mult_22/ab[48][57] ,
         \mult_22/ab[48][58] , \mult_22/ab[48][59] , \mult_22/ab[48][60] ,
         \mult_22/ab[48][61] , \mult_22/ab[48][62] , \mult_22/ab[48][63] ,
         \mult_22/ab[49][0] , \mult_22/ab[49][1] , \mult_22/ab[49][2] ,
         \mult_22/ab[49][3] , \mult_22/ab[49][4] , \mult_22/ab[49][5] ,
         \mult_22/ab[49][6] , \mult_22/ab[49][7] , \mult_22/ab[49][8] ,
         \mult_22/ab[49][9] , \mult_22/ab[49][10] , \mult_22/ab[49][11] ,
         \mult_22/ab[49][12] , \mult_22/ab[49][13] , \mult_22/ab[49][14] ,
         \mult_22/ab[49][15] , \mult_22/ab[49][16] , \mult_22/ab[49][17] ,
         \mult_22/ab[49][18] , \mult_22/ab[49][19] , \mult_22/ab[49][20] ,
         \mult_22/ab[49][21] , \mult_22/ab[49][22] , \mult_22/ab[49][23] ,
         \mult_22/ab[49][24] , \mult_22/ab[49][25] , \mult_22/ab[49][26] ,
         \mult_22/ab[49][27] , \mult_22/ab[49][28] , \mult_22/ab[49][29] ,
         \mult_22/ab[49][30] , \mult_22/ab[49][31] , \mult_22/ab[49][32] ,
         \mult_22/ab[49][33] , \mult_22/ab[49][34] , \mult_22/ab[49][35] ,
         \mult_22/ab[49][36] , \mult_22/ab[49][37] , \mult_22/ab[49][38] ,
         \mult_22/ab[49][39] , \mult_22/ab[49][40] , \mult_22/ab[49][41] ,
         \mult_22/ab[49][42] , \mult_22/ab[49][43] , \mult_22/ab[49][44] ,
         \mult_22/ab[49][45] , \mult_22/ab[49][46] , \mult_22/ab[49][47] ,
         \mult_22/ab[49][48] , \mult_22/ab[49][49] , \mult_22/ab[49][50] ,
         \mult_22/ab[49][51] , \mult_22/ab[49][52] , \mult_22/ab[49][53] ,
         \mult_22/ab[49][54] , \mult_22/ab[49][55] , \mult_22/ab[49][56] ,
         \mult_22/ab[49][57] , \mult_22/ab[49][58] , \mult_22/ab[49][59] ,
         \mult_22/ab[49][60] , \mult_22/ab[49][61] , \mult_22/ab[49][62] ,
         \mult_22/ab[49][63] , \mult_22/ab[50][0] , \mult_22/ab[50][1] ,
         \mult_22/ab[50][2] , \mult_22/ab[50][3] , \mult_22/ab[50][4] ,
         \mult_22/ab[50][5] , \mult_22/ab[50][6] , \mult_22/ab[50][7] ,
         \mult_22/ab[50][8] , \mult_22/ab[50][9] , \mult_22/ab[50][10] ,
         \mult_22/ab[50][11] , \mult_22/ab[50][12] , \mult_22/ab[50][13] ,
         \mult_22/ab[50][14] , \mult_22/ab[50][15] , \mult_22/ab[50][16] ,
         \mult_22/ab[50][17] , \mult_22/ab[50][18] , \mult_22/ab[50][19] ,
         \mult_22/ab[50][20] , \mult_22/ab[50][21] , \mult_22/ab[50][22] ,
         \mult_22/ab[50][23] , \mult_22/ab[50][24] , \mult_22/ab[50][25] ,
         \mult_22/ab[50][26] , \mult_22/ab[50][27] , \mult_22/ab[50][28] ,
         \mult_22/ab[50][29] , \mult_22/ab[50][30] , \mult_22/ab[50][31] ,
         \mult_22/ab[50][32] , \mult_22/ab[50][33] , \mult_22/ab[50][34] ,
         \mult_22/ab[50][35] , \mult_22/ab[50][36] , \mult_22/ab[50][37] ,
         \mult_22/ab[50][38] , \mult_22/ab[50][39] , \mult_22/ab[50][40] ,
         \mult_22/ab[50][41] , \mult_22/ab[50][42] , \mult_22/ab[50][43] ,
         \mult_22/ab[50][44] , \mult_22/ab[50][45] , \mult_22/ab[50][46] ,
         \mult_22/ab[50][47] , \mult_22/ab[50][48] , \mult_22/ab[50][49] ,
         \mult_22/ab[50][50] , \mult_22/ab[50][51] , \mult_22/ab[50][52] ,
         \mult_22/ab[50][53] , \mult_22/ab[50][54] , \mult_22/ab[50][55] ,
         \mult_22/ab[50][56] , \mult_22/ab[50][57] , \mult_22/ab[50][58] ,
         \mult_22/ab[50][59] , \mult_22/ab[50][60] , \mult_22/ab[50][61] ,
         \mult_22/ab[50][62] , \mult_22/ab[50][63] , \mult_22/ab[51][0] ,
         \mult_22/ab[51][1] , \mult_22/ab[51][2] , \mult_22/ab[51][3] ,
         \mult_22/ab[51][4] , \mult_22/ab[51][5] , \mult_22/ab[51][6] ,
         \mult_22/ab[51][7] , \mult_22/ab[51][8] , \mult_22/ab[51][9] ,
         \mult_22/ab[51][10] , \mult_22/ab[51][11] , \mult_22/ab[51][12] ,
         \mult_22/ab[51][13] , \mult_22/ab[51][14] , \mult_22/ab[51][15] ,
         \mult_22/ab[51][16] , \mult_22/ab[51][17] , \mult_22/ab[51][18] ,
         \mult_22/ab[51][19] , \mult_22/ab[51][20] , \mult_22/ab[51][21] ,
         \mult_22/ab[51][22] , \mult_22/ab[51][23] , \mult_22/ab[51][24] ,
         \mult_22/ab[51][25] , \mult_22/ab[51][26] , \mult_22/ab[51][27] ,
         \mult_22/ab[51][28] , \mult_22/ab[51][29] , \mult_22/ab[51][30] ,
         \mult_22/ab[51][31] , \mult_22/ab[51][32] , \mult_22/ab[51][33] ,
         \mult_22/ab[51][34] , \mult_22/ab[51][35] , \mult_22/ab[51][36] ,
         \mult_22/ab[51][37] , \mult_22/ab[51][38] , \mult_22/ab[51][39] ,
         \mult_22/ab[51][40] , \mult_22/ab[51][41] , \mult_22/ab[51][42] ,
         \mult_22/ab[51][43] , \mult_22/ab[51][44] , \mult_22/ab[51][45] ,
         \mult_22/ab[51][46] , \mult_22/ab[51][47] , \mult_22/ab[51][48] ,
         \mult_22/ab[51][49] , \mult_22/ab[51][50] , \mult_22/ab[51][51] ,
         \mult_22/ab[51][52] , \mult_22/ab[51][53] , \mult_22/ab[51][54] ,
         \mult_22/ab[51][55] , \mult_22/ab[51][56] , \mult_22/ab[51][57] ,
         \mult_22/ab[51][58] , \mult_22/ab[51][59] , \mult_22/ab[51][60] ,
         \mult_22/ab[51][61] , \mult_22/ab[51][62] , \mult_22/ab[51][63] ,
         \mult_22/ab[52][0] , \mult_22/ab[52][1] , \mult_22/ab[52][2] ,
         \mult_22/ab[52][3] , \mult_22/ab[52][4] , \mult_22/ab[52][5] ,
         \mult_22/ab[52][6] , \mult_22/ab[52][7] , \mult_22/ab[52][8] ,
         \mult_22/ab[52][9] , \mult_22/ab[52][10] , \mult_22/ab[52][11] ,
         \mult_22/ab[52][12] , \mult_22/ab[52][13] , \mult_22/ab[52][14] ,
         \mult_22/ab[52][15] , \mult_22/ab[52][16] , \mult_22/ab[52][17] ,
         \mult_22/ab[52][18] , \mult_22/ab[52][19] , \mult_22/ab[52][20] ,
         \mult_22/ab[52][21] , \mult_22/ab[52][22] , \mult_22/ab[52][23] ,
         \mult_22/ab[52][24] , \mult_22/ab[52][25] , \mult_22/ab[52][26] ,
         \mult_22/ab[52][27] , \mult_22/ab[52][28] , \mult_22/ab[52][29] ,
         \mult_22/ab[52][30] , \mult_22/ab[52][31] , \mult_22/ab[52][32] ,
         \mult_22/ab[52][33] , \mult_22/ab[52][34] , \mult_22/ab[52][35] ,
         \mult_22/ab[52][36] , \mult_22/ab[52][37] , \mult_22/ab[52][38] ,
         \mult_22/ab[52][39] , \mult_22/ab[52][40] , \mult_22/ab[52][41] ,
         \mult_22/ab[52][42] , \mult_22/ab[52][43] , \mult_22/ab[52][44] ,
         \mult_22/ab[52][45] , \mult_22/ab[52][46] , \mult_22/ab[52][47] ,
         \mult_22/ab[52][48] , \mult_22/ab[52][49] , \mult_22/ab[52][50] ,
         \mult_22/ab[52][51] , \mult_22/ab[52][52] , \mult_22/ab[52][53] ,
         \mult_22/ab[52][54] , \mult_22/ab[52][55] , \mult_22/ab[52][56] ,
         \mult_22/ab[52][57] , \mult_22/ab[52][58] , \mult_22/ab[52][59] ,
         \mult_22/ab[52][60] , \mult_22/ab[52][61] , \mult_22/ab[52][62] ,
         \mult_22/ab[52][63] , \mult_22/ab[53][0] , \mult_22/ab[53][1] ,
         \mult_22/ab[53][2] , \mult_22/ab[53][3] , \mult_22/ab[53][4] ,
         \mult_22/ab[53][5] , \mult_22/ab[53][6] , \mult_22/ab[53][7] ,
         \mult_22/ab[53][8] , \mult_22/ab[53][9] , \mult_22/ab[53][10] ,
         \mult_22/ab[53][11] , \mult_22/ab[53][12] , \mult_22/ab[53][13] ,
         \mult_22/ab[53][14] , \mult_22/ab[53][15] , \mult_22/ab[53][16] ,
         \mult_22/ab[53][17] , \mult_22/ab[53][18] , \mult_22/ab[53][19] ,
         \mult_22/ab[53][20] , \mult_22/ab[53][21] , \mult_22/ab[53][22] ,
         \mult_22/ab[53][23] , \mult_22/ab[53][24] , \mult_22/ab[53][25] ,
         \mult_22/ab[53][26] , \mult_22/ab[53][27] , \mult_22/ab[53][28] ,
         \mult_22/ab[53][29] , \mult_22/ab[53][30] , \mult_22/ab[53][31] ,
         \mult_22/ab[53][32] , \mult_22/ab[53][33] , \mult_22/ab[53][34] ,
         \mult_22/ab[53][35] , \mult_22/ab[53][36] , \mult_22/ab[53][37] ,
         \mult_22/ab[53][38] , \mult_22/ab[53][39] , \mult_22/ab[53][40] ,
         \mult_22/ab[53][41] , \mult_22/ab[53][42] , \mult_22/ab[53][43] ,
         \mult_22/ab[53][44] , \mult_22/ab[53][45] , \mult_22/ab[53][46] ,
         \mult_22/ab[53][47] , \mult_22/ab[53][48] , \mult_22/ab[53][49] ,
         \mult_22/ab[53][50] , \mult_22/ab[53][51] , \mult_22/ab[53][52] ,
         \mult_22/ab[53][53] , \mult_22/ab[53][54] , \mult_22/ab[53][55] ,
         \mult_22/ab[53][56] , \mult_22/ab[53][57] , \mult_22/ab[53][58] ,
         \mult_22/ab[53][59] , \mult_22/ab[53][60] , \mult_22/ab[53][61] ,
         \mult_22/ab[53][62] , \mult_22/ab[53][63] , \mult_22/ab[54][0] ,
         \mult_22/ab[54][1] , \mult_22/ab[54][2] , \mult_22/ab[54][3] ,
         \mult_22/ab[54][4] , \mult_22/ab[54][5] , \mult_22/ab[54][6] ,
         \mult_22/ab[54][7] , \mult_22/ab[54][8] , \mult_22/ab[54][9] ,
         \mult_22/ab[54][10] , \mult_22/ab[54][11] , \mult_22/ab[54][12] ,
         \mult_22/ab[54][13] , \mult_22/ab[54][14] , \mult_22/ab[54][15] ,
         \mult_22/ab[54][16] , \mult_22/ab[54][17] , \mult_22/ab[54][18] ,
         \mult_22/ab[54][19] , \mult_22/ab[54][20] , \mult_22/ab[54][21] ,
         \mult_22/ab[54][22] , \mult_22/ab[54][23] , \mult_22/ab[54][24] ,
         \mult_22/ab[54][25] , \mult_22/ab[54][26] , \mult_22/ab[54][27] ,
         \mult_22/ab[54][28] , \mult_22/ab[54][29] , \mult_22/ab[54][30] ,
         \mult_22/ab[54][31] , \mult_22/ab[54][32] , \mult_22/ab[54][33] ,
         \mult_22/ab[54][34] , \mult_22/ab[54][35] , \mult_22/ab[54][36] ,
         \mult_22/ab[54][37] , \mult_22/ab[54][38] , \mult_22/ab[54][39] ,
         \mult_22/ab[54][40] , \mult_22/ab[54][41] , \mult_22/ab[54][42] ,
         \mult_22/ab[54][43] , \mult_22/ab[54][44] , \mult_22/ab[54][45] ,
         \mult_22/ab[54][46] , \mult_22/ab[54][47] , \mult_22/ab[54][48] ,
         \mult_22/ab[54][49] , \mult_22/ab[54][50] , \mult_22/ab[54][51] ,
         \mult_22/ab[54][52] , \mult_22/ab[54][53] , \mult_22/ab[54][54] ,
         \mult_22/ab[54][55] , \mult_22/ab[54][56] , \mult_22/ab[54][57] ,
         \mult_22/ab[54][58] , \mult_22/ab[54][59] , \mult_22/ab[54][60] ,
         \mult_22/ab[54][61] , \mult_22/ab[54][62] , \mult_22/ab[54][63] ,
         \mult_22/ab[55][0] , \mult_22/ab[55][1] , \mult_22/ab[55][2] ,
         \mult_22/ab[55][3] , \mult_22/ab[55][4] , \mult_22/ab[55][5] ,
         \mult_22/ab[55][6] , \mult_22/ab[55][7] , \mult_22/ab[55][8] ,
         \mult_22/ab[55][9] , \mult_22/ab[55][10] , \mult_22/ab[55][11] ,
         \mult_22/ab[55][12] , \mult_22/ab[55][13] , \mult_22/ab[55][14] ,
         \mult_22/ab[55][15] , \mult_22/ab[55][16] , \mult_22/ab[55][17] ,
         \mult_22/ab[55][18] , \mult_22/ab[55][19] , \mult_22/ab[55][20] ,
         \mult_22/ab[55][21] , \mult_22/ab[55][22] , \mult_22/ab[55][23] ,
         \mult_22/ab[55][24] , \mult_22/ab[55][25] , \mult_22/ab[55][26] ,
         \mult_22/ab[55][27] , \mult_22/ab[55][28] , \mult_22/ab[55][29] ,
         \mult_22/ab[55][30] , \mult_22/ab[55][31] , \mult_22/ab[55][32] ,
         \mult_22/ab[55][33] , \mult_22/ab[55][34] , \mult_22/ab[55][35] ,
         \mult_22/ab[55][36] , \mult_22/ab[55][37] , \mult_22/ab[55][38] ,
         \mult_22/ab[55][39] , \mult_22/ab[55][40] , \mult_22/ab[55][41] ,
         \mult_22/ab[55][42] , \mult_22/ab[55][43] , \mult_22/ab[55][44] ,
         \mult_22/ab[55][45] , \mult_22/ab[55][46] , \mult_22/ab[55][47] ,
         \mult_22/ab[55][48] , \mult_22/ab[55][49] , \mult_22/ab[55][50] ,
         \mult_22/ab[55][51] , \mult_22/ab[55][52] , \mult_22/ab[55][53] ,
         \mult_22/ab[55][54] , \mult_22/ab[55][55] , \mult_22/ab[55][56] ,
         \mult_22/ab[55][57] , \mult_22/ab[55][58] , \mult_22/ab[55][59] ,
         \mult_22/ab[55][60] , \mult_22/ab[55][61] , \mult_22/ab[55][62] ,
         \mult_22/ab[55][63] , \mult_22/ab[56][0] , \mult_22/ab[56][1] ,
         \mult_22/ab[56][2] , \mult_22/ab[56][3] , \mult_22/ab[56][4] ,
         \mult_22/ab[56][5] , \mult_22/ab[56][6] , \mult_22/ab[56][7] ,
         \mult_22/ab[56][8] , \mult_22/ab[56][9] , \mult_22/ab[56][10] ,
         \mult_22/ab[56][11] , \mult_22/ab[56][12] , \mult_22/ab[56][13] ,
         \mult_22/ab[56][14] , \mult_22/ab[56][15] , \mult_22/ab[56][16] ,
         \mult_22/ab[56][17] , \mult_22/ab[56][18] , \mult_22/ab[56][19] ,
         \mult_22/ab[56][20] , \mult_22/ab[56][21] , \mult_22/ab[56][22] ,
         \mult_22/ab[56][23] , \mult_22/ab[56][24] , \mult_22/ab[56][25] ,
         \mult_22/ab[56][26] , \mult_22/ab[56][27] , \mult_22/ab[56][28] ,
         \mult_22/ab[56][29] , \mult_22/ab[56][30] , \mult_22/ab[56][31] ,
         \mult_22/ab[56][32] , \mult_22/ab[56][33] , \mult_22/ab[56][34] ,
         \mult_22/ab[56][35] , \mult_22/ab[56][36] , \mult_22/ab[56][37] ,
         \mult_22/ab[56][38] , \mult_22/ab[56][39] , \mult_22/ab[56][40] ,
         \mult_22/ab[56][41] , \mult_22/ab[56][42] , \mult_22/ab[56][43] ,
         \mult_22/ab[56][44] , \mult_22/ab[56][45] , \mult_22/ab[56][46] ,
         \mult_22/ab[56][47] , \mult_22/ab[56][48] , \mult_22/ab[56][49] ,
         \mult_22/ab[56][50] , \mult_22/ab[56][51] , \mult_22/ab[56][52] ,
         \mult_22/ab[56][53] , \mult_22/ab[56][54] , \mult_22/ab[56][55] ,
         \mult_22/ab[56][56] , \mult_22/ab[56][57] , \mult_22/ab[56][58] ,
         \mult_22/ab[56][59] , \mult_22/ab[56][60] , \mult_22/ab[56][61] ,
         \mult_22/ab[56][62] , \mult_22/ab[56][63] , \mult_22/ab[57][0] ,
         \mult_22/ab[57][1] , \mult_22/ab[57][2] , \mult_22/ab[57][3] ,
         \mult_22/ab[57][4] , \mult_22/ab[57][5] , \mult_22/ab[57][6] ,
         \mult_22/ab[57][7] , \mult_22/ab[57][8] , \mult_22/ab[57][9] ,
         \mult_22/ab[57][10] , \mult_22/ab[57][11] , \mult_22/ab[57][12] ,
         \mult_22/ab[57][13] , \mult_22/ab[57][14] , \mult_22/ab[57][15] ,
         \mult_22/ab[57][16] , \mult_22/ab[57][17] , \mult_22/ab[57][18] ,
         \mult_22/ab[57][19] , \mult_22/ab[57][20] , \mult_22/ab[57][21] ,
         \mult_22/ab[57][22] , \mult_22/ab[57][23] , \mult_22/ab[57][24] ,
         \mult_22/ab[57][25] , \mult_22/ab[57][26] , \mult_22/ab[57][27] ,
         \mult_22/ab[57][28] , \mult_22/ab[57][29] , \mult_22/ab[57][30] ,
         \mult_22/ab[57][31] , \mult_22/ab[57][32] , \mult_22/ab[57][33] ,
         \mult_22/ab[57][34] , \mult_22/ab[57][35] , \mult_22/ab[57][36] ,
         \mult_22/ab[57][37] , \mult_22/ab[57][38] , \mult_22/ab[57][39] ,
         \mult_22/ab[57][40] , \mult_22/ab[57][41] , \mult_22/ab[57][42] ,
         \mult_22/ab[57][43] , \mult_22/ab[57][44] , \mult_22/ab[57][45] ,
         \mult_22/ab[57][46] , \mult_22/ab[57][47] , \mult_22/ab[57][48] ,
         \mult_22/ab[57][49] , \mult_22/ab[57][50] , \mult_22/ab[57][51] ,
         \mult_22/ab[57][52] , \mult_22/ab[57][53] , \mult_22/ab[57][54] ,
         \mult_22/ab[57][55] , \mult_22/ab[57][56] , \mult_22/ab[57][57] ,
         \mult_22/ab[57][58] , \mult_22/ab[57][59] , \mult_22/ab[57][60] ,
         \mult_22/ab[57][61] , \mult_22/ab[57][62] , \mult_22/ab[57][63] ,
         \mult_22/ab[58][0] , \mult_22/ab[58][1] , \mult_22/ab[58][2] ,
         \mult_22/ab[58][3] , \mult_22/ab[58][4] , \mult_22/ab[58][5] ,
         \mult_22/ab[58][6] , \mult_22/ab[58][7] , \mult_22/ab[58][8] ,
         \mult_22/ab[58][9] , \mult_22/ab[58][10] , \mult_22/ab[58][11] ,
         \mult_22/ab[58][12] , \mult_22/ab[58][13] , \mult_22/ab[58][14] ,
         \mult_22/ab[58][15] , \mult_22/ab[58][16] , \mult_22/ab[58][17] ,
         \mult_22/ab[58][18] , \mult_22/ab[58][19] , \mult_22/ab[58][20] ,
         \mult_22/ab[58][21] , \mult_22/ab[58][22] , \mult_22/ab[58][23] ,
         \mult_22/ab[58][24] , \mult_22/ab[58][25] , \mult_22/ab[58][26] ,
         \mult_22/ab[58][27] , \mult_22/ab[58][28] , \mult_22/ab[58][29] ,
         \mult_22/ab[58][30] , \mult_22/ab[58][31] , \mult_22/ab[58][32] ,
         \mult_22/ab[58][33] , \mult_22/ab[58][34] , \mult_22/ab[58][35] ,
         \mult_22/ab[58][36] , \mult_22/ab[58][37] , \mult_22/ab[58][38] ,
         \mult_22/ab[58][39] , \mult_22/ab[58][40] , \mult_22/ab[58][41] ,
         \mult_22/ab[58][42] , \mult_22/ab[58][43] , \mult_22/ab[58][44] ,
         \mult_22/ab[58][45] , \mult_22/ab[58][46] , \mult_22/ab[58][47] ,
         \mult_22/ab[58][48] , \mult_22/ab[58][49] , \mult_22/ab[58][50] ,
         \mult_22/ab[58][51] , \mult_22/ab[58][52] , \mult_22/ab[58][53] ,
         \mult_22/ab[58][54] , \mult_22/ab[58][55] , \mult_22/ab[58][56] ,
         \mult_22/ab[58][57] , \mult_22/ab[58][58] , \mult_22/ab[58][59] ,
         \mult_22/ab[58][60] , \mult_22/ab[58][61] , \mult_22/ab[58][62] ,
         \mult_22/ab[58][63] , \mult_22/ab[59][0] , \mult_22/ab[59][1] ,
         \mult_22/ab[59][2] , \mult_22/ab[59][3] , \mult_22/ab[59][4] ,
         \mult_22/ab[59][5] , \mult_22/ab[59][6] , \mult_22/ab[59][7] ,
         \mult_22/ab[59][8] , \mult_22/ab[59][9] , \mult_22/ab[59][10] ,
         \mult_22/ab[59][11] , \mult_22/ab[59][12] , \mult_22/ab[59][13] ,
         \mult_22/ab[59][14] , \mult_22/ab[59][15] , \mult_22/ab[59][16] ,
         \mult_22/ab[59][17] , \mult_22/ab[59][18] , \mult_22/ab[59][19] ,
         \mult_22/ab[59][20] , \mult_22/ab[59][21] , \mult_22/ab[59][22] ,
         \mult_22/ab[59][23] , \mult_22/ab[59][24] , \mult_22/ab[59][25] ,
         \mult_22/ab[59][26] , \mult_22/ab[59][27] , \mult_22/ab[59][28] ,
         \mult_22/ab[59][29] , \mult_22/ab[59][30] , \mult_22/ab[59][31] ,
         \mult_22/ab[59][32] , \mult_22/ab[59][33] , \mult_22/ab[59][34] ,
         \mult_22/ab[59][35] , \mult_22/ab[59][36] , \mult_22/ab[59][37] ,
         \mult_22/ab[59][38] , \mult_22/ab[59][39] , \mult_22/ab[59][40] ,
         \mult_22/ab[59][41] , \mult_22/ab[59][42] , \mult_22/ab[59][43] ,
         \mult_22/ab[59][44] , \mult_22/ab[59][45] , \mult_22/ab[59][46] ,
         \mult_22/ab[59][47] , \mult_22/ab[59][48] , \mult_22/ab[59][49] ,
         \mult_22/ab[59][50] , \mult_22/ab[59][51] , \mult_22/ab[59][52] ,
         \mult_22/ab[59][53] , \mult_22/ab[59][54] , \mult_22/ab[59][55] ,
         \mult_22/ab[59][56] , \mult_22/ab[59][57] , \mult_22/ab[59][58] ,
         \mult_22/ab[59][59] , \mult_22/ab[59][60] , \mult_22/ab[59][61] ,
         \mult_22/ab[59][62] , \mult_22/ab[59][63] , \mult_22/ab[60][0] ,
         \mult_22/ab[60][1] , \mult_22/ab[60][2] , \mult_22/ab[60][3] ,
         \mult_22/ab[60][4] , \mult_22/ab[60][5] , \mult_22/ab[60][6] ,
         \mult_22/ab[60][7] , \mult_22/ab[60][8] , \mult_22/ab[60][9] ,
         \mult_22/ab[60][10] , \mult_22/ab[60][11] , \mult_22/ab[60][12] ,
         \mult_22/ab[60][13] , \mult_22/ab[60][14] , \mult_22/ab[60][15] ,
         \mult_22/ab[60][16] , \mult_22/ab[60][17] , \mult_22/ab[60][18] ,
         \mult_22/ab[60][19] , \mult_22/ab[60][20] , \mult_22/ab[60][21] ,
         \mult_22/ab[60][22] , \mult_22/ab[60][23] , \mult_22/ab[60][24] ,
         \mult_22/ab[60][25] , \mult_22/ab[60][26] , \mult_22/ab[60][27] ,
         \mult_22/ab[60][28] , \mult_22/ab[60][29] , \mult_22/ab[60][30] ,
         \mult_22/ab[60][31] , \mult_22/ab[60][32] , \mult_22/ab[60][33] ,
         \mult_22/ab[60][34] , \mult_22/ab[60][35] , \mult_22/ab[60][36] ,
         \mult_22/ab[60][37] , \mult_22/ab[60][38] , \mult_22/ab[60][39] ,
         \mult_22/ab[60][40] , \mult_22/ab[60][41] , \mult_22/ab[60][42] ,
         \mult_22/ab[60][43] , \mult_22/ab[60][44] , \mult_22/ab[60][45] ,
         \mult_22/ab[60][46] , \mult_22/ab[60][47] , \mult_22/ab[60][48] ,
         \mult_22/ab[60][49] , \mult_22/ab[60][50] , \mult_22/ab[60][51] ,
         \mult_22/ab[60][52] , \mult_22/ab[60][53] , \mult_22/ab[60][54] ,
         \mult_22/ab[60][55] , \mult_22/ab[60][56] , \mult_22/ab[60][57] ,
         \mult_22/ab[60][58] , \mult_22/ab[60][59] , \mult_22/ab[60][60] ,
         \mult_22/ab[60][61] , \mult_22/ab[60][62] , \mult_22/ab[60][63] ,
         \mult_22/ab[61][0] , \mult_22/ab[61][1] , \mult_22/ab[61][2] ,
         \mult_22/ab[61][3] , \mult_22/ab[61][4] , \mult_22/ab[61][5] ,
         \mult_22/ab[61][6] , \mult_22/ab[61][7] , \mult_22/ab[61][8] ,
         \mult_22/ab[61][9] , \mult_22/ab[61][10] , \mult_22/ab[61][11] ,
         \mult_22/ab[61][12] , \mult_22/ab[61][13] , \mult_22/ab[61][14] ,
         \mult_22/ab[61][15] , \mult_22/ab[61][16] , \mult_22/ab[61][17] ,
         \mult_22/ab[61][18] , \mult_22/ab[61][19] , \mult_22/ab[61][20] ,
         \mult_22/ab[61][21] , \mult_22/ab[61][22] , \mult_22/ab[61][23] ,
         \mult_22/ab[61][24] , \mult_22/ab[61][25] , \mult_22/ab[61][26] ,
         \mult_22/ab[61][27] , \mult_22/ab[61][28] , \mult_22/ab[61][29] ,
         \mult_22/ab[61][30] , \mult_22/ab[61][31] , \mult_22/ab[61][32] ,
         \mult_22/ab[61][33] , \mult_22/ab[61][34] , \mult_22/ab[61][35] ,
         \mult_22/ab[61][36] , \mult_22/ab[61][37] , \mult_22/ab[61][38] ,
         \mult_22/ab[61][39] , \mult_22/ab[61][40] , \mult_22/ab[61][41] ,
         \mult_22/ab[61][42] , \mult_22/ab[61][43] , \mult_22/ab[61][44] ,
         \mult_22/ab[61][45] , \mult_22/ab[61][46] , \mult_22/ab[61][47] ,
         \mult_22/ab[61][48] , \mult_22/ab[61][49] , \mult_22/ab[61][50] ,
         \mult_22/ab[61][51] , \mult_22/ab[61][52] , \mult_22/ab[61][53] ,
         \mult_22/ab[61][54] , \mult_22/ab[61][55] , \mult_22/ab[61][56] ,
         \mult_22/ab[61][57] , \mult_22/ab[61][58] , \mult_22/ab[61][59] ,
         \mult_22/ab[61][60] , \mult_22/ab[61][61] , \mult_22/ab[61][62] ,
         \mult_22/ab[61][63] , \mult_22/ab[62][0] , \mult_22/ab[62][1] ,
         \mult_22/ab[62][2] , \mult_22/ab[62][3] , \mult_22/ab[62][4] ,
         \mult_22/ab[62][5] , \mult_22/ab[62][6] , \mult_22/ab[62][7] ,
         \mult_22/ab[62][8] , \mult_22/ab[62][9] , \mult_22/ab[62][10] ,
         \mult_22/ab[62][11] , \mult_22/ab[62][12] , \mult_22/ab[62][13] ,
         \mult_22/ab[62][14] , \mult_22/ab[62][15] , \mult_22/ab[62][16] ,
         \mult_22/ab[62][17] , \mult_22/ab[62][18] , \mult_22/ab[62][19] ,
         \mult_22/ab[62][20] , \mult_22/ab[62][21] , \mult_22/ab[62][22] ,
         \mult_22/ab[62][23] , \mult_22/ab[62][24] , \mult_22/ab[62][25] ,
         \mult_22/ab[62][26] , \mult_22/ab[62][27] , \mult_22/ab[62][28] ,
         \mult_22/ab[62][29] , \mult_22/ab[62][30] , \mult_22/ab[62][31] ,
         \mult_22/ab[62][32] , \mult_22/ab[62][33] , \mult_22/ab[62][34] ,
         \mult_22/ab[62][35] , \mult_22/ab[62][36] , \mult_22/ab[62][37] ,
         \mult_22/ab[62][38] , \mult_22/ab[62][39] , \mult_22/ab[62][40] ,
         \mult_22/ab[62][41] , \mult_22/ab[62][42] , \mult_22/ab[62][43] ,
         \mult_22/ab[62][44] , \mult_22/ab[62][45] , \mult_22/ab[62][46] ,
         \mult_22/ab[62][47] , \mult_22/ab[62][48] , \mult_22/ab[62][49] ,
         \mult_22/ab[62][50] , \mult_22/ab[62][51] , \mult_22/ab[62][52] ,
         \mult_22/ab[62][53] , \mult_22/ab[62][54] , \mult_22/ab[62][55] ,
         \mult_22/ab[62][56] , \mult_22/ab[62][57] , \mult_22/ab[62][58] ,
         \mult_22/ab[62][59] , \mult_22/ab[62][60] , \mult_22/ab[62][61] ,
         \mult_22/ab[62][62] , \mult_22/ab[62][63] , \mult_22/ab[63][0] ,
         \mult_22/ab[63][1] , \mult_22/ab[63][2] , \mult_22/ab[63][3] ,
         \mult_22/ab[63][4] , \mult_22/ab[63][5] , \mult_22/ab[63][6] ,
         \mult_22/ab[63][7] , \mult_22/ab[63][8] , \mult_22/ab[63][9] ,
         \mult_22/ab[63][10] , \mult_22/ab[63][11] , \mult_22/ab[63][12] ,
         \mult_22/ab[63][13] , \mult_22/ab[63][14] , \mult_22/ab[63][15] ,
         \mult_22/ab[63][16] , \mult_22/ab[63][17] , \mult_22/ab[63][18] ,
         \mult_22/ab[63][19] , \mult_22/ab[63][20] , \mult_22/ab[63][21] ,
         \mult_22/ab[63][22] , \mult_22/ab[63][23] , \mult_22/ab[63][24] ,
         \mult_22/ab[63][25] , \mult_22/ab[63][26] , \mult_22/ab[63][27] ,
         \mult_22/ab[63][28] , \mult_22/ab[63][29] , \mult_22/ab[63][30] ,
         \mult_22/ab[63][31] , \mult_22/ab[63][32] , \mult_22/ab[63][33] ,
         \mult_22/ab[63][34] , \mult_22/ab[63][35] , \mult_22/ab[63][36] ,
         \mult_22/ab[63][37] , \mult_22/ab[63][38] , \mult_22/ab[63][39] ,
         \mult_22/ab[63][40] , \mult_22/ab[63][41] , \mult_22/ab[63][42] ,
         \mult_22/ab[63][43] , \mult_22/ab[63][44] , \mult_22/ab[63][45] ,
         \mult_22/ab[63][46] , \mult_22/ab[63][47] , \mult_22/ab[63][48] ,
         \mult_22/ab[63][49] , \mult_22/ab[63][50] , \mult_22/ab[63][51] ,
         \mult_22/ab[63][52] , \mult_22/ab[63][53] , \mult_22/ab[63][54] ,
         \mult_22/ab[63][55] , \mult_22/ab[63][56] , \mult_22/ab[63][57] ,
         \mult_22/ab[63][58] , \mult_22/ab[63][59] , \mult_22/ab[63][60] ,
         \mult_22/ab[63][61] , \mult_22/ab[63][62] , n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n686, n687, n693,
         n694, n696, n698, n700, n701, n703, n704, n706, n708, n709, n712,
         n713, n717, n718, n726, n727, n731, n732, n737, n738, n740, n741,
         n746, n748, n751, n752, n753, n754, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n903, n905, n906, n907, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n935, n938, n939, n941, n942, n945,
         n946, n947, n948, n950, n951, n952, n953, n956, n958, n959, n960,
         n961, n962, n963, n964, n967, n968, n969, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
         n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
         n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
         n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
         n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
         n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
         n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
         n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
         n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
         n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
         n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
         n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
         n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
         n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
         n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
         n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
         n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
         n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
         n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1227, n1228,
         n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
         n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
         n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
         n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
         n1269, n1270, n1271, n1272, n1274, n1275, n1276, n1277, n1278, n1279,
         n1280, n1281, n1282, n1283, n1284, n1285, n1287, n1288, n1289, n1290,
         n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1299, n1300, n1301,
         n1302, n1304, n1305, n1306, n1307, n1308, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1320, n1321, n1322, n1323, n1325,
         n1326, n1327, n1328, n1330, n1331, n1332, n1333, n1335, n1336, n1337,
         n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
         n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
         n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
         n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
         n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
         n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1397, n1398,
         n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
         n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
         n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1437, n1438, n1439, n1440,
         n1441, n1442, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451,
         n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461,
         n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471,
         n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481,
         n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491,
         n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501,
         n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511,
         n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521,
         n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531,
         n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541,
         n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
         n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
         n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
         n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
         n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
         n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1802, n1803, n1804, n1805,
         n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815,
         n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825,
         n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835,
         n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845,
         n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855,
         n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865,
         n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875,
         n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885,
         n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895,
         n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905,
         n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915,
         n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925,
         n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935,
         n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945,
         n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955,
         n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965,
         n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975,
         n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985,
         n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995,
         n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005,
         n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015,
         n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025,
         n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035,
         n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045,
         n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2055, n2056,
         n2057, n2058, n2060, n2061, n2062, n2064, n2065, n2066, n2068, n2069,
         n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
         n2080, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
         n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
         n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
         n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
         n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
         n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
         n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
         n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
         n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170,
         n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180,
         n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190,
         n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200,
         n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
         n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220,
         n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
         n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240,
         n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250,
         n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260,
         n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270,
         n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280,
         n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290,
         n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300,
         n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310,
         n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320,
         n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330,
         n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340,
         n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350,
         n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360,
         n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370,
         n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380,
         n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390,
         n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400,
         n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410,
         n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420,
         n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430,
         n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440,
         n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450,
         n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460,
         n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470,
         n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480,
         n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490,
         n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500,
         n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510,
         n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520,
         n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530,
         n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540,
         n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550,
         n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560,
         n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570,
         n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580,
         n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590,
         n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600,
         n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610,
         n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620,
         n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630,
         n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640,
         n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650,
         n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660,
         n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670,
         n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680,
         n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690,
         n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700,
         n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710,
         n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720,
         n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730,
         n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740,
         n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750,
         n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760,
         n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770,
         n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780,
         n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790,
         n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800,
         n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810,
         n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820,
         n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830,
         n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840,
         n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850,
         n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860,
         n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870,
         n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880,
         n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890,
         n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900,
         n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910,
         n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920,
         n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930,
         n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940,
         n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950,
         n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960,
         n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970,
         n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980,
         n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990,
         n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000,
         n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010,
         n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020,
         n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030,
         n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040,
         n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050,
         n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060,
         n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070,
         n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080,
         n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090,
         n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100,
         n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110,
         n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120,
         n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130,
         n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140,
         n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150,
         n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160,
         n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170,
         n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180,
         n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190,
         n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200,
         n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210,
         n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220,
         n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230,
         n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240,
         n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250,
         n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260,
         n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270,
         n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280,
         n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290,
         n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300,
         n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310,
         n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320,
         n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330,
         n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340,
         n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350,
         n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360,
         n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370,
         n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380,
         n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390,
         n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400,
         n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410,
         n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420,
         n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430,
         n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440,
         n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450,
         n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460,
         n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470,
         n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480,
         n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490,
         n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500,
         n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510,
         n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520,
         n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530,
         n3531, n3532, n3533, n3534;
  wire   [31:0] reg_ini_0;
  wire   [31:0] reg_ini_1;
  wire   [31:0] reg_ini_2;
  wire   [31:0] reg_ini_3;
  wire   [63:0] reg_mid_0;
  wire   [63:0] reg_mid_1;

  DFF_X1 \reg_ini_3_reg[31]  ( .D(g_inA3[31]), .CK(g_inClk), .Q(reg_ini_3[31]), 
        .QN(n1902) );
  DFF_X1 \reg_ini_3_reg[30]  ( .D(g_inA3[30]), .CK(g_inClk), .Q(reg_ini_3[30]), 
        .QN(n1910) );
  DFF_X1 \reg_ini_3_reg[29]  ( .D(g_inA3[29]), .CK(g_inClk), .Q(reg_ini_3[29]), 
        .QN(n1905) );
  DFF_X1 \reg_ini_3_reg[28]  ( .D(g_inA3[28]), .CK(g_inClk), .Q(reg_ini_3[28]), 
        .QN(n1913) );
  DFF_X1 \reg_ini_3_reg[27]  ( .D(g_inA3[27]), .CK(g_inClk), .Q(reg_ini_3[27]), 
        .QN(n1912) );
  DFF_X1 \reg_ini_3_reg[26]  ( .D(g_inA3[26]), .CK(g_inClk), .Q(reg_ini_3[26]), 
        .QN(n1915) );
  DFF_X1 \reg_ini_3_reg[25]  ( .D(g_inA3[25]), .CK(g_inClk), .Q(reg_ini_3[25]), 
        .QN(n1914) );
  DFF_X1 \reg_ini_3_reg[24]  ( .D(g_inA3[24]), .CK(g_inClk), .Q(reg_ini_3[24]), 
        .QN(n1906) );
  DFF_X1 \reg_ini_3_reg[23]  ( .D(g_inA3[23]), .CK(g_inClk), .Q(reg_ini_3[23]), 
        .QN(n1901) );
  DFF_X1 \reg_ini_3_reg[22]  ( .D(g_inA3[22]), .CK(g_inClk), .Q(reg_ini_3[22]), 
        .QN(n1907) );
  DFF_X1 \reg_ini_3_reg[21]  ( .D(g_inA3[21]), .CK(g_inClk), .Q(reg_ini_3[21]), 
        .QN(n1916) );
  DFF_X1 \reg_ini_3_reg[20]  ( .D(g_inA3[20]), .CK(g_inClk), .Q(reg_ini_3[20]), 
        .QN(n1966) );
  DFF_X1 \reg_ini_3_reg[19]  ( .D(g_inA3[19]), .CK(g_inClk), .Q(reg_ini_3[19]), 
        .QN(n1963) );
  DFF_X1 \reg_ini_3_reg[18]  ( .D(g_inA3[18]), .CK(g_inClk), .Q(reg_ini_3[18]), 
        .QN(n1967) );
  DFF_X1 \reg_ini_3_reg[17]  ( .D(g_inA3[17]), .CK(g_inClk), .Q(reg_ini_3[17]), 
        .QN(n1964) );
  DFF_X1 \reg_ini_3_reg[16]  ( .D(g_inA3[16]), .CK(g_inClk), .Q(reg_ini_3[16]), 
        .QN(n1968) );
  DFF_X1 \reg_ini_3_reg[15]  ( .D(g_inA3[15]), .CK(g_inClk), .Q(reg_ini_3[15]), 
        .QN(n1965) );
  DFF_X1 \reg_ini_3_reg[14]  ( .D(g_inA3[14]), .CK(g_inClk), .Q(reg_ini_3[14]), 
        .QN(n1937) );
  DFF_X1 \reg_ini_3_reg[13]  ( .D(g_inA3[13]), .CK(g_inClk), .Q(reg_ini_3[13]), 
        .QN(n1938) );
  DFF_X1 \reg_ini_3_reg[12]  ( .D(g_inA3[12]), .CK(g_inClk), .Q(reg_ini_3[12]), 
        .QN(n1939) );
  DFF_X1 \reg_ini_3_reg[11]  ( .D(g_inA3[11]), .CK(g_inClk), .Q(reg_ini_3[11]), 
        .QN(n1940) );
  DFF_X1 \reg_ini_3_reg[10]  ( .D(g_inA3[10]), .CK(g_inClk), .Q(reg_ini_3[10]), 
        .QN(n1941) );
  DFF_X1 \reg_ini_3_reg[9]  ( .D(g_inA3[9]), .CK(g_inClk), .Q(reg_ini_3[9]), 
        .QN(n1947) );
  DFF_X1 \reg_ini_3_reg[8]  ( .D(g_inA3[8]), .CK(g_inClk), .Q(reg_ini_3[8]), 
        .QN(n1948) );
  DFF_X1 \reg_ini_3_reg[7]  ( .D(g_inA3[7]), .CK(g_inClk), .Q(reg_ini_3[7]), 
        .QN(n1949) );
  DFF_X1 \reg_ini_3_reg[6]  ( .D(g_inA3[6]), .CK(g_inClk), .Q(reg_ini_3[6]), 
        .QN(n1950) );
  DFF_X1 \reg_ini_3_reg[5]  ( .D(g_inA3[5]), .CK(g_inClk), .Q(reg_ini_3[5]), 
        .QN(n1951) );
  DFF_X1 \reg_ini_3_reg[4]  ( .D(g_inA3[4]), .CK(g_inClk), .Q(reg_ini_3[4]), 
        .QN(n1960) );
  DFF_X1 \reg_ini_3_reg[3]  ( .D(g_inA3[3]), .CK(g_inClk), .Q(reg_ini_3[3]), 
        .QN(n1961) );
  DFF_X1 \reg_ini_3_reg[2]  ( .D(g_inA3[2]), .CK(g_inClk), .Q(reg_ini_3[2]), 
        .QN(n1962) );
  DFF_X1 \reg_ini_3_reg[1]  ( .D(g_inA3[1]), .CK(g_inClk), .Q(reg_ini_3[1]), 
        .QN(n1975) );
  DFF_X1 \reg_ini_3_reg[0]  ( .D(g_inA3[0]), .CK(g_inClk), .Q(reg_ini_3[0]), 
        .QN(n1977) );
  DFF_X1 \reg_ini_2_reg[31]  ( .D(g_inA2[31]), .CK(g_inClk), .Q(reg_ini_2[31]), 
        .QN(n2044) );
  DFF_X1 \reg_ini_2_reg[30]  ( .D(g_inA2[30]), .CK(g_inClk), .Q(reg_ini_2[30]), 
        .QN(n2050) );
  DFF_X1 \reg_ini_2_reg[29]  ( .D(g_inA2[29]), .CK(g_inClk), .Q(reg_ini_2[29]), 
        .QN(n2048) );
  DFF_X1 \reg_ini_2_reg[28]  ( .D(g_inA2[28]), .CK(g_inClk), .Q(reg_ini_2[28]), 
        .QN(n2046) );
  DFF_X1 \reg_ini_2_reg[27]  ( .D(g_inA2[27]), .CK(g_inClk), .Q(reg_ini_2[27]), 
        .QN(n2042) );
  DFF_X1 \reg_ini_2_reg[26]  ( .D(g_inA2[26]), .CK(g_inClk), .Q(reg_ini_2[26]), 
        .QN(n2040) );
  DFF_X1 \reg_ini_2_reg[25]  ( .D(g_inA2[25]), .CK(g_inClk), .Q(reg_ini_2[25]), 
        .QN(n2038) );
  DFF_X1 \reg_ini_2_reg[24]  ( .D(g_inA2[24]), .CK(g_inClk), .Q(reg_ini_2[24]), 
        .QN(n2036) );
  DFF_X1 \reg_ini_2_reg[23]  ( .D(g_inA2[23]), .CK(g_inClk), .Q(reg_ini_2[23]), 
        .QN(n2034) );
  DFF_X1 \reg_ini_2_reg[22]  ( .D(g_inA2[22]), .CK(g_inClk), .Q(reg_ini_2[22]), 
        .QN(n2032) );
  DFF_X1 \reg_ini_2_reg[21]  ( .D(g_inA2[21]), .CK(g_inClk), .Q(reg_ini_2[21]), 
        .QN(n2030) );
  DFF_X1 \reg_ini_2_reg[20]  ( .D(g_inA2[20]), .CK(g_inClk), .Q(reg_ini_2[20]), 
        .QN(n2028) );
  DFF_X1 \reg_ini_2_reg[19]  ( .D(g_inA2[19]), .CK(g_inClk), .Q(reg_ini_2[19]), 
        .QN(n2018) );
  DFF_X1 \reg_ini_2_reg[18]  ( .D(g_inA2[18]), .CK(g_inClk), .Q(reg_ini_2[18]), 
        .QN(n2016) );
  DFF_X1 \reg_ini_2_reg[17]  ( .D(g_inA2[17]), .CK(g_inClk), .Q(reg_ini_2[17]), 
        .QN(n2014) );
  DFF_X1 \reg_ini_2_reg[16]  ( .D(g_inA2[16]), .CK(g_inClk), .Q(reg_ini_2[16]), 
        .QN(n2012) );
  DFF_X1 \reg_ini_2_reg[15]  ( .D(g_inA2[15]), .CK(g_inClk), .Q(reg_ini_2[15]), 
        .QN(n2010) );
  DFF_X1 \reg_ini_2_reg[14]  ( .D(g_inA2[14]), .CK(g_inClk), .Q(reg_ini_2[14]), 
        .QN(n2008) );
  DFF_X1 \reg_ini_2_reg[13]  ( .D(g_inA2[13]), .CK(g_inClk), .Q(reg_ini_2[13]), 
        .QN(n2006) );
  DFF_X1 \reg_ini_2_reg[12]  ( .D(g_inA2[12]), .CK(g_inClk), .Q(reg_ini_2[12]), 
        .QN(n2004) );
  DFF_X1 \reg_ini_2_reg[11]  ( .D(g_inA2[11]), .CK(g_inClk), .Q(reg_ini_2[11]), 
        .QN(n1984) );
  DFF_X1 \reg_ini_2_reg[10]  ( .D(g_inA2[10]), .CK(g_inClk), .Q(reg_ini_2[10]), 
        .QN(n1983) );
  DFF_X1 \reg_ini_2_reg[9]  ( .D(g_inA2[9]), .CK(g_inClk), .Q(reg_ini_2[9]), 
        .QN(n1982) );
  DFF_X1 \reg_ini_2_reg[8]  ( .D(g_inA2[8]), .CK(g_inClk), .Q(reg_ini_2[8]), 
        .QN(n1981) );
  DFF_X1 \reg_ini_2_reg[7]  ( .D(g_inA2[7]), .CK(g_inClk), .Q(reg_ini_2[7]), 
        .QN(n1980) );
  DFF_X1 \reg_ini_2_reg[6]  ( .D(g_inA2[6]), .CK(g_inClk), .Q(reg_ini_2[6]), 
        .QN(n1979) );
  DFF_X1 \reg_ini_2_reg[5]  ( .D(g_inA2[5]), .CK(g_inClk), .Q(reg_ini_2[5]), 
        .QN(n1992) );
  DFF_X1 \reg_ini_2_reg[4]  ( .D(g_inA2[4]), .CK(g_inClk), .Q(reg_ini_2[4]), 
        .QN(n1991) );
  DFF_X1 \reg_ini_2_reg[3]  ( .D(g_inA2[3]), .CK(g_inClk), .Q(reg_ini_2[3]), 
        .QN(n1923) );
  DFF_X1 \reg_ini_2_reg[2]  ( .D(g_inA2[2]), .CK(g_inClk), .Q(reg_ini_2[2]), 
        .QN(n1925) );
  DFF_X1 \reg_ini_2_reg[1]  ( .D(g_inA2[1]), .CK(g_inClk), .Q(n1806), .QN(
        n1807) );
  DFF_X1 \reg_ini_2_reg[0]  ( .D(g_inA2[0]), .CK(g_inClk), .Q(reg_ini_2[0]), 
        .QN(n1935) );
  DFF_X1 \reg_ini_1_reg[31]  ( .D(g_inA1[31]), .CK(g_inClk), .Q(reg_ini_1[31]), 
        .QN(n1903) );
  DFF_X1 \reg_ini_1_reg[30]  ( .D(g_inA1[30]), .CK(g_inClk), .Q(reg_ini_1[30]), 
        .QN(n1911) );
  DFF_X1 \reg_ini_1_reg[29]  ( .D(g_inA1[29]), .CK(g_inClk), .Q(reg_ini_1[29]), 
        .QN(n1908) );
  DFF_X1 \reg_ini_1_reg[28]  ( .D(g_inA1[28]), .CK(g_inClk), .Q(reg_ini_1[28]), 
        .QN(n1917) );
  DFF_X1 \reg_ini_1_reg[27]  ( .D(g_inA1[27]), .CK(g_inClk), .Q(reg_ini_1[27]), 
        .QN(n1918) );
  DFF_X1 \reg_ini_1_reg[26]  ( .D(g_inA1[26]), .CK(g_inClk), .Q(reg_ini_1[26]), 
        .QN(n1920) );
  DFF_X1 \reg_ini_1_reg[25]  ( .D(g_inA1[25]), .CK(g_inClk), .Q(reg_ini_1[25]), 
        .QN(n1919) );
  DFF_X1 \reg_ini_1_reg[24]  ( .D(g_inA1[24]), .CK(g_inClk), .Q(reg_ini_1[24]), 
        .QN(n1921) );
  DFF_X1 \reg_ini_1_reg[23]  ( .D(g_inA1[23]), .CK(g_inClk), .Q(reg_ini_1[23]), 
        .QN(n1904) );
  DFF_X1 \reg_ini_1_reg[22]  ( .D(g_inA1[22]), .CK(g_inClk), .Q(reg_ini_1[22]), 
        .QN(n1909) );
  DFF_X1 \reg_ini_1_reg[21]  ( .D(g_inA1[21]), .CK(g_inClk), .Q(reg_ini_1[21]), 
        .QN(n1922) );
  DFF_X1 \reg_ini_1_reg[20]  ( .D(g_inA1[20]), .CK(g_inClk), .Q(reg_ini_1[20]), 
        .QN(n1969) );
  DFF_X1 \reg_ini_1_reg[19]  ( .D(g_inA1[19]), .CK(g_inClk), .Q(reg_ini_1[19]), 
        .QN(n1970) );
  DFF_X1 \reg_ini_1_reg[18]  ( .D(g_inA1[18]), .CK(g_inClk), .Q(reg_ini_1[18]), 
        .QN(n1971) );
  DFF_X1 \reg_ini_1_reg[17]  ( .D(g_inA1[17]), .CK(g_inClk), .Q(reg_ini_1[17]), 
        .QN(n1972) );
  DFF_X1 \reg_ini_1_reg[16]  ( .D(g_inA1[16]), .CK(g_inClk), .Q(reg_ini_1[16]), 
        .QN(n1973) );
  DFF_X1 \reg_ini_1_reg[15]  ( .D(g_inA1[15]), .CK(g_inClk), .Q(reg_ini_1[15]), 
        .QN(n1974) );
  DFF_X1 \reg_ini_1_reg[14]  ( .D(g_inA1[14]), .CK(g_inClk), .Q(reg_ini_1[14]), 
        .QN(n1942) );
  DFF_X1 \reg_ini_1_reg[13]  ( .D(g_inA1[13]), .CK(g_inClk), .Q(reg_ini_1[13]), 
        .QN(n1943) );
  DFF_X1 \reg_ini_1_reg[12]  ( .D(g_inA1[12]), .CK(g_inClk), .Q(reg_ini_1[12]), 
        .QN(n1944) );
  DFF_X1 \reg_ini_1_reg[11]  ( .D(g_inA1[11]), .CK(g_inClk), .Q(reg_ini_1[11]), 
        .QN(n1945) );
  DFF_X1 \reg_ini_1_reg[10]  ( .D(g_inA1[10]), .CK(g_inClk), .Q(reg_ini_1[10]), 
        .QN(n1946) );
  DFF_X1 \reg_ini_1_reg[9]  ( .D(g_inA1[9]), .CK(g_inClk), .Q(reg_ini_1[9]), 
        .QN(n1955) );
  DFF_X1 \reg_ini_1_reg[8]  ( .D(g_inA1[8]), .CK(g_inClk), .Q(reg_ini_1[8]), 
        .QN(n1956) );
  DFF_X1 \reg_ini_1_reg[7]  ( .D(g_inA1[7]), .CK(g_inClk), .Q(reg_ini_1[7]), 
        .QN(n1957) );
  DFF_X1 \reg_ini_1_reg[6]  ( .D(g_inA1[6]), .CK(g_inClk), .Q(reg_ini_1[6]), 
        .QN(n1958) );
  DFF_X1 \reg_ini_1_reg[5]  ( .D(g_inA1[5]), .CK(g_inClk), .Q(reg_ini_1[5]), 
        .QN(n1959) );
  DFF_X1 \reg_ini_1_reg[4]  ( .D(g_inA1[4]), .CK(g_inClk), .Q(reg_ini_1[4]), 
        .QN(n1952) );
  DFF_X1 \reg_ini_1_reg[3]  ( .D(g_inA1[3]), .CK(g_inClk), .Q(reg_ini_1[3]), 
        .QN(n1953) );
  DFF_X1 \reg_ini_1_reg[2]  ( .D(g_inA1[2]), .CK(g_inClk), .Q(reg_ini_1[2]), 
        .QN(n1954) );
  DFF_X1 \reg_ini_1_reg[1]  ( .D(g_inA1[1]), .CK(g_inClk), .Q(reg_ini_1[1]), 
        .QN(n1976) );
  DFF_X1 \reg_ini_1_reg[0]  ( .D(g_inA1[0]), .CK(g_inClk), .Q(reg_ini_1[0]), 
        .QN(n1978) );
  DFF_X1 \reg_ini_0_reg[31]  ( .D(g_inA0[31]), .CK(g_inClk), .Q(reg_ini_0[31]), 
        .QN(n2045) );
  DFF_X1 \reg_ini_0_reg[30]  ( .D(g_inA0[30]), .CK(g_inClk), .Q(reg_ini_0[30]), 
        .QN(n2051) );
  DFF_X1 \reg_ini_0_reg[29]  ( .D(g_inA0[29]), .CK(g_inClk), .Q(reg_ini_0[29]), 
        .QN(n2049) );
  DFF_X1 \reg_ini_0_reg[28]  ( .D(g_inA0[28]), .CK(g_inClk), .Q(reg_ini_0[28]), 
        .QN(n2047) );
  DFF_X1 \reg_ini_0_reg[27]  ( .D(g_inA0[27]), .CK(g_inClk), .Q(reg_ini_0[27]), 
        .QN(n2043) );
  DFF_X1 \reg_ini_0_reg[26]  ( .D(g_inA0[26]), .CK(g_inClk), .Q(reg_ini_0[26]), 
        .QN(n2041) );
  DFF_X1 \reg_ini_0_reg[25]  ( .D(g_inA0[25]), .CK(g_inClk), .Q(reg_ini_0[25]), 
        .QN(n2039) );
  DFF_X1 \reg_ini_0_reg[24]  ( .D(g_inA0[24]), .CK(g_inClk), .Q(reg_ini_0[24]), 
        .QN(n2037) );
  DFF_X1 \reg_ini_0_reg[23]  ( .D(g_inA0[23]), .CK(g_inClk), .Q(reg_ini_0[23]), 
        .QN(n2035) );
  DFF_X1 \reg_ini_0_reg[22]  ( .D(g_inA0[22]), .CK(g_inClk), .Q(reg_ini_0[22]), 
        .QN(n2033) );
  DFF_X1 \reg_ini_0_reg[21]  ( .D(g_inA0[21]), .CK(g_inClk), .Q(reg_ini_0[21]), 
        .QN(n2031) );
  DFF_X1 \reg_ini_0_reg[20]  ( .D(g_inA0[20]), .CK(g_inClk), .Q(reg_ini_0[20]), 
        .QN(n2029) );
  DFF_X1 \reg_ini_0_reg[19]  ( .D(g_inA0[19]), .CK(g_inClk), .Q(reg_ini_0[19]), 
        .QN(n2019) );
  DFF_X1 \reg_ini_0_reg[18]  ( .D(g_inA0[18]), .CK(g_inClk), .Q(reg_ini_0[18]), 
        .QN(n2017) );
  DFF_X1 \reg_ini_0_reg[17]  ( .D(g_inA0[17]), .CK(g_inClk), .Q(reg_ini_0[17]), 
        .QN(n2015) );
  DFF_X1 \reg_ini_0_reg[16]  ( .D(g_inA0[16]), .CK(g_inClk), .Q(reg_ini_0[16]), 
        .QN(n2013) );
  DFF_X1 \reg_ini_0_reg[15]  ( .D(g_inA0[15]), .CK(g_inClk), .Q(reg_ini_0[15]), 
        .QN(n2011) );
  DFF_X1 \reg_ini_0_reg[14]  ( .D(g_inA0[14]), .CK(g_inClk), .Q(reg_ini_0[14]), 
        .QN(n2009) );
  DFF_X1 \reg_ini_0_reg[13]  ( .D(g_inA0[13]), .CK(g_inClk), .Q(reg_ini_0[13]), 
        .QN(n2007) );
  DFF_X1 \reg_ini_0_reg[12]  ( .D(g_inA0[12]), .CK(g_inClk), .Q(reg_ini_0[12]), 
        .QN(n2005) );
  DFF_X1 \reg_ini_0_reg[11]  ( .D(g_inA0[11]), .CK(g_inClk), .Q(reg_ini_0[11]), 
        .QN(n1990) );
  DFF_X1 \reg_ini_0_reg[10]  ( .D(g_inA0[10]), .CK(g_inClk), .Q(reg_ini_0[10]), 
        .QN(n1989) );
  DFF_X1 \reg_ini_0_reg[9]  ( .D(g_inA0[9]), .CK(g_inClk), .Q(reg_ini_0[9]), 
        .QN(n1988) );
  DFF_X1 \reg_ini_0_reg[8]  ( .D(g_inA0[8]), .CK(g_inClk), .Q(reg_ini_0[8]), 
        .QN(n1987) );
  DFF_X1 \reg_ini_0_reg[7]  ( .D(g_inA0[7]), .CK(g_inClk), .Q(reg_ini_0[7]), 
        .QN(n1986) );
  DFF_X1 \reg_ini_0_reg[6]  ( .D(g_inA0[6]), .CK(g_inClk), .Q(reg_ini_0[6]), 
        .QN(n1985) );
  DFF_X1 \reg_ini_0_reg[5]  ( .D(g_inA0[5]), .CK(g_inClk), .Q(reg_ini_0[5]), 
        .QN(n1994) );
  DFF_X1 \reg_ini_0_reg[4]  ( .D(g_inA0[4]), .CK(g_inClk), .Q(reg_ini_0[4]), 
        .QN(n1993) );
  DFF_X1 \reg_ini_0_reg[3]  ( .D(g_inA0[3]), .CK(g_inClk), .Q(reg_ini_0[3]), 
        .QN(n1924) );
  DFF_X1 \reg_ini_0_reg[2]  ( .D(g_inA0[2]), .CK(g_inClk), .Q(reg_ini_0[2]), 
        .QN(n1926) );
  DFF_X1 \reg_ini_0_reg[1]  ( .D(g_inA0[1]), .CK(g_inClk), .Q(n1805), .QN(
        n1808) );
  DFF_X1 \reg_ini_0_reg[0]  ( .D(g_inA0[0]), .CK(g_inClk), .Q(reg_ini_0[0]), 
        .QN(n1936) );
  DFF_X1 \reg_mid_0_reg[63]  ( .D(N63), .CK(g_inClk), .Q(reg_mid_0[63]), .QN(
        n2022) );
  DFF_X1 \reg_mid_0_reg[62]  ( .D(N62), .CK(g_inClk), .Q(reg_mid_0[62]), .QN(
        n2023) );
  DFF_X1 \reg_mid_0_reg[61]  ( .D(N61), .CK(g_inClk), .Q(reg_mid_0[61]), .QN(
        n2024) );
  DFF_X1 \reg_mid_0_reg[60]  ( .D(N60), .CK(g_inClk), .Q(reg_mid_0[60]), .QN(
        n2025) );
  DFF_X1 \reg_mid_0_reg[59]  ( .D(N59), .CK(g_inClk), .Q(reg_mid_0[59]), .QN(
        n2026) );
  DFF_X1 \reg_mid_0_reg[58]  ( .D(N58), .CK(g_inClk), .Q(reg_mid_0[58]), .QN(
        n2027) );
  DFF_X1 \reg_mid_0_reg[57]  ( .D(N57), .CK(g_inClk), .Q(reg_mid_0[57]), .QN(
        n2020) );
  DFF_X1 \reg_mid_0_reg[56]  ( .D(N56), .CK(g_inClk), .Q(reg_mid_0[56]), .QN(
        n2021) );
  DFF_X1 \reg_mid_0_reg[55]  ( .D(N55), .CK(g_inClk), .Q(reg_mid_0[55]), .QN(
        n2002) );
  DFF_X1 \reg_mid_0_reg[54]  ( .D(N54), .CK(g_inClk), .Q(reg_mid_0[54]), .QN(
        n2003) );
  DFF_X1 \reg_mid_0_reg[53]  ( .D(N53), .CK(g_inClk), .Q(reg_mid_0[53]), .QN(
        n2001) );
  DFF_X1 \reg_mid_0_reg[52]  ( .D(N52), .CK(g_inClk), .Q(reg_mid_0[52]), .QN(
        n2000) );
  DFF_X1 \reg_mid_0_reg[51]  ( .D(N51), .CK(g_inClk), .Q(reg_mid_0[51]), .QN(
        n1999) );
  DFF_X1 \reg_mid_0_reg[50]  ( .D(N50), .CK(g_inClk), .Q(reg_mid_0[50]), .QN(
        n1998) );
  DFF_X1 \reg_mid_0_reg[49]  ( .D(N49), .CK(g_inClk), .Q(reg_mid_0[49]), .QN(
        n1996) );
  DFF_X1 \reg_mid_0_reg[48]  ( .D(N48), .CK(g_inClk), .Q(reg_mid_0[48]), .QN(
        n1997) );
  DFF_X1 \reg_mid_0_reg[47]  ( .D(N47), .CK(g_inClk), .Q(reg_mid_0[47]), .QN(
        n1995) );
  DFF_X1 \reg_mid_0_reg[46]  ( .D(N46), .CK(g_inClk), .Q(reg_mid_0[46]), .QN(
        n1933) );
  DFF_X1 \reg_mid_0_reg[45]  ( .D(N45), .CK(g_inClk), .Q(reg_mid_0[45]), .QN(
        n1934) );
  DFF_X1 \reg_mid_0_reg[44]  ( .D(N44), .CK(g_inClk), .Q(reg_mid_0[44]), .QN(
        n1932) );
  DFF_X1 \reg_mid_0_reg[43]  ( .D(N43), .CK(g_inClk), .Q(reg_mid_0[43]), .QN(
        n1931) );
  DFF_X1 \reg_mid_0_reg[42]  ( .D(N42), .CK(g_inClk), .Q(reg_mid_0[42]), .QN(
        n1930) );
  DFF_X1 \reg_mid_0_reg[41]  ( .D(N41), .CK(g_inClk), .Q(reg_mid_0[41]), .QN(
        n1929) );
  DFF_X1 \reg_mid_0_reg[40]  ( .D(N40), .CK(g_inClk), .Q(reg_mid_0[40]), .QN(
        n1928) );
  DFF_X1 \reg_mid_0_reg[39]  ( .D(N39), .CK(g_inClk), .Q(reg_mid_0[39]), .QN(
        n1927) );
  DFF_X1 \reg_mid_0_reg[38]  ( .D(N38), .CK(g_inClk), .Q(reg_mid_0[38]), .QN(
        n1896) );
  DFF_X1 \reg_mid_0_reg[37]  ( .D(N37), .CK(g_inClk), .Q(reg_mid_0[37]), .QN(
        n1895) );
  DFF_X1 \reg_mid_0_reg[36]  ( .D(N36), .CK(g_inClk), .Q(reg_mid_0[36]), .QN(
        n1894) );
  DFF_X1 \reg_mid_0_reg[35]  ( .D(N35), .CK(g_inClk), .Q(reg_mid_0[35]), .QN(
        n1897) );
  DFF_X1 \reg_mid_0_reg[34]  ( .D(N34), .CK(g_inClk), .Q(reg_mid_0[34]), .QN(
        n1898) );
  DFF_X1 \reg_mid_0_reg[33]  ( .D(N33), .CK(g_inClk), .Q(reg_mid_0[33]), .QN(
        n1899) );
  DFF_X1 \reg_mid_0_reg[32]  ( .D(N32), .CK(g_inClk), .Q(reg_mid_0[32]), .QN(
        n1888) );
  DFF_X1 \reg_mid_0_reg[31]  ( .D(N31), .CK(g_inClk), .Q(reg_mid_0[31]), .QN(
        n1900) );
  DFF_X1 \reg_mid_0_reg[30]  ( .D(N30), .CK(g_inClk), .Q(reg_mid_0[30]), .QN(
        n1889) );
  DFF_X1 \reg_mid_0_reg[29]  ( .D(N29), .CK(g_inClk), .Q(reg_mid_0[29]), .QN(
        n1890) );
  DFF_X1 \reg_mid_0_reg[28]  ( .D(N28), .CK(g_inClk), .Q(reg_mid_0[28]), .QN(
        n1891) );
  DFF_X1 \reg_mid_0_reg[27]  ( .D(N27), .CK(g_inClk), .Q(reg_mid_0[27]), .QN(
        n1892) );
  DFF_X1 \reg_mid_0_reg[26]  ( .D(N26), .CK(g_inClk), .Q(reg_mid_0[26]), .QN(
        n1860) );
  DFF_X1 \reg_mid_0_reg[25]  ( .D(N25), .CK(g_inClk), .Q(reg_mid_0[25]), .QN(
        n1893) );
  DFF_X1 \reg_mid_0_reg[24]  ( .D(N24), .CK(g_inClk), .Q(reg_mid_0[24]), .QN(
        n1886) );
  DFF_X1 \reg_mid_0_reg[23]  ( .D(N23), .CK(g_inClk), .Q(reg_mid_0[23]), .QN(
        n1887) );
  DFF_X1 \reg_mid_0_reg[22]  ( .D(N22), .CK(g_inClk), .Q(reg_mid_0[22]), .QN(
        n1858) );
  DFF_X1 \reg_mid_0_reg[21]  ( .D(N21), .CK(g_inClk), .Q(reg_mid_0[21]), .QN(
        n1857) );
  DFF_X1 \reg_mid_0_reg[20]  ( .D(N20), .CK(g_inClk), .Q(reg_mid_0[20]), .QN(
        n1859) );
  DFF_X1 \reg_mid_0_reg[19]  ( .D(N19), .CK(g_inClk), .Q(reg_mid_0[19]), .QN(
        n1852) );
  DFF_X1 \reg_mid_0_reg[18]  ( .D(N18), .CK(g_inClk), .Q(reg_mid_0[18]), .QN(
        n1869) );
  DFF_X1 \reg_mid_0_reg[17]  ( .D(N17), .CK(g_inClk), .Q(reg_mid_0[17]), .QN(
        n1870) );
  DFF_X1 \reg_mid_0_reg[16]  ( .D(N16), .CK(g_inClk), .Q(reg_mid_0[16]), .QN(
        n1867) );
  DFF_X1 \reg_mid_0_reg[15]  ( .D(N15), .CK(g_inClk), .Q(reg_mid_0[15]), .QN(
        n1848) );
  DFF_X1 \reg_mid_0_reg[14]  ( .D(N14), .CK(g_inClk), .Q(reg_mid_0[14]), .QN(
        n1849) );
  DFF_X1 \reg_mid_0_reg[13]  ( .D(N13), .CK(g_inClk), .Q(reg_mid_0[13]), .QN(
        n1850) );
  DFF_X1 \reg_mid_0_reg[12]  ( .D(N12), .CK(g_inClk), .Q(reg_mid_0[12]), .QN(
        n1851) );
  DFF_X1 \reg_mid_0_reg[11]  ( .D(N11), .CK(g_inClk), .Q(reg_mid_0[11]), .QN(
        n1871) );
  DFF_X1 \reg_mid_0_reg[10]  ( .D(N10), .CK(g_inClk), .Q(reg_mid_0[10]), .QN(
        n1872) );
  DFF_X1 \reg_mid_0_reg[9]  ( .D(N9), .CK(g_inClk), .Q(reg_mid_0[9]), .QN(
        n1866) );
  DFF_X1 \reg_mid_0_reg[8]  ( .D(N8), .CK(g_inClk), .Q(reg_mid_0[8]), .QN(
        n1877) );
  DFF_X1 \reg_mid_0_reg[7]  ( .D(N7), .CK(g_inClk), .Q(reg_mid_0[7]), .QN(
        n1878) );
  DFF_X1 \reg_mid_0_reg[6]  ( .D(N6), .CK(g_inClk), .Q(reg_mid_0[6]), .QN(
        n1828) );
  DFF_X1 \reg_mid_0_reg[5]  ( .D(N5), .CK(g_inClk), .Q(reg_mid_0[5]), .QN(
        n1829) );
  DFF_X1 \reg_mid_0_reg[4]  ( .D(N4), .CK(g_inClk), .Q(reg_mid_0[4]), .QN(
        n1827) );
  DFF_X1 \reg_mid_0_reg[3]  ( .D(N3), .CK(g_inClk), .Q(reg_mid_0[3]), .QN(
        n1810) );
  DFF_X1 \reg_mid_0_reg[2]  ( .D(N2), .CK(g_inClk), .Q(reg_mid_0[2]), .QN(
        n2152) );
  DFF_X1 \reg_mid_1_reg[63]  ( .D(N127), .CK(g_inClk), .Q(reg_mid_1[63]), .QN(
        n2111) );
  DFF_X1 \reg_mid_1_reg[62]  ( .D(N126), .CK(g_inClk), .Q(reg_mid_1[62]), .QN(
        n2193) );
  DFF_X1 \reg_mid_1_reg[61]  ( .D(N125), .CK(g_inClk), .Q(reg_mid_1[61]), .QN(
        n2158) );
  DFF_X1 \reg_mid_1_reg[60]  ( .D(N124), .CK(g_inClk), .Q(reg_mid_1[60]), .QN(
        n2238) );
  DFF_X1 \reg_mid_1_reg[59]  ( .D(N123), .CK(g_inClk), .Q(reg_mid_1[59]), .QN(
        n2140) );
  DFF_X1 \reg_mid_1_reg[58]  ( .D(N122), .CK(g_inClk), .Q(reg_mid_1[58]), .QN(
        n1822) );
  DFF_X1 \reg_mid_1_reg[57]  ( .D(N121), .CK(g_inClk), .Q(reg_mid_1[57]), .QN(
        n2372) );
  DFF_X1 \reg_mid_1_reg[56]  ( .D(N120), .CK(g_inClk), .Q(reg_mid_1[56]), .QN(
        n2375) );
  DFF_X1 \reg_mid_1_reg[55]  ( .D(N119), .CK(g_inClk), .Q(reg_mid_1[55]), .QN(
        n2376) );
  DFF_X1 \reg_mid_1_reg[54]  ( .D(N118), .CK(g_inClk), .Q(reg_mid_1[54]), .QN(
        n2370) );
  DFF_X1 \reg_mid_1_reg[53]  ( .D(N117), .CK(g_inClk), .Q(reg_mid_1[53]), .QN(
        n1809) );
  DFF_X1 \reg_mid_1_reg[52]  ( .D(N116), .CK(g_inClk), .Q(reg_mid_1[52]), .QN(
        n1881) );
  DFF_X1 \reg_mid_1_reg[51]  ( .D(N115), .CK(g_inClk), .Q(reg_mid_1[51]), .QN(
        n1821) );
  DFF_X1 \reg_mid_1_reg[50]  ( .D(N114), .CK(g_inClk), .Q(reg_mid_1[50]), .QN(
        n2359) );
  DFF_X1 \reg_mid_1_reg[49]  ( .D(N113), .CK(g_inClk), .Q(reg_mid_1[49]), .QN(
        n1826) );
  DFF_X1 \reg_mid_1_reg[48]  ( .D(N112), .CK(g_inClk), .Q(reg_mid_1[48]), .QN(
        n2360) );
  DFF_X1 \reg_mid_1_reg[47]  ( .D(N111), .CK(g_inClk), .Q(reg_mid_1[47]), .QN(
        n2361) );
  DFF_X1 \reg_mid_1_reg[46]  ( .D(N110), .CK(g_inClk), .Q(reg_mid_1[46]), .QN(
        n2363) );
  DFF_X1 \reg_mid_1_reg[45]  ( .D(N109), .CK(g_inClk), .Q(reg_mid_1[45]), .QN(
        n2362) );
  DFF_X1 \reg_mid_1_reg[44]  ( .D(N108), .CK(g_inClk), .Q(reg_mid_1[44]), .QN(
        n1813) );
  DFF_X1 \reg_mid_1_reg[43]  ( .D(N107), .CK(g_inClk), .Q(reg_mid_1[43]), .QN(
        n1825) );
  DFF_X1 \reg_mid_1_reg[42]  ( .D(N106), .CK(g_inClk), .Q(reg_mid_1[42]), .QN(
        n1818) );
  DFF_X1 \reg_mid_1_reg[41]  ( .D(N105), .CK(g_inClk), .Q(reg_mid_1[41]), .QN(
        n1824) );
  DFF_X1 \reg_mid_1_reg[40]  ( .D(N104), .CK(g_inClk), .Q(reg_mid_1[40]), .QN(
        n1812) );
  DFF_X1 \reg_mid_1_reg[39]  ( .D(N103), .CK(g_inClk), .Q(reg_mid_1[39]), .QN(
        n1820) );
  DFF_X1 \reg_mid_1_reg[38]  ( .D(N102), .CK(g_inClk), .Q(reg_mid_1[38]), .QN(
        n1882) );
  DFF_X1 \reg_mid_1_reg[37]  ( .D(N101), .CK(g_inClk), .Q(reg_mid_1[37]), .QN(
        n1814) );
  DFF_X1 \reg_mid_1_reg[36]  ( .D(N100), .CK(g_inClk), .Q(reg_mid_1[36]), .QN(
        n1815) );
  DFF_X1 \reg_mid_1_reg[35]  ( .D(N99), .CK(g_inClk), .Q(reg_mid_1[35]), .QN(
        n1811) );
  DFF_X1 \reg_mid_1_reg[34]  ( .D(N98), .CK(g_inClk), .Q(reg_mid_1[34]), .QN(
        n1819) );
  DFF_X1 \reg_mid_1_reg[33]  ( .D(N97), .CK(g_inClk), .Q(reg_mid_1[33]), .QN(
        n1817) );
  DFF_X1 \reg_mid_1_reg[32]  ( .D(N96), .CK(g_inClk), .Q(reg_mid_1[32]), .QN(
        n1883) );
  DFF_X1 \reg_mid_1_reg[31]  ( .D(N95), .CK(g_inClk), .Q(reg_mid_1[31]), .QN(
        n1816) );
  DFF_X1 \reg_mid_1_reg[30]  ( .D(N94), .CK(g_inClk), .Q(reg_mid_1[30]), .QN(
        n1823) );
  DFF_X1 \reg_mid_1_reg[29]  ( .D(N93), .CK(g_inClk), .Q(reg_mid_1[29]), .QN(
        n1856) );
  DFF_X1 \reg_mid_1_reg[28]  ( .D(N92), .CK(g_inClk), .Q(reg_mid_1[28]), .QN(
        n1868) );
  DFF_X1 \reg_mid_1_reg[27]  ( .D(N91), .CK(g_inClk), .Q(reg_mid_1[27]), .QN(
        n1865) );
  DFF_X1 \reg_mid_1_reg[26]  ( .D(N90), .CK(g_inClk), .Q(reg_mid_1[26]), .QN(
        n1862) );
  DFF_X1 \reg_mid_1_reg[25]  ( .D(N89), .CK(g_inClk), .Q(reg_mid_1[25]), .QN(
        n1864) );
  DFF_X1 \reg_mid_1_reg[24]  ( .D(N88), .CK(g_inClk), .Q(reg_mid_1[24]), .QN(
        n1873) );
  DFF_X1 \reg_mid_1_reg[23]  ( .D(N87), .CK(g_inClk), .Q(reg_mid_1[23]), .QN(
        n1833) );
  DFF_X1 \reg_mid_1_reg[22]  ( .D(N86), .CK(g_inClk), .Q(reg_mid_1[22]), .QN(
        n1834) );
  DFF_X1 \reg_mid_1_reg[21]  ( .D(N85), .CK(g_inClk), .Q(reg_mid_1[21]), .QN(
        n1838) );
  DFF_X1 \reg_mid_1_reg[20]  ( .D(N84), .CK(g_inClk), .Q(reg_mid_1[20]), .QN(
        n1839) );
  DFF_X1 \reg_mid_1_reg[19]  ( .D(N83), .CK(g_inClk), .Q(reg_mid_1[19]), .QN(
        n1840) );
  DFF_X1 \reg_mid_1_reg[18]  ( .D(N82), .CK(g_inClk), .Q(reg_mid_1[18]), .QN(
        n1841) );
  DFF_X1 \reg_mid_1_reg[17]  ( .D(N81), .CK(g_inClk), .Q(reg_mid_1[17]), .QN(
        n1842) );
  DFF_X1 \reg_mid_1_reg[16]  ( .D(N80), .CK(g_inClk), .Q(reg_mid_1[16]), .QN(
        n1836) );
  DFF_X1 \reg_mid_1_reg[15]  ( .D(N79), .CK(g_inClk), .Q(reg_mid_1[15]), .QN(
        n1835) );
  DFF_X1 \reg_mid_1_reg[14]  ( .D(N78), .CK(g_inClk), .Q(reg_mid_1[14]), .QN(
        n1843) );
  DFF_X1 \reg_mid_1_reg[13]  ( .D(N77), .CK(g_inClk), .Q(reg_mid_1[13]), .QN(
        n1837) );
  DFF_X1 \reg_mid_1_reg[12]  ( .D(N76), .CK(g_inClk), .Q(reg_mid_1[12]), .QN(
        n1863) );
  DFF_X1 \reg_mid_1_reg[11]  ( .D(N75), .CK(g_inClk), .Q(reg_mid_1[11]), .QN(
        n1861) );
  DFF_X1 \reg_mid_1_reg[10]  ( .D(N74), .CK(g_inClk), .Q(reg_mid_1[10]), .QN(
        n1874) );
  DFF_X1 \reg_mid_1_reg[9]  ( .D(N73), .CK(g_inClk), .Q(reg_mid_1[9]), .QN(
        n1844) );
  DFF_X1 \reg_mid_1_reg[8]  ( .D(N72), .CK(g_inClk), .Q(reg_mid_1[8]), .QN(
        n1845) );
  DFF_X1 \reg_mid_1_reg[7]  ( .D(N71), .CK(g_inClk), .Q(reg_mid_1[7]), .QN(
        n1832) );
  DFF_X1 \reg_mid_1_reg[6]  ( .D(N70), .CK(g_inClk), .Q(reg_mid_1[6]), .QN(
        n1846) );
  DFF_X1 \reg_mid_1_reg[5]  ( .D(N69), .CK(g_inClk), .Q(reg_mid_1[5]), .QN(
        n1847) );
  DFF_X1 \reg_mid_1_reg[4]  ( .D(N68), .CK(g_inClk), .Q(reg_mid_1[4]), .QN(
        n1875) );
  DFF_X1 \reg_mid_1_reg[3]  ( .D(N67), .CK(g_inClk), .Q(reg_mid_1[3]), .QN(
        n1853) );
  DFF_X1 \reg_mid_1_reg[2]  ( .D(N66), .CK(g_inClk), .Q(reg_mid_1[2]), .QN(
        n1854) );
  DFF_X1 \reg_mid_1_reg[1]  ( .D(N65), .CK(g_inClk), .Q(reg_mid_1[1]), .QN(
        n1855) );
  DFF_X1 \reg_mid_1_reg[0]  ( .D(N64), .CK(g_inClk), .Q(reg_mid_1[0]), .QN(
        n1876) );
  DFF_X1 \reg_out_reg[126]  ( .D(N254), .CK(g_inClk), .Q(g_outM[126]) );
  DFF_X1 \reg_out_reg[124]  ( .D(N252), .CK(g_inClk), .Q(g_outM[124]) );
  DFF_X1 \reg_out_reg[122]  ( .D(N250), .CK(g_inClk), .Q(g_outM[122]) );
  DFF_X1 \reg_out_reg[120]  ( .D(N248), .CK(g_inClk), .Q(g_outM[120]) );
  DFF_X1 \reg_out_reg[118]  ( .D(N246), .CK(g_inClk), .Q(g_outM[118]) );
  DFF_X1 \reg_out_reg[116]  ( .D(N244), .CK(g_inClk), .Q(g_outM[116]) );
  DFF_X1 \reg_out_reg[115]  ( .D(N243), .CK(g_inClk), .Q(g_outM[115]) );
  DFF_X1 \reg_out_reg[114]  ( .D(N242), .CK(g_inClk), .Q(g_outM[114]) );
  DFF_X1 \reg_out_reg[113]  ( .D(N241), .CK(g_inClk), .Q(g_outM[113]) );
  DFF_X1 \reg_out_reg[112]  ( .D(N240), .CK(g_inClk), .Q(g_outM[112]) );
  DFF_X1 \reg_out_reg[111]  ( .D(N239), .CK(g_inClk), .Q(g_outM[111]) );
  DFF_X1 \reg_out_reg[110]  ( .D(N238), .CK(g_inClk), .Q(g_outM[110]) );
  DFF_X1 \reg_out_reg[109]  ( .D(N237), .CK(g_inClk), .Q(g_outM[109]) );
  DFF_X1 \reg_out_reg[108]  ( .D(N236), .CK(g_inClk), .Q(g_outM[108]) );
  DFF_X1 \reg_out_reg[107]  ( .D(N235), .CK(g_inClk), .Q(g_outM[107]) );
  DFF_X1 \reg_out_reg[106]  ( .D(N234), .CK(g_inClk), .Q(g_outM[106]) );
  DFF_X1 \reg_out_reg[105]  ( .D(N233), .CK(g_inClk), .Q(g_outM[105]) );
  DFF_X1 \reg_out_reg[104]  ( .D(N232), .CK(g_inClk), .Q(g_outM[104]) );
  DFF_X1 \reg_out_reg[103]  ( .D(N231), .CK(g_inClk), .Q(g_outM[103]) );
  DFF_X1 \reg_out_reg[102]  ( .D(N230), .CK(g_inClk), .Q(g_outM[102]) );
  DFF_X1 \reg_out_reg[101]  ( .D(N229), .CK(g_inClk), .Q(g_outM[101]) );
  DFF_X1 \reg_out_reg[100]  ( .D(N228), .CK(g_inClk), .Q(g_outM[100]) );
  DFF_X1 \reg_out_reg[99]  ( .D(N227), .CK(g_inClk), .Q(g_outM[99]) );
  DFF_X1 \reg_out_reg[98]  ( .D(N226), .CK(g_inClk), .Q(g_outM[98]) );
  DFF_X1 \reg_out_reg[97]  ( .D(N225), .CK(g_inClk), .Q(g_outM[97]) );
  DFF_X1 \reg_out_reg[96]  ( .D(N224), .CK(g_inClk), .Q(g_outM[96]) );
  DFF_X1 \reg_out_reg[95]  ( .D(N223), .CK(g_inClk), .Q(g_outM[95]) );
  DFF_X1 \reg_out_reg[94]  ( .D(N222), .CK(g_inClk), .Q(g_outM[94]) );
  DFF_X1 \reg_out_reg[93]  ( .D(N221), .CK(g_inClk), .Q(g_outM[93]) );
  DFF_X1 \reg_out_reg[92]  ( .D(N220), .CK(g_inClk), .Q(g_outM[92]) );
  DFF_X1 \reg_out_reg[91]  ( .D(N219), .CK(g_inClk), .Q(g_outM[91]) );
  DFF_X1 \reg_out_reg[90]  ( .D(N218), .CK(g_inClk), .Q(g_outM[90]) );
  DFF_X1 \reg_out_reg[89]  ( .D(N217), .CK(g_inClk), .Q(g_outM[89]) );
  DFF_X1 \reg_out_reg[88]  ( .D(N216), .CK(g_inClk), .Q(g_outM[88]) );
  DFF_X1 \reg_out_reg[87]  ( .D(N215), .CK(g_inClk), .Q(g_outM[87]) );
  DFF_X1 \reg_out_reg[86]  ( .D(N214), .CK(g_inClk), .Q(g_outM[86]) );
  DFF_X1 \reg_out_reg[85]  ( .D(N213), .CK(g_inClk), .Q(g_outM[85]) );
  DFF_X1 \reg_out_reg[84]  ( .D(N212), .CK(g_inClk), .Q(g_outM[84]) );
  DFF_X1 \reg_out_reg[83]  ( .D(N211), .CK(g_inClk), .Q(g_outM[83]) );
  DFF_X1 \reg_out_reg[82]  ( .D(N210), .CK(g_inClk), .Q(g_outM[82]) );
  DFF_X1 \reg_out_reg[81]  ( .D(N209), .CK(g_inClk), .Q(g_outM[81]) );
  DFF_X1 \reg_out_reg[80]  ( .D(N208), .CK(g_inClk), .Q(g_outM[80]) );
  DFF_X1 \reg_out_reg[79]  ( .D(N207), .CK(g_inClk), .Q(g_outM[79]) );
  DFF_X1 \reg_out_reg[78]  ( .D(N206), .CK(g_inClk), .Q(g_outM[78]) );
  DFF_X1 \reg_out_reg[77]  ( .D(N205), .CK(g_inClk), .Q(g_outM[77]) );
  DFF_X1 \reg_out_reg[76]  ( .D(N204), .CK(g_inClk), .Q(g_outM[76]) );
  DFF_X1 \reg_out_reg[75]  ( .D(N203), .CK(g_inClk), .Q(g_outM[75]) );
  DFF_X1 \reg_out_reg[74]  ( .D(N202), .CK(g_inClk), .Q(g_outM[74]) );
  DFF_X1 \reg_out_reg[73]  ( .D(N201), .CK(g_inClk), .Q(g_outM[73]) );
  DFF_X1 \reg_out_reg[72]  ( .D(N200), .CK(g_inClk), .Q(g_outM[72]) );
  DFF_X1 \reg_out_reg[71]  ( .D(N199), .CK(g_inClk), .Q(g_outM[71]) );
  DFF_X1 \reg_out_reg[70]  ( .D(N198), .CK(g_inClk), .Q(g_outM[70]) );
  DFF_X1 \reg_out_reg[69]  ( .D(N197), .CK(g_inClk), .Q(g_outM[69]) );
  DFF_X1 \reg_out_reg[68]  ( .D(N196), .CK(g_inClk), .Q(g_outM[68]) );
  DFF_X1 \reg_out_reg[67]  ( .D(N195), .CK(g_inClk), .Q(g_outM[67]) );
  DFF_X1 \reg_out_reg[66]  ( .D(N194), .CK(g_inClk), .Q(g_outM[66]) );
  DFF_X1 \reg_out_reg[65]  ( .D(N193), .CK(g_inClk), .Q(g_outM[65]) );
  DFF_X1 \reg_out_reg[64]  ( .D(N192), .CK(g_inClk), .Q(g_outM[64]) );
  DFF_X1 \reg_out_reg[63]  ( .D(N191), .CK(g_inClk), .Q(g_outM[63]) );
  DFF_X1 \reg_out_reg[62]  ( .D(N190), .CK(g_inClk), .Q(g_outM[62]) );
  DFF_X1 \reg_out_reg[61]  ( .D(N189), .CK(g_inClk), .Q(g_outM[61]) );
  DFF_X1 \reg_out_reg[60]  ( .D(N188), .CK(g_inClk), .Q(g_outM[60]) );
  DFF_X1 \reg_out_reg[59]  ( .D(N187), .CK(g_inClk), .Q(g_outM[59]) );
  DFF_X1 \reg_out_reg[58]  ( .D(N186), .CK(g_inClk), .Q(g_outM[58]) );
  DFF_X1 \reg_out_reg[57]  ( .D(N185), .CK(g_inClk), .Q(g_outM[57]) );
  DFF_X1 \reg_out_reg[56]  ( .D(N184), .CK(g_inClk), .Q(g_outM[56]) );
  DFF_X1 \reg_out_reg[55]  ( .D(N183), .CK(g_inClk), .Q(g_outM[55]) );
  DFF_X1 \reg_out_reg[54]  ( .D(N182), .CK(g_inClk), .Q(g_outM[54]) );
  DFF_X1 \reg_out_reg[53]  ( .D(N181), .CK(g_inClk), .Q(g_outM[53]) );
  DFF_X1 \reg_out_reg[52]  ( .D(N180), .CK(g_inClk), .Q(g_outM[52]) );
  DFF_X1 \reg_out_reg[51]  ( .D(N179), .CK(g_inClk), .Q(g_outM[51]) );
  DFF_X1 \reg_out_reg[50]  ( .D(N178), .CK(g_inClk), .Q(g_outM[50]) );
  DFF_X1 \reg_out_reg[49]  ( .D(N177), .CK(g_inClk), .Q(g_outM[49]) );
  DFF_X1 \reg_out_reg[48]  ( .D(N176), .CK(g_inClk), .Q(g_outM[48]) );
  DFF_X1 \reg_out_reg[47]  ( .D(N175), .CK(g_inClk), .Q(g_outM[47]) );
  DFF_X1 \reg_out_reg[46]  ( .D(N174), .CK(g_inClk), .Q(g_outM[46]) );
  DFF_X1 \reg_out_reg[45]  ( .D(N173), .CK(g_inClk), .Q(g_outM[45]) );
  DFF_X1 \reg_out_reg[44]  ( .D(N172), .CK(g_inClk), .Q(g_outM[44]) );
  DFF_X1 \reg_out_reg[43]  ( .D(N171), .CK(g_inClk), .Q(g_outM[43]) );
  DFF_X1 \reg_out_reg[42]  ( .D(N170), .CK(g_inClk), .Q(g_outM[42]) );
  DFF_X1 \reg_out_reg[41]  ( .D(N169), .CK(g_inClk), .Q(g_outM[41]) );
  DFF_X1 \reg_out_reg[40]  ( .D(N168), .CK(g_inClk), .Q(g_outM[40]) );
  DFF_X1 \reg_out_reg[39]  ( .D(N167), .CK(g_inClk), .Q(g_outM[39]) );
  DFF_X1 \reg_out_reg[38]  ( .D(N166), .CK(g_inClk), .Q(g_outM[38]) );
  DFF_X1 \reg_out_reg[37]  ( .D(N165), .CK(g_inClk), .Q(g_outM[37]) );
  DFF_X1 \reg_out_reg[36]  ( .D(N164), .CK(g_inClk), .Q(g_outM[36]) );
  DFF_X1 \reg_out_reg[35]  ( .D(N163), .CK(g_inClk), .Q(g_outM[35]) );
  DFF_X1 \reg_out_reg[34]  ( .D(N162), .CK(g_inClk), .Q(g_outM[34]) );
  DFF_X1 \reg_out_reg[33]  ( .D(N161), .CK(g_inClk), .Q(g_outM[33]) );
  DFF_X1 \reg_out_reg[32]  ( .D(N160), .CK(g_inClk), .Q(g_outM[32]) );
  DFF_X1 \reg_out_reg[31]  ( .D(N159), .CK(g_inClk), .Q(g_outM[31]) );
  DFF_X1 \reg_out_reg[30]  ( .D(N158), .CK(g_inClk), .Q(g_outM[30]) );
  DFF_X1 \reg_out_reg[29]  ( .D(N157), .CK(g_inClk), .Q(g_outM[29]) );
  DFF_X1 \reg_out_reg[28]  ( .D(N156), .CK(g_inClk), .Q(g_outM[28]) );
  DFF_X1 \reg_out_reg[27]  ( .D(N155), .CK(g_inClk), .Q(g_outM[27]) );
  DFF_X1 \reg_out_reg[26]  ( .D(N154), .CK(g_inClk), .Q(g_outM[26]) );
  DFF_X1 \reg_out_reg[25]  ( .D(N153), .CK(g_inClk), .Q(g_outM[25]) );
  DFF_X1 \reg_out_reg[24]  ( .D(N152), .CK(g_inClk), .Q(g_outM[24]) );
  DFF_X1 \reg_out_reg[23]  ( .D(N151), .CK(g_inClk), .Q(g_outM[23]) );
  DFF_X1 \reg_out_reg[22]  ( .D(N150), .CK(g_inClk), .Q(g_outM[22]) );
  DFF_X1 \reg_out_reg[21]  ( .D(N149), .CK(g_inClk), .Q(g_outM[21]) );
  DFF_X1 \reg_out_reg[20]  ( .D(N148), .CK(g_inClk), .Q(g_outM[20]) );
  DFF_X1 \reg_out_reg[19]  ( .D(N147), .CK(g_inClk), .Q(g_outM[19]) );
  DFF_X1 \reg_out_reg[18]  ( .D(N146), .CK(g_inClk), .Q(g_outM[18]) );
  DFF_X1 \reg_out_reg[17]  ( .D(N145), .CK(g_inClk), .Q(g_outM[17]) );
  DFF_X1 \reg_out_reg[16]  ( .D(N144), .CK(g_inClk), .Q(g_outM[16]) );
  DFF_X1 \reg_out_reg[15]  ( .D(N143), .CK(g_inClk), .Q(g_outM[15]) );
  DFF_X1 \reg_out_reg[14]  ( .D(N142), .CK(g_inClk), .Q(g_outM[14]) );
  DFF_X1 \reg_out_reg[13]  ( .D(N141), .CK(g_inClk), .Q(g_outM[13]) );
  DFF_X1 \reg_out_reg[12]  ( .D(N140), .CK(g_inClk), .Q(g_outM[12]) );
  DFF_X1 \reg_out_reg[11]  ( .D(N139), .CK(g_inClk), .Q(g_outM[11]) );
  DFF_X1 \reg_out_reg[10]  ( .D(N138), .CK(g_inClk), .Q(g_outM[10]) );
  DFF_X1 \reg_out_reg[9]  ( .D(N137), .CK(g_inClk), .Q(g_outM[9]) );
  DFF_X1 \reg_out_reg[8]  ( .D(N136), .CK(g_inClk), .Q(g_outM[8]) );
  DFF_X1 \reg_out_reg[7]  ( .D(N135), .CK(g_inClk), .Q(g_outM[7]) );
  DFF_X1 \reg_out_reg[6]  ( .D(N134), .CK(g_inClk), .Q(g_outM[6]) );
  DFF_X1 \reg_out_reg[5]  ( .D(N133), .CK(g_inClk), .Q(g_outM[5]) );
  DFF_X1 \reg_out_reg[4]  ( .D(N132), .CK(g_inClk), .Q(g_outM[4]) );
  DFF_X1 \reg_out_reg[3]  ( .D(N131), .CK(g_inClk), .Q(g_outM[3]) );
  DFF_X1 \reg_out_reg[2]  ( .D(N130), .CK(g_inClk), .Q(g_outM[2]) );
  DFF_X1 \reg_out_reg[1]  ( .D(N129), .CK(g_inClk), .Q(g_outM[1]) );
  DFF_X1 \reg_out_reg[0]  ( .D(N128), .CK(g_inClk), .Q(g_outM[0]) );
  FA_X1 \mult_20/S3_2_30  ( .A(\mult_20/ab[2][30] ), .B(\mult_20/n33 ), .CI(
        \mult_20/ab[1][31] ), .CO(\mult_20/CARRYB[2][30] ), .S(
        \mult_20/SUMB[2][30] ) );
  FA_X1 \mult_20/S2_2_29  ( .A(\mult_20/ab[2][29] ), .B(\mult_20/n3 ), .CI(
        \mult_20/n34 ), .CO(\mult_20/CARRYB[2][29] ), .S(\mult_20/SUMB[2][29] ) );
  FA_X1 \mult_20/S2_2_28  ( .A(\mult_20/ab[2][28] ), .B(\mult_20/n4 ), .CI(
        \mult_20/n35 ), .CO(\mult_20/CARRYB[2][28] ), .S(\mult_20/SUMB[2][28] ) );
  FA_X1 \mult_20/S2_2_27  ( .A(\mult_20/ab[2][27] ), .B(\mult_20/n5 ), .CI(
        \mult_20/n36 ), .CO(\mult_20/CARRYB[2][27] ), .S(\mult_20/SUMB[2][27] ) );
  FA_X1 \mult_20/S2_2_26  ( .A(\mult_20/ab[2][26] ), .B(\mult_20/n6 ), .CI(
        \mult_20/n37 ), .CO(\mult_20/CARRYB[2][26] ), .S(\mult_20/SUMB[2][26] ) );
  FA_X1 \mult_20/S2_2_25  ( .A(\mult_20/ab[2][25] ), .B(\mult_20/n7 ), .CI(
        \mult_20/n38 ), .CO(\mult_20/CARRYB[2][25] ), .S(\mult_20/SUMB[2][25] ) );
  FA_X1 \mult_20/S2_2_24  ( .A(\mult_20/ab[2][24] ), .B(\mult_20/n8 ), .CI(
        \mult_20/n39 ), .CO(\mult_20/CARRYB[2][24] ), .S(\mult_20/SUMB[2][24] ) );
  FA_X1 \mult_20/S2_2_23  ( .A(\mult_20/ab[2][23] ), .B(\mult_20/n9 ), .CI(
        \mult_20/n40 ), .CO(\mult_20/CARRYB[2][23] ), .S(\mult_20/SUMB[2][23] ) );
  FA_X1 \mult_20/S2_2_22  ( .A(\mult_20/ab[2][22] ), .B(\mult_20/n10 ), .CI(
        \mult_20/n41 ), .CO(\mult_20/CARRYB[2][22] ), .S(\mult_20/SUMB[2][22] ) );
  FA_X1 \mult_20/S2_2_21  ( .A(\mult_20/ab[2][21] ), .B(\mult_20/n11 ), .CI(
        \mult_20/n42 ), .CO(\mult_20/CARRYB[2][21] ), .S(\mult_20/SUMB[2][21] ) );
  FA_X1 \mult_20/S2_2_20  ( .A(\mult_20/ab[2][20] ), .B(\mult_20/n12 ), .CI(
        \mult_20/n43 ), .CO(\mult_20/CARRYB[2][20] ), .S(\mult_20/SUMB[2][20] ) );
  FA_X1 \mult_20/S2_2_19  ( .A(\mult_20/ab[2][19] ), .B(\mult_20/n13 ), .CI(
        \mult_20/n44 ), .CO(\mult_20/CARRYB[2][19] ), .S(\mult_20/SUMB[2][19] ) );
  FA_X1 \mult_20/S2_2_18  ( .A(\mult_20/ab[2][18] ), .B(\mult_20/n14 ), .CI(
        \mult_20/n45 ), .CO(\mult_20/CARRYB[2][18] ), .S(\mult_20/SUMB[2][18] ) );
  FA_X1 \mult_20/S2_2_17  ( .A(\mult_20/ab[2][17] ), .B(\mult_20/n15 ), .CI(
        \mult_20/n46 ), .CO(\mult_20/CARRYB[2][17] ), .S(\mult_20/SUMB[2][17] ) );
  FA_X1 \mult_20/S2_2_16  ( .A(\mult_20/ab[2][16] ), .B(\mult_20/n16 ), .CI(
        \mult_20/n47 ), .CO(\mult_20/CARRYB[2][16] ), .S(\mult_20/SUMB[2][16] ) );
  FA_X1 \mult_20/S2_2_15  ( .A(\mult_20/ab[2][15] ), .B(\mult_20/n17 ), .CI(
        \mult_20/n48 ), .CO(\mult_20/CARRYB[2][15] ), .S(\mult_20/SUMB[2][15] ) );
  FA_X1 \mult_20/S2_2_14  ( .A(\mult_20/ab[2][14] ), .B(\mult_20/n18 ), .CI(
        \mult_20/n49 ), .CO(\mult_20/CARRYB[2][14] ), .S(\mult_20/SUMB[2][14] ) );
  FA_X1 \mult_20/S2_2_13  ( .A(\mult_20/ab[2][13] ), .B(\mult_20/n19 ), .CI(
        \mult_20/n50 ), .CO(\mult_20/CARRYB[2][13] ), .S(\mult_20/SUMB[2][13] ) );
  FA_X1 \mult_20/S2_2_12  ( .A(\mult_20/ab[2][12] ), .B(\mult_20/n20 ), .CI(
        \mult_20/n51 ), .CO(\mult_20/CARRYB[2][12] ), .S(\mult_20/SUMB[2][12] ) );
  FA_X1 \mult_20/S2_2_11  ( .A(\mult_20/ab[2][11] ), .B(\mult_20/n21 ), .CI(
        \mult_20/n52 ), .CO(\mult_20/CARRYB[2][11] ), .S(\mult_20/SUMB[2][11] ) );
  FA_X1 \mult_20/S2_2_10  ( .A(\mult_20/ab[2][10] ), .B(\mult_20/n22 ), .CI(
        \mult_20/n53 ), .CO(\mult_20/CARRYB[2][10] ), .S(\mult_20/SUMB[2][10] ) );
  FA_X1 \mult_20/S2_2_9  ( .A(\mult_20/ab[2][9] ), .B(\mult_20/n23 ), .CI(
        \mult_20/n54 ), .CO(\mult_20/CARRYB[2][9] ), .S(\mult_20/SUMB[2][9] )
         );
  FA_X1 \mult_20/S2_2_8  ( .A(\mult_20/ab[2][8] ), .B(\mult_20/n24 ), .CI(
        \mult_20/n55 ), .CO(\mult_20/CARRYB[2][8] ), .S(\mult_20/SUMB[2][8] )
         );
  FA_X1 \mult_20/S2_2_7  ( .A(\mult_20/ab[2][7] ), .B(\mult_20/n25 ), .CI(
        \mult_20/n56 ), .CO(\mult_20/CARRYB[2][7] ), .S(\mult_20/SUMB[2][7] )
         );
  FA_X1 \mult_20/S2_2_6  ( .A(\mult_20/ab[2][6] ), .B(\mult_20/n26 ), .CI(
        \mult_20/n57 ), .CO(\mult_20/CARRYB[2][6] ), .S(\mult_20/SUMB[2][6] )
         );
  FA_X1 \mult_20/S2_2_5  ( .A(\mult_20/ab[2][5] ), .B(\mult_20/n27 ), .CI(
        \mult_20/n58 ), .CO(\mult_20/CARRYB[2][5] ), .S(\mult_20/SUMB[2][5] )
         );
  FA_X1 \mult_20/S2_2_4  ( .A(\mult_20/ab[2][4] ), .B(\mult_20/n28 ), .CI(
        \mult_20/n59 ), .CO(\mult_20/CARRYB[2][4] ), .S(\mult_20/SUMB[2][4] )
         );
  FA_X1 \mult_20/S2_2_3  ( .A(\mult_20/ab[2][3] ), .B(\mult_20/n29 ), .CI(
        \mult_20/n60 ), .CO(\mult_20/CARRYB[2][3] ), .S(\mult_20/SUMB[2][3] )
         );
  FA_X1 \mult_20/S2_2_2  ( .A(\mult_20/ab[2][2] ), .B(\mult_20/n30 ), .CI(
        \mult_20/n61 ), .CO(\mult_20/CARRYB[2][2] ), .S(\mult_20/SUMB[2][2] )
         );
  FA_X1 \mult_20/S2_2_1  ( .A(\mult_20/ab[2][1] ), .B(\mult_20/n31 ), .CI(
        \mult_20/n62 ), .CO(\mult_20/CARRYB[2][1] ), .S(\mult_20/SUMB[2][1] )
         );
  FA_X1 \mult_20/S1_2_0  ( .A(\mult_20/ab[2][0] ), .B(\mult_20/n32 ), .CI(
        \mult_20/n63 ), .CO(\mult_20/CARRYB[2][0] ), .S(N66) );
  FA_X1 \mult_20/S3_3_30  ( .A(\mult_20/ab[3][30] ), .B(
        \mult_20/CARRYB[2][30] ), .CI(\mult_20/ab[2][31] ), .CO(
        \mult_20/CARRYB[3][30] ), .S(\mult_20/SUMB[3][30] ) );
  FA_X1 \mult_20/S2_3_29  ( .A(\mult_20/ab[3][29] ), .B(
        \mult_20/CARRYB[2][29] ), .CI(\mult_20/SUMB[2][30] ), .CO(
        \mult_20/CARRYB[3][29] ), .S(\mult_20/SUMB[3][29] ) );
  FA_X1 \mult_20/S2_3_28  ( .A(\mult_20/ab[3][28] ), .B(
        \mult_20/CARRYB[2][28] ), .CI(\mult_20/SUMB[2][29] ), .CO(
        \mult_20/CARRYB[3][28] ), .S(\mult_20/SUMB[3][28] ) );
  FA_X1 \mult_20/S2_3_27  ( .A(\mult_20/ab[3][27] ), .B(
        \mult_20/CARRYB[2][27] ), .CI(\mult_20/SUMB[2][28] ), .CO(
        \mult_20/CARRYB[3][27] ), .S(\mult_20/SUMB[3][27] ) );
  FA_X1 \mult_20/S2_3_26  ( .A(\mult_20/ab[3][26] ), .B(
        \mult_20/CARRYB[2][26] ), .CI(\mult_20/SUMB[2][27] ), .CO(
        \mult_20/CARRYB[3][26] ), .S(\mult_20/SUMB[3][26] ) );
  FA_X1 \mult_20/S2_3_25  ( .A(\mult_20/ab[3][25] ), .B(
        \mult_20/CARRYB[2][25] ), .CI(\mult_20/SUMB[2][26] ), .CO(
        \mult_20/CARRYB[3][25] ), .S(\mult_20/SUMB[3][25] ) );
  FA_X1 \mult_20/S2_3_24  ( .A(\mult_20/ab[3][24] ), .B(
        \mult_20/CARRYB[2][24] ), .CI(\mult_20/SUMB[2][25] ), .CO(
        \mult_20/CARRYB[3][24] ), .S(\mult_20/SUMB[3][24] ) );
  FA_X1 \mult_20/S2_3_23  ( .A(\mult_20/ab[3][23] ), .B(
        \mult_20/CARRYB[2][23] ), .CI(\mult_20/SUMB[2][24] ), .CO(
        \mult_20/CARRYB[3][23] ), .S(\mult_20/SUMB[3][23] ) );
  FA_X1 \mult_20/S2_3_22  ( .A(\mult_20/ab[3][22] ), .B(
        \mult_20/CARRYB[2][22] ), .CI(\mult_20/SUMB[2][23] ), .CO(
        \mult_20/CARRYB[3][22] ), .S(\mult_20/SUMB[3][22] ) );
  FA_X1 \mult_20/S2_3_21  ( .A(\mult_20/ab[3][21] ), .B(
        \mult_20/CARRYB[2][21] ), .CI(\mult_20/SUMB[2][22] ), .CO(
        \mult_20/CARRYB[3][21] ), .S(\mult_20/SUMB[3][21] ) );
  FA_X1 \mult_20/S2_3_20  ( .A(\mult_20/ab[3][20] ), .B(
        \mult_20/CARRYB[2][20] ), .CI(\mult_20/SUMB[2][21] ), .CO(
        \mult_20/CARRYB[3][20] ), .S(\mult_20/SUMB[3][20] ) );
  FA_X1 \mult_20/S2_3_19  ( .A(\mult_20/ab[3][19] ), .B(
        \mult_20/CARRYB[2][19] ), .CI(\mult_20/SUMB[2][20] ), .CO(
        \mult_20/CARRYB[3][19] ), .S(\mult_20/SUMB[3][19] ) );
  FA_X1 \mult_20/S2_3_18  ( .A(\mult_20/ab[3][18] ), .B(
        \mult_20/CARRYB[2][18] ), .CI(\mult_20/SUMB[2][19] ), .CO(
        \mult_20/CARRYB[3][18] ), .S(\mult_20/SUMB[3][18] ) );
  FA_X1 \mult_20/S2_3_17  ( .A(\mult_20/ab[3][17] ), .B(
        \mult_20/CARRYB[2][17] ), .CI(\mult_20/SUMB[2][18] ), .CO(
        \mult_20/CARRYB[3][17] ), .S(\mult_20/SUMB[3][17] ) );
  FA_X1 \mult_20/S2_3_16  ( .A(\mult_20/ab[3][16] ), .B(
        \mult_20/CARRYB[2][16] ), .CI(\mult_20/SUMB[2][17] ), .CO(
        \mult_20/CARRYB[3][16] ), .S(\mult_20/SUMB[3][16] ) );
  FA_X1 \mult_20/S2_3_15  ( .A(\mult_20/ab[3][15] ), .B(
        \mult_20/CARRYB[2][15] ), .CI(\mult_20/SUMB[2][16] ), .CO(
        \mult_20/CARRYB[3][15] ), .S(\mult_20/SUMB[3][15] ) );
  FA_X1 \mult_20/S2_3_14  ( .A(\mult_20/ab[3][14] ), .B(
        \mult_20/CARRYB[2][14] ), .CI(\mult_20/SUMB[2][15] ), .CO(
        \mult_20/CARRYB[3][14] ), .S(\mult_20/SUMB[3][14] ) );
  FA_X1 \mult_20/S2_3_13  ( .A(\mult_20/ab[3][13] ), .B(
        \mult_20/CARRYB[2][13] ), .CI(\mult_20/SUMB[2][14] ), .CO(
        \mult_20/CARRYB[3][13] ), .S(\mult_20/SUMB[3][13] ) );
  FA_X1 \mult_20/S2_3_12  ( .A(\mult_20/ab[3][12] ), .B(
        \mult_20/CARRYB[2][12] ), .CI(\mult_20/SUMB[2][13] ), .CO(
        \mult_20/CARRYB[3][12] ), .S(\mult_20/SUMB[3][12] ) );
  FA_X1 \mult_20/S2_3_11  ( .A(\mult_20/ab[3][11] ), .B(
        \mult_20/CARRYB[2][11] ), .CI(\mult_20/SUMB[2][12] ), .CO(
        \mult_20/CARRYB[3][11] ), .S(\mult_20/SUMB[3][11] ) );
  FA_X1 \mult_20/S2_3_10  ( .A(\mult_20/ab[3][10] ), .B(
        \mult_20/CARRYB[2][10] ), .CI(\mult_20/SUMB[2][11] ), .CO(
        \mult_20/CARRYB[3][10] ), .S(\mult_20/SUMB[3][10] ) );
  FA_X1 \mult_20/S2_3_9  ( .A(\mult_20/ab[3][9] ), .B(\mult_20/CARRYB[2][9] ), 
        .CI(\mult_20/SUMB[2][10] ), .CO(\mult_20/CARRYB[3][9] ), .S(
        \mult_20/SUMB[3][9] ) );
  FA_X1 \mult_20/S2_3_8  ( .A(\mult_20/ab[3][8] ), .B(\mult_20/CARRYB[2][8] ), 
        .CI(\mult_20/SUMB[2][9] ), .CO(\mult_20/CARRYB[3][8] ), .S(
        \mult_20/SUMB[3][8] ) );
  FA_X1 \mult_20/S2_3_7  ( .A(\mult_20/ab[3][7] ), .B(\mult_20/CARRYB[2][7] ), 
        .CI(\mult_20/SUMB[2][8] ), .CO(\mult_20/CARRYB[3][7] ), .S(
        \mult_20/SUMB[3][7] ) );
  FA_X1 \mult_20/S2_3_6  ( .A(\mult_20/ab[3][6] ), .B(\mult_20/CARRYB[2][6] ), 
        .CI(\mult_20/SUMB[2][7] ), .CO(\mult_20/CARRYB[3][6] ), .S(
        \mult_20/SUMB[3][6] ) );
  FA_X1 \mult_20/S2_3_5  ( .A(\mult_20/ab[3][5] ), .B(\mult_20/CARRYB[2][5] ), 
        .CI(\mult_20/SUMB[2][6] ), .CO(\mult_20/CARRYB[3][5] ), .S(
        \mult_20/SUMB[3][5] ) );
  FA_X1 \mult_20/S2_3_4  ( .A(\mult_20/ab[3][4] ), .B(\mult_20/CARRYB[2][4] ), 
        .CI(\mult_20/SUMB[2][5] ), .CO(\mult_20/CARRYB[3][4] ), .S(
        \mult_20/SUMB[3][4] ) );
  FA_X1 \mult_20/S2_3_3  ( .A(\mult_20/ab[3][3] ), .B(\mult_20/CARRYB[2][3] ), 
        .CI(\mult_20/SUMB[2][4] ), .CO(\mult_20/CARRYB[3][3] ), .S(
        \mult_20/SUMB[3][3] ) );
  FA_X1 \mult_20/S2_3_2  ( .A(\mult_20/ab[3][2] ), .B(\mult_20/CARRYB[2][2] ), 
        .CI(\mult_20/SUMB[2][3] ), .CO(\mult_20/CARRYB[3][2] ), .S(
        \mult_20/SUMB[3][2] ) );
  FA_X1 \mult_20/S2_3_1  ( .A(\mult_20/ab[3][1] ), .B(\mult_20/CARRYB[2][1] ), 
        .CI(\mult_20/SUMB[2][2] ), .CO(\mult_20/CARRYB[3][1] ), .S(
        \mult_20/SUMB[3][1] ) );
  FA_X1 \mult_20/S1_3_0  ( .A(\mult_20/ab[3][0] ), .B(\mult_20/CARRYB[2][0] ), 
        .CI(\mult_20/SUMB[2][1] ), .CO(\mult_20/CARRYB[3][0] ), .S(N67) );
  FA_X1 \mult_20/S3_4_30  ( .A(\mult_20/ab[4][30] ), .B(
        \mult_20/CARRYB[3][30] ), .CI(\mult_20/ab[3][31] ), .CO(
        \mult_20/CARRYB[4][30] ), .S(\mult_20/SUMB[4][30] ) );
  FA_X1 \mult_20/S2_4_29  ( .A(\mult_20/ab[4][29] ), .B(
        \mult_20/CARRYB[3][29] ), .CI(\mult_20/SUMB[3][30] ), .CO(
        \mult_20/CARRYB[4][29] ), .S(\mult_20/SUMB[4][29] ) );
  FA_X1 \mult_20/S2_4_28  ( .A(\mult_20/ab[4][28] ), .B(
        \mult_20/CARRYB[3][28] ), .CI(\mult_20/SUMB[3][29] ), .CO(
        \mult_20/CARRYB[4][28] ), .S(\mult_20/SUMB[4][28] ) );
  FA_X1 \mult_20/S2_4_27  ( .A(\mult_20/ab[4][27] ), .B(
        \mult_20/CARRYB[3][27] ), .CI(\mult_20/SUMB[3][28] ), .CO(
        \mult_20/CARRYB[4][27] ), .S(\mult_20/SUMB[4][27] ) );
  FA_X1 \mult_20/S2_4_26  ( .A(\mult_20/ab[4][26] ), .B(
        \mult_20/CARRYB[3][26] ), .CI(\mult_20/SUMB[3][27] ), .CO(
        \mult_20/CARRYB[4][26] ), .S(\mult_20/SUMB[4][26] ) );
  FA_X1 \mult_20/S2_4_25  ( .A(\mult_20/ab[4][25] ), .B(
        \mult_20/CARRYB[3][25] ), .CI(\mult_20/SUMB[3][26] ), .CO(
        \mult_20/CARRYB[4][25] ), .S(\mult_20/SUMB[4][25] ) );
  FA_X1 \mult_20/S2_4_24  ( .A(\mult_20/ab[4][24] ), .B(
        \mult_20/CARRYB[3][24] ), .CI(\mult_20/SUMB[3][25] ), .CO(
        \mult_20/CARRYB[4][24] ), .S(\mult_20/SUMB[4][24] ) );
  FA_X1 \mult_20/S2_4_23  ( .A(\mult_20/ab[4][23] ), .B(
        \mult_20/CARRYB[3][23] ), .CI(\mult_20/SUMB[3][24] ), .CO(
        \mult_20/CARRYB[4][23] ), .S(\mult_20/SUMB[4][23] ) );
  FA_X1 \mult_20/S2_4_22  ( .A(\mult_20/ab[4][22] ), .B(
        \mult_20/CARRYB[3][22] ), .CI(\mult_20/SUMB[3][23] ), .CO(
        \mult_20/CARRYB[4][22] ), .S(\mult_20/SUMB[4][22] ) );
  FA_X1 \mult_20/S2_4_21  ( .A(\mult_20/ab[4][21] ), .B(
        \mult_20/CARRYB[3][21] ), .CI(\mult_20/SUMB[3][22] ), .CO(
        \mult_20/CARRYB[4][21] ), .S(\mult_20/SUMB[4][21] ) );
  FA_X1 \mult_20/S2_4_20  ( .A(\mult_20/ab[4][20] ), .B(
        \mult_20/CARRYB[3][20] ), .CI(\mult_20/SUMB[3][21] ), .CO(
        \mult_20/CARRYB[4][20] ), .S(\mult_20/SUMB[4][20] ) );
  FA_X1 \mult_20/S2_4_19  ( .A(\mult_20/ab[4][19] ), .B(
        \mult_20/CARRYB[3][19] ), .CI(\mult_20/SUMB[3][20] ), .CO(
        \mult_20/CARRYB[4][19] ), .S(\mult_20/SUMB[4][19] ) );
  FA_X1 \mult_20/S2_4_18  ( .A(\mult_20/ab[4][18] ), .B(
        \mult_20/CARRYB[3][18] ), .CI(\mult_20/SUMB[3][19] ), .CO(
        \mult_20/CARRYB[4][18] ), .S(\mult_20/SUMB[4][18] ) );
  FA_X1 \mult_20/S2_4_17  ( .A(\mult_20/ab[4][17] ), .B(
        \mult_20/CARRYB[3][17] ), .CI(\mult_20/SUMB[3][18] ), .CO(
        \mult_20/CARRYB[4][17] ), .S(\mult_20/SUMB[4][17] ) );
  FA_X1 \mult_20/S2_4_16  ( .A(\mult_20/ab[4][16] ), .B(
        \mult_20/CARRYB[3][16] ), .CI(\mult_20/SUMB[3][17] ), .CO(
        \mult_20/CARRYB[4][16] ), .S(\mult_20/SUMB[4][16] ) );
  FA_X1 \mult_20/S2_4_15  ( .A(\mult_20/ab[4][15] ), .B(
        \mult_20/CARRYB[3][15] ), .CI(\mult_20/SUMB[3][16] ), .CO(
        \mult_20/CARRYB[4][15] ), .S(\mult_20/SUMB[4][15] ) );
  FA_X1 \mult_20/S2_4_14  ( .A(\mult_20/ab[4][14] ), .B(
        \mult_20/CARRYB[3][14] ), .CI(\mult_20/SUMB[3][15] ), .CO(
        \mult_20/CARRYB[4][14] ), .S(\mult_20/SUMB[4][14] ) );
  FA_X1 \mult_20/S2_4_13  ( .A(\mult_20/ab[4][13] ), .B(
        \mult_20/CARRYB[3][13] ), .CI(\mult_20/SUMB[3][14] ), .CO(
        \mult_20/CARRYB[4][13] ), .S(\mult_20/SUMB[4][13] ) );
  FA_X1 \mult_20/S2_4_12  ( .A(\mult_20/ab[4][12] ), .B(
        \mult_20/CARRYB[3][12] ), .CI(\mult_20/SUMB[3][13] ), .CO(
        \mult_20/CARRYB[4][12] ), .S(\mult_20/SUMB[4][12] ) );
  FA_X1 \mult_20/S2_4_11  ( .A(\mult_20/ab[4][11] ), .B(
        \mult_20/CARRYB[3][11] ), .CI(\mult_20/SUMB[3][12] ), .CO(
        \mult_20/CARRYB[4][11] ), .S(\mult_20/SUMB[4][11] ) );
  FA_X1 \mult_20/S2_4_10  ( .A(\mult_20/ab[4][10] ), .B(
        \mult_20/CARRYB[3][10] ), .CI(\mult_20/SUMB[3][11] ), .CO(
        \mult_20/CARRYB[4][10] ), .S(\mult_20/SUMB[4][10] ) );
  FA_X1 \mult_20/S2_4_9  ( .A(\mult_20/ab[4][9] ), .B(\mult_20/CARRYB[3][9] ), 
        .CI(\mult_20/SUMB[3][10] ), .CO(\mult_20/CARRYB[4][9] ), .S(
        \mult_20/SUMB[4][9] ) );
  FA_X1 \mult_20/S2_4_8  ( .A(\mult_20/ab[4][8] ), .B(\mult_20/CARRYB[3][8] ), 
        .CI(\mult_20/SUMB[3][9] ), .CO(\mult_20/CARRYB[4][8] ), .S(
        \mult_20/SUMB[4][8] ) );
  FA_X1 \mult_20/S2_4_7  ( .A(\mult_20/ab[4][7] ), .B(\mult_20/CARRYB[3][7] ), 
        .CI(\mult_20/SUMB[3][8] ), .CO(\mult_20/CARRYB[4][7] ), .S(
        \mult_20/SUMB[4][7] ) );
  FA_X1 \mult_20/S2_4_6  ( .A(\mult_20/ab[4][6] ), .B(\mult_20/CARRYB[3][6] ), 
        .CI(\mult_20/SUMB[3][7] ), .CO(\mult_20/CARRYB[4][6] ), .S(
        \mult_20/SUMB[4][6] ) );
  FA_X1 \mult_20/S2_4_5  ( .A(\mult_20/ab[4][5] ), .B(\mult_20/CARRYB[3][5] ), 
        .CI(\mult_20/SUMB[3][6] ), .CO(\mult_20/CARRYB[4][5] ), .S(
        \mult_20/SUMB[4][5] ) );
  FA_X1 \mult_20/S2_4_4  ( .A(\mult_20/ab[4][4] ), .B(\mult_20/CARRYB[3][4] ), 
        .CI(\mult_20/SUMB[3][5] ), .CO(\mult_20/CARRYB[4][4] ), .S(
        \mult_20/SUMB[4][4] ) );
  FA_X1 \mult_20/S2_4_3  ( .A(\mult_20/ab[4][3] ), .B(\mult_20/CARRYB[3][3] ), 
        .CI(\mult_20/SUMB[3][4] ), .CO(\mult_20/CARRYB[4][3] ), .S(
        \mult_20/SUMB[4][3] ) );
  FA_X1 \mult_20/S2_4_2  ( .A(\mult_20/ab[4][2] ), .B(\mult_20/CARRYB[3][2] ), 
        .CI(\mult_20/SUMB[3][3] ), .CO(\mult_20/CARRYB[4][2] ), .S(
        \mult_20/SUMB[4][2] ) );
  FA_X1 \mult_20/S2_4_1  ( .A(\mult_20/ab[4][1] ), .B(\mult_20/CARRYB[3][1] ), 
        .CI(\mult_20/SUMB[3][2] ), .CO(\mult_20/CARRYB[4][1] ), .S(
        \mult_20/SUMB[4][1] ) );
  FA_X1 \mult_20/S1_4_0  ( .A(\mult_20/ab[4][0] ), .B(\mult_20/CARRYB[3][0] ), 
        .CI(\mult_20/SUMB[3][1] ), .CO(\mult_20/CARRYB[4][0] ), .S(N68) );
  FA_X1 \mult_20/S3_5_30  ( .A(\mult_20/ab[5][30] ), .B(
        \mult_20/CARRYB[4][30] ), .CI(\mult_20/ab[4][31] ), .CO(
        \mult_20/CARRYB[5][30] ), .S(\mult_20/SUMB[5][30] ) );
  FA_X1 \mult_20/S2_5_29  ( .A(\mult_20/ab[5][29] ), .B(
        \mult_20/CARRYB[4][29] ), .CI(\mult_20/SUMB[4][30] ), .CO(
        \mult_20/CARRYB[5][29] ), .S(\mult_20/SUMB[5][29] ) );
  FA_X1 \mult_20/S2_5_28  ( .A(\mult_20/ab[5][28] ), .B(
        \mult_20/CARRYB[4][28] ), .CI(\mult_20/SUMB[4][29] ), .CO(
        \mult_20/CARRYB[5][28] ), .S(\mult_20/SUMB[5][28] ) );
  FA_X1 \mult_20/S2_5_27  ( .A(\mult_20/ab[5][27] ), .B(
        \mult_20/CARRYB[4][27] ), .CI(\mult_20/SUMB[4][28] ), .CO(
        \mult_20/CARRYB[5][27] ), .S(\mult_20/SUMB[5][27] ) );
  FA_X1 \mult_20/S2_5_26  ( .A(\mult_20/ab[5][26] ), .B(
        \mult_20/CARRYB[4][26] ), .CI(\mult_20/SUMB[4][27] ), .CO(
        \mult_20/CARRYB[5][26] ), .S(\mult_20/SUMB[5][26] ) );
  FA_X1 \mult_20/S2_5_25  ( .A(\mult_20/ab[5][25] ), .B(
        \mult_20/CARRYB[4][25] ), .CI(\mult_20/SUMB[4][26] ), .CO(
        \mult_20/CARRYB[5][25] ), .S(\mult_20/SUMB[5][25] ) );
  FA_X1 \mult_20/S2_5_24  ( .A(\mult_20/ab[5][24] ), .B(
        \mult_20/CARRYB[4][24] ), .CI(\mult_20/SUMB[4][25] ), .CO(
        \mult_20/CARRYB[5][24] ), .S(\mult_20/SUMB[5][24] ) );
  FA_X1 \mult_20/S2_5_23  ( .A(\mult_20/ab[5][23] ), .B(
        \mult_20/CARRYB[4][23] ), .CI(\mult_20/SUMB[4][24] ), .CO(
        \mult_20/CARRYB[5][23] ), .S(\mult_20/SUMB[5][23] ) );
  FA_X1 \mult_20/S2_5_22  ( .A(\mult_20/ab[5][22] ), .B(
        \mult_20/CARRYB[4][22] ), .CI(\mult_20/SUMB[4][23] ), .CO(
        \mult_20/CARRYB[5][22] ), .S(\mult_20/SUMB[5][22] ) );
  FA_X1 \mult_20/S2_5_21  ( .A(\mult_20/ab[5][21] ), .B(
        \mult_20/CARRYB[4][21] ), .CI(\mult_20/SUMB[4][22] ), .CO(
        \mult_20/CARRYB[5][21] ), .S(\mult_20/SUMB[5][21] ) );
  FA_X1 \mult_20/S2_5_20  ( .A(\mult_20/ab[5][20] ), .B(
        \mult_20/CARRYB[4][20] ), .CI(\mult_20/SUMB[4][21] ), .CO(
        \mult_20/CARRYB[5][20] ), .S(\mult_20/SUMB[5][20] ) );
  FA_X1 \mult_20/S2_5_19  ( .A(\mult_20/ab[5][19] ), .B(
        \mult_20/CARRYB[4][19] ), .CI(\mult_20/SUMB[4][20] ), .CO(
        \mult_20/CARRYB[5][19] ), .S(\mult_20/SUMB[5][19] ) );
  FA_X1 \mult_20/S2_5_18  ( .A(\mult_20/ab[5][18] ), .B(
        \mult_20/CARRYB[4][18] ), .CI(\mult_20/SUMB[4][19] ), .CO(
        \mult_20/CARRYB[5][18] ), .S(\mult_20/SUMB[5][18] ) );
  FA_X1 \mult_20/S2_5_17  ( .A(\mult_20/ab[5][17] ), .B(
        \mult_20/CARRYB[4][17] ), .CI(\mult_20/SUMB[4][18] ), .CO(
        \mult_20/CARRYB[5][17] ), .S(\mult_20/SUMB[5][17] ) );
  FA_X1 \mult_20/S2_5_16  ( .A(\mult_20/ab[5][16] ), .B(
        \mult_20/CARRYB[4][16] ), .CI(\mult_20/SUMB[4][17] ), .CO(
        \mult_20/CARRYB[5][16] ), .S(\mult_20/SUMB[5][16] ) );
  FA_X1 \mult_20/S2_5_15  ( .A(\mult_20/ab[5][15] ), .B(
        \mult_20/CARRYB[4][15] ), .CI(\mult_20/SUMB[4][16] ), .CO(
        \mult_20/CARRYB[5][15] ), .S(\mult_20/SUMB[5][15] ) );
  FA_X1 \mult_20/S2_5_14  ( .A(\mult_20/ab[5][14] ), .B(
        \mult_20/CARRYB[4][14] ), .CI(\mult_20/SUMB[4][15] ), .CO(
        \mult_20/CARRYB[5][14] ), .S(\mult_20/SUMB[5][14] ) );
  FA_X1 \mult_20/S2_5_13  ( .A(\mult_20/ab[5][13] ), .B(
        \mult_20/CARRYB[4][13] ), .CI(\mult_20/SUMB[4][14] ), .CO(
        \mult_20/CARRYB[5][13] ), .S(\mult_20/SUMB[5][13] ) );
  FA_X1 \mult_20/S2_5_12  ( .A(\mult_20/ab[5][12] ), .B(
        \mult_20/CARRYB[4][12] ), .CI(\mult_20/SUMB[4][13] ), .CO(
        \mult_20/CARRYB[5][12] ), .S(\mult_20/SUMB[5][12] ) );
  FA_X1 \mult_20/S2_5_11  ( .A(\mult_20/ab[5][11] ), .B(
        \mult_20/CARRYB[4][11] ), .CI(\mult_20/SUMB[4][12] ), .CO(
        \mult_20/CARRYB[5][11] ), .S(\mult_20/SUMB[5][11] ) );
  FA_X1 \mult_20/S2_5_10  ( .A(\mult_20/ab[5][10] ), .B(
        \mult_20/CARRYB[4][10] ), .CI(\mult_20/SUMB[4][11] ), .CO(
        \mult_20/CARRYB[5][10] ), .S(\mult_20/SUMB[5][10] ) );
  FA_X1 \mult_20/S2_5_9  ( .A(\mult_20/ab[5][9] ), .B(\mult_20/CARRYB[4][9] ), 
        .CI(\mult_20/SUMB[4][10] ), .CO(\mult_20/CARRYB[5][9] ), .S(
        \mult_20/SUMB[5][9] ) );
  FA_X1 \mult_20/S2_5_8  ( .A(\mult_20/ab[5][8] ), .B(\mult_20/CARRYB[4][8] ), 
        .CI(\mult_20/SUMB[4][9] ), .CO(\mult_20/CARRYB[5][8] ), .S(
        \mult_20/SUMB[5][8] ) );
  FA_X1 \mult_20/S2_5_7  ( .A(\mult_20/ab[5][7] ), .B(\mult_20/CARRYB[4][7] ), 
        .CI(\mult_20/SUMB[4][8] ), .CO(\mult_20/CARRYB[5][7] ), .S(
        \mult_20/SUMB[5][7] ) );
  FA_X1 \mult_20/S2_5_6  ( .A(\mult_20/ab[5][6] ), .B(\mult_20/CARRYB[4][6] ), 
        .CI(\mult_20/SUMB[4][7] ), .CO(\mult_20/CARRYB[5][6] ), .S(
        \mult_20/SUMB[5][6] ) );
  FA_X1 \mult_20/S2_5_5  ( .A(\mult_20/ab[5][5] ), .B(\mult_20/CARRYB[4][5] ), 
        .CI(\mult_20/SUMB[4][6] ), .CO(\mult_20/CARRYB[5][5] ), .S(
        \mult_20/SUMB[5][5] ) );
  FA_X1 \mult_20/S2_5_4  ( .A(\mult_20/ab[5][4] ), .B(\mult_20/CARRYB[4][4] ), 
        .CI(\mult_20/SUMB[4][5] ), .CO(\mult_20/CARRYB[5][4] ), .S(
        \mult_20/SUMB[5][4] ) );
  FA_X1 \mult_20/S2_5_3  ( .A(\mult_20/ab[5][3] ), .B(\mult_20/CARRYB[4][3] ), 
        .CI(\mult_20/SUMB[4][4] ), .CO(\mult_20/CARRYB[5][3] ), .S(
        \mult_20/SUMB[5][3] ) );
  FA_X1 \mult_20/S2_5_2  ( .A(\mult_20/ab[5][2] ), .B(\mult_20/CARRYB[4][2] ), 
        .CI(\mult_20/SUMB[4][3] ), .CO(\mult_20/CARRYB[5][2] ), .S(
        \mult_20/SUMB[5][2] ) );
  FA_X1 \mult_20/S2_5_1  ( .A(\mult_20/ab[5][1] ), .B(\mult_20/CARRYB[4][1] ), 
        .CI(\mult_20/SUMB[4][2] ), .CO(\mult_20/CARRYB[5][1] ), .S(
        \mult_20/SUMB[5][1] ) );
  FA_X1 \mult_20/S1_5_0  ( .A(\mult_20/ab[5][0] ), .B(\mult_20/CARRYB[4][0] ), 
        .CI(\mult_20/SUMB[4][1] ), .CO(\mult_20/CARRYB[5][0] ), .S(N69) );
  FA_X1 \mult_20/S3_6_30  ( .A(\mult_20/ab[6][30] ), .B(
        \mult_20/CARRYB[5][30] ), .CI(\mult_20/ab[5][31] ), .CO(
        \mult_20/CARRYB[6][30] ), .S(\mult_20/SUMB[6][30] ) );
  FA_X1 \mult_20/S2_6_29  ( .A(\mult_20/ab[6][29] ), .B(
        \mult_20/CARRYB[5][29] ), .CI(\mult_20/SUMB[5][30] ), .CO(
        \mult_20/CARRYB[6][29] ), .S(\mult_20/SUMB[6][29] ) );
  FA_X1 \mult_20/S2_6_28  ( .A(\mult_20/ab[6][28] ), .B(
        \mult_20/CARRYB[5][28] ), .CI(\mult_20/SUMB[5][29] ), .CO(
        \mult_20/CARRYB[6][28] ), .S(\mult_20/SUMB[6][28] ) );
  FA_X1 \mult_20/S2_6_27  ( .A(\mult_20/ab[6][27] ), .B(
        \mult_20/CARRYB[5][27] ), .CI(\mult_20/SUMB[5][28] ), .CO(
        \mult_20/CARRYB[6][27] ), .S(\mult_20/SUMB[6][27] ) );
  FA_X1 \mult_20/S2_6_26  ( .A(\mult_20/ab[6][26] ), .B(
        \mult_20/CARRYB[5][26] ), .CI(\mult_20/SUMB[5][27] ), .CO(
        \mult_20/CARRYB[6][26] ), .S(\mult_20/SUMB[6][26] ) );
  FA_X1 \mult_20/S2_6_25  ( .A(\mult_20/ab[6][25] ), .B(
        \mult_20/CARRYB[5][25] ), .CI(\mult_20/SUMB[5][26] ), .CO(
        \mult_20/CARRYB[6][25] ), .S(\mult_20/SUMB[6][25] ) );
  FA_X1 \mult_20/S2_6_24  ( .A(\mult_20/ab[6][24] ), .B(
        \mult_20/CARRYB[5][24] ), .CI(\mult_20/SUMB[5][25] ), .CO(
        \mult_20/CARRYB[6][24] ), .S(\mult_20/SUMB[6][24] ) );
  FA_X1 \mult_20/S2_6_23  ( .A(\mult_20/ab[6][23] ), .B(
        \mult_20/CARRYB[5][23] ), .CI(\mult_20/SUMB[5][24] ), .CO(
        \mult_20/CARRYB[6][23] ), .S(\mult_20/SUMB[6][23] ) );
  FA_X1 \mult_20/S2_6_22  ( .A(\mult_20/ab[6][22] ), .B(
        \mult_20/CARRYB[5][22] ), .CI(\mult_20/SUMB[5][23] ), .CO(
        \mult_20/CARRYB[6][22] ), .S(\mult_20/SUMB[6][22] ) );
  FA_X1 \mult_20/S2_6_21  ( .A(\mult_20/ab[6][21] ), .B(
        \mult_20/CARRYB[5][21] ), .CI(\mult_20/SUMB[5][22] ), .CO(
        \mult_20/CARRYB[6][21] ), .S(\mult_20/SUMB[6][21] ) );
  FA_X1 \mult_20/S2_6_20  ( .A(\mult_20/ab[6][20] ), .B(
        \mult_20/CARRYB[5][20] ), .CI(\mult_20/SUMB[5][21] ), .CO(
        \mult_20/CARRYB[6][20] ), .S(\mult_20/SUMB[6][20] ) );
  FA_X1 \mult_20/S2_6_19  ( .A(\mult_20/ab[6][19] ), .B(
        \mult_20/CARRYB[5][19] ), .CI(\mult_20/SUMB[5][20] ), .CO(
        \mult_20/CARRYB[6][19] ), .S(\mult_20/SUMB[6][19] ) );
  FA_X1 \mult_20/S2_6_18  ( .A(\mult_20/ab[6][18] ), .B(
        \mult_20/CARRYB[5][18] ), .CI(\mult_20/SUMB[5][19] ), .CO(
        \mult_20/CARRYB[6][18] ), .S(\mult_20/SUMB[6][18] ) );
  FA_X1 \mult_20/S2_6_17  ( .A(\mult_20/ab[6][17] ), .B(
        \mult_20/CARRYB[5][17] ), .CI(\mult_20/SUMB[5][18] ), .CO(
        \mult_20/CARRYB[6][17] ), .S(\mult_20/SUMB[6][17] ) );
  FA_X1 \mult_20/S2_6_16  ( .A(\mult_20/ab[6][16] ), .B(
        \mult_20/CARRYB[5][16] ), .CI(\mult_20/SUMB[5][17] ), .CO(
        \mult_20/CARRYB[6][16] ), .S(\mult_20/SUMB[6][16] ) );
  FA_X1 \mult_20/S2_6_15  ( .A(\mult_20/ab[6][15] ), .B(
        \mult_20/CARRYB[5][15] ), .CI(\mult_20/SUMB[5][16] ), .CO(
        \mult_20/CARRYB[6][15] ), .S(\mult_20/SUMB[6][15] ) );
  FA_X1 \mult_20/S2_6_14  ( .A(\mult_20/ab[6][14] ), .B(
        \mult_20/CARRYB[5][14] ), .CI(\mult_20/SUMB[5][15] ), .CO(
        \mult_20/CARRYB[6][14] ), .S(\mult_20/SUMB[6][14] ) );
  FA_X1 \mult_20/S2_6_13  ( .A(\mult_20/ab[6][13] ), .B(
        \mult_20/CARRYB[5][13] ), .CI(\mult_20/SUMB[5][14] ), .CO(
        \mult_20/CARRYB[6][13] ), .S(\mult_20/SUMB[6][13] ) );
  FA_X1 \mult_20/S2_6_12  ( .A(\mult_20/ab[6][12] ), .B(
        \mult_20/CARRYB[5][12] ), .CI(\mult_20/SUMB[5][13] ), .CO(
        \mult_20/CARRYB[6][12] ), .S(\mult_20/SUMB[6][12] ) );
  FA_X1 \mult_20/S2_6_11  ( .A(\mult_20/ab[6][11] ), .B(
        \mult_20/CARRYB[5][11] ), .CI(\mult_20/SUMB[5][12] ), .CO(
        \mult_20/CARRYB[6][11] ), .S(\mult_20/SUMB[6][11] ) );
  FA_X1 \mult_20/S2_6_10  ( .A(\mult_20/ab[6][10] ), .B(
        \mult_20/CARRYB[5][10] ), .CI(\mult_20/SUMB[5][11] ), .CO(
        \mult_20/CARRYB[6][10] ), .S(\mult_20/SUMB[6][10] ) );
  FA_X1 \mult_20/S2_6_9  ( .A(\mult_20/ab[6][9] ), .B(\mult_20/CARRYB[5][9] ), 
        .CI(\mult_20/SUMB[5][10] ), .CO(\mult_20/CARRYB[6][9] ), .S(
        \mult_20/SUMB[6][9] ) );
  FA_X1 \mult_20/S2_6_8  ( .A(\mult_20/ab[6][8] ), .B(\mult_20/CARRYB[5][8] ), 
        .CI(\mult_20/SUMB[5][9] ), .CO(\mult_20/CARRYB[6][8] ), .S(
        \mult_20/SUMB[6][8] ) );
  FA_X1 \mult_20/S2_6_7  ( .A(\mult_20/ab[6][7] ), .B(\mult_20/CARRYB[5][7] ), 
        .CI(\mult_20/SUMB[5][8] ), .CO(\mult_20/CARRYB[6][7] ), .S(
        \mult_20/SUMB[6][7] ) );
  FA_X1 \mult_20/S2_6_6  ( .A(\mult_20/ab[6][6] ), .B(\mult_20/CARRYB[5][6] ), 
        .CI(\mult_20/SUMB[5][7] ), .CO(\mult_20/CARRYB[6][6] ), .S(
        \mult_20/SUMB[6][6] ) );
  FA_X1 \mult_20/S2_6_5  ( .A(\mult_20/ab[6][5] ), .B(\mult_20/CARRYB[5][5] ), 
        .CI(\mult_20/SUMB[5][6] ), .CO(\mult_20/CARRYB[6][5] ), .S(
        \mult_20/SUMB[6][5] ) );
  FA_X1 \mult_20/S2_6_4  ( .A(\mult_20/ab[6][4] ), .B(\mult_20/CARRYB[5][4] ), 
        .CI(\mult_20/SUMB[5][5] ), .CO(\mult_20/CARRYB[6][4] ), .S(
        \mult_20/SUMB[6][4] ) );
  FA_X1 \mult_20/S2_6_3  ( .A(\mult_20/ab[6][3] ), .B(\mult_20/CARRYB[5][3] ), 
        .CI(\mult_20/SUMB[5][4] ), .CO(\mult_20/CARRYB[6][3] ), .S(
        \mult_20/SUMB[6][3] ) );
  FA_X1 \mult_20/S2_6_2  ( .A(\mult_20/ab[6][2] ), .B(\mult_20/CARRYB[5][2] ), 
        .CI(\mult_20/SUMB[5][3] ), .CO(\mult_20/CARRYB[6][2] ), .S(
        \mult_20/SUMB[6][2] ) );
  FA_X1 \mult_20/S2_6_1  ( .A(\mult_20/ab[6][1] ), .B(\mult_20/CARRYB[5][1] ), 
        .CI(\mult_20/SUMB[5][2] ), .CO(\mult_20/CARRYB[6][1] ), .S(
        \mult_20/SUMB[6][1] ) );
  FA_X1 \mult_20/S1_6_0  ( .A(\mult_20/ab[6][0] ), .B(\mult_20/CARRYB[5][0] ), 
        .CI(\mult_20/SUMB[5][1] ), .CO(\mult_20/CARRYB[6][0] ), .S(N70) );
  FA_X1 \mult_20/S3_7_30  ( .A(\mult_20/ab[7][30] ), .B(
        \mult_20/CARRYB[6][30] ), .CI(\mult_20/ab[6][31] ), .CO(
        \mult_20/CARRYB[7][30] ), .S(\mult_20/SUMB[7][30] ) );
  FA_X1 \mult_20/S2_7_29  ( .A(\mult_20/ab[7][29] ), .B(
        \mult_20/CARRYB[6][29] ), .CI(\mult_20/SUMB[6][30] ), .CO(
        \mult_20/CARRYB[7][29] ), .S(\mult_20/SUMB[7][29] ) );
  FA_X1 \mult_20/S2_7_28  ( .A(\mult_20/ab[7][28] ), .B(
        \mult_20/CARRYB[6][28] ), .CI(\mult_20/SUMB[6][29] ), .CO(
        \mult_20/CARRYB[7][28] ), .S(\mult_20/SUMB[7][28] ) );
  FA_X1 \mult_20/S2_7_27  ( .A(\mult_20/ab[7][27] ), .B(
        \mult_20/CARRYB[6][27] ), .CI(\mult_20/SUMB[6][28] ), .CO(
        \mult_20/CARRYB[7][27] ), .S(\mult_20/SUMB[7][27] ) );
  FA_X1 \mult_20/S2_7_26  ( .A(\mult_20/ab[7][26] ), .B(
        \mult_20/CARRYB[6][26] ), .CI(\mult_20/SUMB[6][27] ), .CO(
        \mult_20/CARRYB[7][26] ), .S(\mult_20/SUMB[7][26] ) );
  FA_X1 \mult_20/S2_7_25  ( .A(\mult_20/ab[7][25] ), .B(
        \mult_20/CARRYB[6][25] ), .CI(\mult_20/SUMB[6][26] ), .CO(
        \mult_20/CARRYB[7][25] ), .S(\mult_20/SUMB[7][25] ) );
  FA_X1 \mult_20/S2_7_24  ( .A(\mult_20/ab[7][24] ), .B(
        \mult_20/CARRYB[6][24] ), .CI(\mult_20/SUMB[6][25] ), .CO(
        \mult_20/CARRYB[7][24] ), .S(\mult_20/SUMB[7][24] ) );
  FA_X1 \mult_20/S2_7_23  ( .A(\mult_20/ab[7][23] ), .B(
        \mult_20/CARRYB[6][23] ), .CI(\mult_20/SUMB[6][24] ), .CO(
        \mult_20/CARRYB[7][23] ), .S(\mult_20/SUMB[7][23] ) );
  FA_X1 \mult_20/S2_7_22  ( .A(\mult_20/ab[7][22] ), .B(
        \mult_20/CARRYB[6][22] ), .CI(\mult_20/SUMB[6][23] ), .CO(
        \mult_20/CARRYB[7][22] ), .S(\mult_20/SUMB[7][22] ) );
  FA_X1 \mult_20/S2_7_21  ( .A(\mult_20/ab[7][21] ), .B(
        \mult_20/CARRYB[6][21] ), .CI(\mult_20/SUMB[6][22] ), .CO(
        \mult_20/CARRYB[7][21] ), .S(\mult_20/SUMB[7][21] ) );
  FA_X1 \mult_20/S2_7_20  ( .A(\mult_20/ab[7][20] ), .B(
        \mult_20/CARRYB[6][20] ), .CI(\mult_20/SUMB[6][21] ), .CO(
        \mult_20/CARRYB[7][20] ), .S(\mult_20/SUMB[7][20] ) );
  FA_X1 \mult_20/S2_7_19  ( .A(\mult_20/ab[7][19] ), .B(
        \mult_20/CARRYB[6][19] ), .CI(\mult_20/SUMB[6][20] ), .CO(
        \mult_20/CARRYB[7][19] ), .S(\mult_20/SUMB[7][19] ) );
  FA_X1 \mult_20/S2_7_18  ( .A(\mult_20/ab[7][18] ), .B(
        \mult_20/CARRYB[6][18] ), .CI(\mult_20/SUMB[6][19] ), .CO(
        \mult_20/CARRYB[7][18] ), .S(\mult_20/SUMB[7][18] ) );
  FA_X1 \mult_20/S2_7_17  ( .A(\mult_20/ab[7][17] ), .B(
        \mult_20/CARRYB[6][17] ), .CI(\mult_20/SUMB[6][18] ), .CO(
        \mult_20/CARRYB[7][17] ), .S(\mult_20/SUMB[7][17] ) );
  FA_X1 \mult_20/S2_7_16  ( .A(\mult_20/ab[7][16] ), .B(
        \mult_20/CARRYB[6][16] ), .CI(\mult_20/SUMB[6][17] ), .CO(
        \mult_20/CARRYB[7][16] ), .S(\mult_20/SUMB[7][16] ) );
  FA_X1 \mult_20/S2_7_15  ( .A(\mult_20/ab[7][15] ), .B(
        \mult_20/CARRYB[6][15] ), .CI(\mult_20/SUMB[6][16] ), .CO(
        \mult_20/CARRYB[7][15] ), .S(\mult_20/SUMB[7][15] ) );
  FA_X1 \mult_20/S2_7_14  ( .A(\mult_20/ab[7][14] ), .B(
        \mult_20/CARRYB[6][14] ), .CI(\mult_20/SUMB[6][15] ), .CO(
        \mult_20/CARRYB[7][14] ), .S(\mult_20/SUMB[7][14] ) );
  FA_X1 \mult_20/S2_7_13  ( .A(\mult_20/ab[7][13] ), .B(
        \mult_20/CARRYB[6][13] ), .CI(\mult_20/SUMB[6][14] ), .CO(
        \mult_20/CARRYB[7][13] ), .S(\mult_20/SUMB[7][13] ) );
  FA_X1 \mult_20/S2_7_12  ( .A(\mult_20/ab[7][12] ), .B(
        \mult_20/CARRYB[6][12] ), .CI(\mult_20/SUMB[6][13] ), .CO(
        \mult_20/CARRYB[7][12] ), .S(\mult_20/SUMB[7][12] ) );
  FA_X1 \mult_20/S2_7_11  ( .A(\mult_20/ab[7][11] ), .B(
        \mult_20/CARRYB[6][11] ), .CI(\mult_20/SUMB[6][12] ), .CO(
        \mult_20/CARRYB[7][11] ), .S(\mult_20/SUMB[7][11] ) );
  FA_X1 \mult_20/S2_7_10  ( .A(\mult_20/ab[7][10] ), .B(
        \mult_20/CARRYB[6][10] ), .CI(\mult_20/SUMB[6][11] ), .CO(
        \mult_20/CARRYB[7][10] ), .S(\mult_20/SUMB[7][10] ) );
  FA_X1 \mult_20/S2_7_9  ( .A(\mult_20/ab[7][9] ), .B(\mult_20/CARRYB[6][9] ), 
        .CI(\mult_20/SUMB[6][10] ), .CO(\mult_20/CARRYB[7][9] ), .S(
        \mult_20/SUMB[7][9] ) );
  FA_X1 \mult_20/S2_7_8  ( .A(\mult_20/ab[7][8] ), .B(\mult_20/CARRYB[6][8] ), 
        .CI(\mult_20/SUMB[6][9] ), .CO(\mult_20/CARRYB[7][8] ), .S(
        \mult_20/SUMB[7][8] ) );
  FA_X1 \mult_20/S2_7_7  ( .A(\mult_20/ab[7][7] ), .B(\mult_20/CARRYB[6][7] ), 
        .CI(\mult_20/SUMB[6][8] ), .CO(\mult_20/CARRYB[7][7] ), .S(
        \mult_20/SUMB[7][7] ) );
  FA_X1 \mult_20/S2_7_6  ( .A(\mult_20/ab[7][6] ), .B(\mult_20/CARRYB[6][6] ), 
        .CI(\mult_20/SUMB[6][7] ), .CO(\mult_20/CARRYB[7][6] ), .S(
        \mult_20/SUMB[7][6] ) );
  FA_X1 \mult_20/S2_7_5  ( .A(\mult_20/ab[7][5] ), .B(\mult_20/CARRYB[6][5] ), 
        .CI(\mult_20/SUMB[6][6] ), .CO(\mult_20/CARRYB[7][5] ), .S(
        \mult_20/SUMB[7][5] ) );
  FA_X1 \mult_20/S2_7_4  ( .A(\mult_20/ab[7][4] ), .B(\mult_20/CARRYB[6][4] ), 
        .CI(\mult_20/SUMB[6][5] ), .CO(\mult_20/CARRYB[7][4] ), .S(
        \mult_20/SUMB[7][4] ) );
  FA_X1 \mult_20/S2_7_3  ( .A(\mult_20/ab[7][3] ), .B(\mult_20/CARRYB[6][3] ), 
        .CI(\mult_20/SUMB[6][4] ), .CO(\mult_20/CARRYB[7][3] ), .S(
        \mult_20/SUMB[7][3] ) );
  FA_X1 \mult_20/S2_7_2  ( .A(\mult_20/ab[7][2] ), .B(\mult_20/CARRYB[6][2] ), 
        .CI(\mult_20/SUMB[6][3] ), .CO(\mult_20/CARRYB[7][2] ), .S(
        \mult_20/SUMB[7][2] ) );
  FA_X1 \mult_20/S2_7_1  ( .A(\mult_20/ab[7][1] ), .B(\mult_20/CARRYB[6][1] ), 
        .CI(\mult_20/SUMB[6][2] ), .CO(\mult_20/CARRYB[7][1] ), .S(
        \mult_20/SUMB[7][1] ) );
  FA_X1 \mult_20/S1_7_0  ( .A(\mult_20/ab[7][0] ), .B(\mult_20/CARRYB[6][0] ), 
        .CI(\mult_20/SUMB[6][1] ), .CO(\mult_20/CARRYB[7][0] ), .S(N71) );
  FA_X1 \mult_20/S3_8_30  ( .A(\mult_20/ab[8][30] ), .B(
        \mult_20/CARRYB[7][30] ), .CI(\mult_20/ab[7][31] ), .CO(
        \mult_20/CARRYB[8][30] ), .S(\mult_20/SUMB[8][30] ) );
  FA_X1 \mult_20/S2_8_29  ( .A(\mult_20/ab[8][29] ), .B(
        \mult_20/CARRYB[7][29] ), .CI(\mult_20/SUMB[7][30] ), .CO(
        \mult_20/CARRYB[8][29] ), .S(\mult_20/SUMB[8][29] ) );
  FA_X1 \mult_20/S2_8_28  ( .A(\mult_20/ab[8][28] ), .B(
        \mult_20/CARRYB[7][28] ), .CI(\mult_20/SUMB[7][29] ), .CO(
        \mult_20/CARRYB[8][28] ), .S(\mult_20/SUMB[8][28] ) );
  FA_X1 \mult_20/S2_8_27  ( .A(\mult_20/ab[8][27] ), .B(
        \mult_20/CARRYB[7][27] ), .CI(\mult_20/SUMB[7][28] ), .CO(
        \mult_20/CARRYB[8][27] ), .S(\mult_20/SUMB[8][27] ) );
  FA_X1 \mult_20/S2_8_26  ( .A(\mult_20/ab[8][26] ), .B(
        \mult_20/CARRYB[7][26] ), .CI(\mult_20/SUMB[7][27] ), .CO(
        \mult_20/CARRYB[8][26] ), .S(\mult_20/SUMB[8][26] ) );
  FA_X1 \mult_20/S2_8_25  ( .A(\mult_20/ab[8][25] ), .B(
        \mult_20/CARRYB[7][25] ), .CI(\mult_20/SUMB[7][26] ), .CO(
        \mult_20/CARRYB[8][25] ), .S(\mult_20/SUMB[8][25] ) );
  FA_X1 \mult_20/S2_8_24  ( .A(\mult_20/ab[8][24] ), .B(
        \mult_20/CARRYB[7][24] ), .CI(\mult_20/SUMB[7][25] ), .CO(
        \mult_20/CARRYB[8][24] ), .S(\mult_20/SUMB[8][24] ) );
  FA_X1 \mult_20/S2_8_23  ( .A(\mult_20/ab[8][23] ), .B(
        \mult_20/CARRYB[7][23] ), .CI(\mult_20/SUMB[7][24] ), .CO(
        \mult_20/CARRYB[8][23] ), .S(\mult_20/SUMB[8][23] ) );
  FA_X1 \mult_20/S2_8_22  ( .A(\mult_20/ab[8][22] ), .B(
        \mult_20/CARRYB[7][22] ), .CI(\mult_20/SUMB[7][23] ), .CO(
        \mult_20/CARRYB[8][22] ), .S(\mult_20/SUMB[8][22] ) );
  FA_X1 \mult_20/S2_8_21  ( .A(\mult_20/ab[8][21] ), .B(
        \mult_20/CARRYB[7][21] ), .CI(\mult_20/SUMB[7][22] ), .CO(
        \mult_20/CARRYB[8][21] ), .S(\mult_20/SUMB[8][21] ) );
  FA_X1 \mult_20/S2_8_20  ( .A(\mult_20/ab[8][20] ), .B(
        \mult_20/CARRYB[7][20] ), .CI(\mult_20/SUMB[7][21] ), .CO(
        \mult_20/CARRYB[8][20] ), .S(\mult_20/SUMB[8][20] ) );
  FA_X1 \mult_20/S2_8_19  ( .A(\mult_20/ab[8][19] ), .B(
        \mult_20/CARRYB[7][19] ), .CI(\mult_20/SUMB[7][20] ), .CO(
        \mult_20/CARRYB[8][19] ), .S(\mult_20/SUMB[8][19] ) );
  FA_X1 \mult_20/S2_8_18  ( .A(\mult_20/ab[8][18] ), .B(
        \mult_20/CARRYB[7][18] ), .CI(\mult_20/SUMB[7][19] ), .CO(
        \mult_20/CARRYB[8][18] ), .S(\mult_20/SUMB[8][18] ) );
  FA_X1 \mult_20/S2_8_17  ( .A(\mult_20/ab[8][17] ), .B(
        \mult_20/CARRYB[7][17] ), .CI(\mult_20/SUMB[7][18] ), .CO(
        \mult_20/CARRYB[8][17] ), .S(\mult_20/SUMB[8][17] ) );
  FA_X1 \mult_20/S2_8_16  ( .A(\mult_20/ab[8][16] ), .B(
        \mult_20/CARRYB[7][16] ), .CI(\mult_20/SUMB[7][17] ), .CO(
        \mult_20/CARRYB[8][16] ), .S(\mult_20/SUMB[8][16] ) );
  FA_X1 \mult_20/S2_8_15  ( .A(\mult_20/ab[8][15] ), .B(
        \mult_20/CARRYB[7][15] ), .CI(\mult_20/SUMB[7][16] ), .CO(
        \mult_20/CARRYB[8][15] ), .S(\mult_20/SUMB[8][15] ) );
  FA_X1 \mult_20/S2_8_14  ( .A(\mult_20/ab[8][14] ), .B(
        \mult_20/CARRYB[7][14] ), .CI(\mult_20/SUMB[7][15] ), .CO(
        \mult_20/CARRYB[8][14] ), .S(\mult_20/SUMB[8][14] ) );
  FA_X1 \mult_20/S2_8_13  ( .A(\mult_20/ab[8][13] ), .B(
        \mult_20/CARRYB[7][13] ), .CI(\mult_20/SUMB[7][14] ), .CO(
        \mult_20/CARRYB[8][13] ), .S(\mult_20/SUMB[8][13] ) );
  FA_X1 \mult_20/S2_8_12  ( .A(\mult_20/ab[8][12] ), .B(
        \mult_20/CARRYB[7][12] ), .CI(\mult_20/SUMB[7][13] ), .CO(
        \mult_20/CARRYB[8][12] ), .S(\mult_20/SUMB[8][12] ) );
  FA_X1 \mult_20/S2_8_11  ( .A(\mult_20/ab[8][11] ), .B(
        \mult_20/CARRYB[7][11] ), .CI(\mult_20/SUMB[7][12] ), .CO(
        \mult_20/CARRYB[8][11] ), .S(\mult_20/SUMB[8][11] ) );
  FA_X1 \mult_20/S2_8_10  ( .A(\mult_20/ab[8][10] ), .B(
        \mult_20/CARRYB[7][10] ), .CI(\mult_20/SUMB[7][11] ), .CO(
        \mult_20/CARRYB[8][10] ), .S(\mult_20/SUMB[8][10] ) );
  FA_X1 \mult_20/S2_8_9  ( .A(\mult_20/ab[8][9] ), .B(\mult_20/CARRYB[7][9] ), 
        .CI(\mult_20/SUMB[7][10] ), .CO(\mult_20/CARRYB[8][9] ), .S(
        \mult_20/SUMB[8][9] ) );
  FA_X1 \mult_20/S2_8_8  ( .A(\mult_20/ab[8][8] ), .B(\mult_20/CARRYB[7][8] ), 
        .CI(\mult_20/SUMB[7][9] ), .CO(\mult_20/CARRYB[8][8] ), .S(
        \mult_20/SUMB[8][8] ) );
  FA_X1 \mult_20/S2_8_7  ( .A(\mult_20/ab[8][7] ), .B(\mult_20/CARRYB[7][7] ), 
        .CI(\mult_20/SUMB[7][8] ), .CO(\mult_20/CARRYB[8][7] ), .S(
        \mult_20/SUMB[8][7] ) );
  FA_X1 \mult_20/S2_8_6  ( .A(\mult_20/ab[8][6] ), .B(\mult_20/CARRYB[7][6] ), 
        .CI(\mult_20/SUMB[7][7] ), .CO(\mult_20/CARRYB[8][6] ), .S(
        \mult_20/SUMB[8][6] ) );
  FA_X1 \mult_20/S2_8_5  ( .A(\mult_20/ab[8][5] ), .B(\mult_20/CARRYB[7][5] ), 
        .CI(\mult_20/SUMB[7][6] ), .CO(\mult_20/CARRYB[8][5] ), .S(
        \mult_20/SUMB[8][5] ) );
  FA_X1 \mult_20/S2_8_4  ( .A(\mult_20/ab[8][4] ), .B(\mult_20/CARRYB[7][4] ), 
        .CI(\mult_20/SUMB[7][5] ), .CO(\mult_20/CARRYB[8][4] ), .S(
        \mult_20/SUMB[8][4] ) );
  FA_X1 \mult_20/S2_8_3  ( .A(\mult_20/ab[8][3] ), .B(\mult_20/CARRYB[7][3] ), 
        .CI(\mult_20/SUMB[7][4] ), .CO(\mult_20/CARRYB[8][3] ), .S(
        \mult_20/SUMB[8][3] ) );
  FA_X1 \mult_20/S2_8_2  ( .A(\mult_20/ab[8][2] ), .B(\mult_20/CARRYB[7][2] ), 
        .CI(\mult_20/SUMB[7][3] ), .CO(\mult_20/CARRYB[8][2] ), .S(
        \mult_20/SUMB[8][2] ) );
  FA_X1 \mult_20/S2_8_1  ( .A(\mult_20/ab[8][1] ), .B(\mult_20/CARRYB[7][1] ), 
        .CI(\mult_20/SUMB[7][2] ), .CO(\mult_20/CARRYB[8][1] ), .S(
        \mult_20/SUMB[8][1] ) );
  FA_X1 \mult_20/S1_8_0  ( .A(\mult_20/ab[8][0] ), .B(\mult_20/CARRYB[7][0] ), 
        .CI(\mult_20/SUMB[7][1] ), .CO(\mult_20/CARRYB[8][0] ), .S(N72) );
  FA_X1 \mult_20/S3_9_30  ( .A(\mult_20/ab[9][30] ), .B(
        \mult_20/CARRYB[8][30] ), .CI(\mult_20/ab[8][31] ), .CO(
        \mult_20/CARRYB[9][30] ), .S(\mult_20/SUMB[9][30] ) );
  FA_X1 \mult_20/S2_9_29  ( .A(\mult_20/ab[9][29] ), .B(
        \mult_20/CARRYB[8][29] ), .CI(\mult_20/SUMB[8][30] ), .CO(
        \mult_20/CARRYB[9][29] ), .S(\mult_20/SUMB[9][29] ) );
  FA_X1 \mult_20/S2_9_28  ( .A(\mult_20/ab[9][28] ), .B(
        \mult_20/CARRYB[8][28] ), .CI(\mult_20/SUMB[8][29] ), .CO(
        \mult_20/CARRYB[9][28] ), .S(\mult_20/SUMB[9][28] ) );
  FA_X1 \mult_20/S2_9_27  ( .A(\mult_20/ab[9][27] ), .B(
        \mult_20/CARRYB[8][27] ), .CI(\mult_20/SUMB[8][28] ), .CO(
        \mult_20/CARRYB[9][27] ), .S(\mult_20/SUMB[9][27] ) );
  FA_X1 \mult_20/S2_9_26  ( .A(\mult_20/ab[9][26] ), .B(
        \mult_20/CARRYB[8][26] ), .CI(\mult_20/SUMB[8][27] ), .CO(
        \mult_20/CARRYB[9][26] ), .S(\mult_20/SUMB[9][26] ) );
  FA_X1 \mult_20/S2_9_25  ( .A(\mult_20/ab[9][25] ), .B(
        \mult_20/CARRYB[8][25] ), .CI(\mult_20/SUMB[8][26] ), .CO(
        \mult_20/CARRYB[9][25] ), .S(\mult_20/SUMB[9][25] ) );
  FA_X1 \mult_20/S2_9_24  ( .A(\mult_20/ab[9][24] ), .B(
        \mult_20/CARRYB[8][24] ), .CI(\mult_20/SUMB[8][25] ), .CO(
        \mult_20/CARRYB[9][24] ), .S(\mult_20/SUMB[9][24] ) );
  FA_X1 \mult_20/S2_9_23  ( .A(\mult_20/ab[9][23] ), .B(
        \mult_20/CARRYB[8][23] ), .CI(\mult_20/SUMB[8][24] ), .CO(
        \mult_20/CARRYB[9][23] ), .S(\mult_20/SUMB[9][23] ) );
  FA_X1 \mult_20/S2_9_22  ( .A(\mult_20/ab[9][22] ), .B(
        \mult_20/CARRYB[8][22] ), .CI(\mult_20/SUMB[8][23] ), .CO(
        \mult_20/CARRYB[9][22] ), .S(\mult_20/SUMB[9][22] ) );
  FA_X1 \mult_20/S2_9_21  ( .A(\mult_20/ab[9][21] ), .B(
        \mult_20/CARRYB[8][21] ), .CI(\mult_20/SUMB[8][22] ), .CO(
        \mult_20/CARRYB[9][21] ), .S(\mult_20/SUMB[9][21] ) );
  FA_X1 \mult_20/S2_9_20  ( .A(\mult_20/ab[9][20] ), .B(
        \mult_20/CARRYB[8][20] ), .CI(\mult_20/SUMB[8][21] ), .CO(
        \mult_20/CARRYB[9][20] ), .S(\mult_20/SUMB[9][20] ) );
  FA_X1 \mult_20/S2_9_19  ( .A(\mult_20/ab[9][19] ), .B(
        \mult_20/CARRYB[8][19] ), .CI(\mult_20/SUMB[8][20] ), .CO(
        \mult_20/CARRYB[9][19] ), .S(\mult_20/SUMB[9][19] ) );
  FA_X1 \mult_20/S2_9_18  ( .A(\mult_20/ab[9][18] ), .B(
        \mult_20/CARRYB[8][18] ), .CI(\mult_20/SUMB[8][19] ), .CO(
        \mult_20/CARRYB[9][18] ), .S(\mult_20/SUMB[9][18] ) );
  FA_X1 \mult_20/S2_9_17  ( .A(\mult_20/ab[9][17] ), .B(
        \mult_20/CARRYB[8][17] ), .CI(\mult_20/SUMB[8][18] ), .CO(
        \mult_20/CARRYB[9][17] ), .S(\mult_20/SUMB[9][17] ) );
  FA_X1 \mult_20/S2_9_16  ( .A(\mult_20/ab[9][16] ), .B(
        \mult_20/CARRYB[8][16] ), .CI(\mult_20/SUMB[8][17] ), .CO(
        \mult_20/CARRYB[9][16] ), .S(\mult_20/SUMB[9][16] ) );
  FA_X1 \mult_20/S2_9_15  ( .A(\mult_20/ab[9][15] ), .B(
        \mult_20/CARRYB[8][15] ), .CI(\mult_20/SUMB[8][16] ), .CO(
        \mult_20/CARRYB[9][15] ), .S(\mult_20/SUMB[9][15] ) );
  FA_X1 \mult_20/S2_9_14  ( .A(\mult_20/ab[9][14] ), .B(
        \mult_20/CARRYB[8][14] ), .CI(\mult_20/SUMB[8][15] ), .CO(
        \mult_20/CARRYB[9][14] ), .S(\mult_20/SUMB[9][14] ) );
  FA_X1 \mult_20/S2_9_13  ( .A(\mult_20/ab[9][13] ), .B(
        \mult_20/CARRYB[8][13] ), .CI(\mult_20/SUMB[8][14] ), .CO(
        \mult_20/CARRYB[9][13] ), .S(\mult_20/SUMB[9][13] ) );
  FA_X1 \mult_20/S2_9_12  ( .A(\mult_20/ab[9][12] ), .B(
        \mult_20/CARRYB[8][12] ), .CI(\mult_20/SUMB[8][13] ), .CO(
        \mult_20/CARRYB[9][12] ), .S(\mult_20/SUMB[9][12] ) );
  FA_X1 \mult_20/S2_9_11  ( .A(\mult_20/ab[9][11] ), .B(
        \mult_20/CARRYB[8][11] ), .CI(\mult_20/SUMB[8][12] ), .CO(
        \mult_20/CARRYB[9][11] ), .S(\mult_20/SUMB[9][11] ) );
  FA_X1 \mult_20/S2_9_10  ( .A(\mult_20/ab[9][10] ), .B(
        \mult_20/CARRYB[8][10] ), .CI(\mult_20/SUMB[8][11] ), .CO(
        \mult_20/CARRYB[9][10] ), .S(\mult_20/SUMB[9][10] ) );
  FA_X1 \mult_20/S2_9_9  ( .A(\mult_20/ab[9][9] ), .B(\mult_20/CARRYB[8][9] ), 
        .CI(\mult_20/SUMB[8][10] ), .CO(\mult_20/CARRYB[9][9] ), .S(
        \mult_20/SUMB[9][9] ) );
  FA_X1 \mult_20/S2_9_8  ( .A(\mult_20/ab[9][8] ), .B(\mult_20/CARRYB[8][8] ), 
        .CI(\mult_20/SUMB[8][9] ), .CO(\mult_20/CARRYB[9][8] ), .S(
        \mult_20/SUMB[9][8] ) );
  FA_X1 \mult_20/S2_9_7  ( .A(\mult_20/ab[9][7] ), .B(\mult_20/CARRYB[8][7] ), 
        .CI(\mult_20/SUMB[8][8] ), .CO(\mult_20/CARRYB[9][7] ), .S(
        \mult_20/SUMB[9][7] ) );
  FA_X1 \mult_20/S2_9_6  ( .A(\mult_20/ab[9][6] ), .B(\mult_20/CARRYB[8][6] ), 
        .CI(\mult_20/SUMB[8][7] ), .CO(\mult_20/CARRYB[9][6] ), .S(
        \mult_20/SUMB[9][6] ) );
  FA_X1 \mult_20/S2_9_5  ( .A(\mult_20/ab[9][5] ), .B(\mult_20/CARRYB[8][5] ), 
        .CI(\mult_20/SUMB[8][6] ), .CO(\mult_20/CARRYB[9][5] ), .S(
        \mult_20/SUMB[9][5] ) );
  FA_X1 \mult_20/S2_9_4  ( .A(\mult_20/ab[9][4] ), .B(\mult_20/CARRYB[8][4] ), 
        .CI(\mult_20/SUMB[8][5] ), .CO(\mult_20/CARRYB[9][4] ), .S(
        \mult_20/SUMB[9][4] ) );
  FA_X1 \mult_20/S2_9_3  ( .A(\mult_20/ab[9][3] ), .B(\mult_20/CARRYB[8][3] ), 
        .CI(\mult_20/SUMB[8][4] ), .CO(\mult_20/CARRYB[9][3] ), .S(
        \mult_20/SUMB[9][3] ) );
  FA_X1 \mult_20/S2_9_2  ( .A(\mult_20/ab[9][2] ), .B(\mult_20/CARRYB[8][2] ), 
        .CI(\mult_20/SUMB[8][3] ), .CO(\mult_20/CARRYB[9][2] ), .S(
        \mult_20/SUMB[9][2] ) );
  FA_X1 \mult_20/S2_9_1  ( .A(\mult_20/ab[9][1] ), .B(\mult_20/CARRYB[8][1] ), 
        .CI(\mult_20/SUMB[8][2] ), .CO(\mult_20/CARRYB[9][1] ), .S(
        \mult_20/SUMB[9][1] ) );
  FA_X1 \mult_20/S1_9_0  ( .A(\mult_20/ab[9][0] ), .B(\mult_20/CARRYB[8][0] ), 
        .CI(\mult_20/SUMB[8][1] ), .CO(\mult_20/CARRYB[9][0] ), .S(N73) );
  FA_X1 \mult_20/S3_10_30  ( .A(\mult_20/ab[10][30] ), .B(
        \mult_20/CARRYB[9][30] ), .CI(\mult_20/ab[9][31] ), .CO(
        \mult_20/CARRYB[10][30] ), .S(\mult_20/SUMB[10][30] ) );
  FA_X1 \mult_20/S2_10_29  ( .A(\mult_20/ab[10][29] ), .B(
        \mult_20/CARRYB[9][29] ), .CI(\mult_20/SUMB[9][30] ), .CO(
        \mult_20/CARRYB[10][29] ), .S(\mult_20/SUMB[10][29] ) );
  FA_X1 \mult_20/S2_10_28  ( .A(\mult_20/ab[10][28] ), .B(
        \mult_20/CARRYB[9][28] ), .CI(\mult_20/SUMB[9][29] ), .CO(
        \mult_20/CARRYB[10][28] ), .S(\mult_20/SUMB[10][28] ) );
  FA_X1 \mult_20/S2_10_27  ( .A(\mult_20/ab[10][27] ), .B(
        \mult_20/CARRYB[9][27] ), .CI(\mult_20/SUMB[9][28] ), .CO(
        \mult_20/CARRYB[10][27] ), .S(\mult_20/SUMB[10][27] ) );
  FA_X1 \mult_20/S2_10_26  ( .A(\mult_20/ab[10][26] ), .B(
        \mult_20/CARRYB[9][26] ), .CI(\mult_20/SUMB[9][27] ), .CO(
        \mult_20/CARRYB[10][26] ), .S(\mult_20/SUMB[10][26] ) );
  FA_X1 \mult_20/S2_10_25  ( .A(\mult_20/ab[10][25] ), .B(
        \mult_20/CARRYB[9][25] ), .CI(\mult_20/SUMB[9][26] ), .CO(
        \mult_20/CARRYB[10][25] ), .S(\mult_20/SUMB[10][25] ) );
  FA_X1 \mult_20/S2_10_24  ( .A(\mult_20/ab[10][24] ), .B(
        \mult_20/CARRYB[9][24] ), .CI(\mult_20/SUMB[9][25] ), .CO(
        \mult_20/CARRYB[10][24] ), .S(\mult_20/SUMB[10][24] ) );
  FA_X1 \mult_20/S2_10_23  ( .A(\mult_20/ab[10][23] ), .B(
        \mult_20/CARRYB[9][23] ), .CI(\mult_20/SUMB[9][24] ), .CO(
        \mult_20/CARRYB[10][23] ), .S(\mult_20/SUMB[10][23] ) );
  FA_X1 \mult_20/S2_10_22  ( .A(\mult_20/ab[10][22] ), .B(
        \mult_20/CARRYB[9][22] ), .CI(\mult_20/SUMB[9][23] ), .CO(
        \mult_20/CARRYB[10][22] ), .S(\mult_20/SUMB[10][22] ) );
  FA_X1 \mult_20/S2_10_21  ( .A(\mult_20/ab[10][21] ), .B(
        \mult_20/CARRYB[9][21] ), .CI(\mult_20/SUMB[9][22] ), .CO(
        \mult_20/CARRYB[10][21] ), .S(\mult_20/SUMB[10][21] ) );
  FA_X1 \mult_20/S2_10_20  ( .A(\mult_20/ab[10][20] ), .B(
        \mult_20/CARRYB[9][20] ), .CI(\mult_20/SUMB[9][21] ), .CO(
        \mult_20/CARRYB[10][20] ), .S(\mult_20/SUMB[10][20] ) );
  FA_X1 \mult_20/S2_10_19  ( .A(\mult_20/ab[10][19] ), .B(
        \mult_20/CARRYB[9][19] ), .CI(\mult_20/SUMB[9][20] ), .CO(
        \mult_20/CARRYB[10][19] ), .S(\mult_20/SUMB[10][19] ) );
  FA_X1 \mult_20/S2_10_18  ( .A(\mult_20/ab[10][18] ), .B(
        \mult_20/CARRYB[9][18] ), .CI(\mult_20/SUMB[9][19] ), .CO(
        \mult_20/CARRYB[10][18] ), .S(\mult_20/SUMB[10][18] ) );
  FA_X1 \mult_20/S2_10_17  ( .A(\mult_20/ab[10][17] ), .B(
        \mult_20/CARRYB[9][17] ), .CI(\mult_20/SUMB[9][18] ), .CO(
        \mult_20/CARRYB[10][17] ), .S(\mult_20/SUMB[10][17] ) );
  FA_X1 \mult_20/S2_10_16  ( .A(\mult_20/ab[10][16] ), .B(
        \mult_20/CARRYB[9][16] ), .CI(\mult_20/SUMB[9][17] ), .CO(
        \mult_20/CARRYB[10][16] ), .S(\mult_20/SUMB[10][16] ) );
  FA_X1 \mult_20/S2_10_15  ( .A(\mult_20/ab[10][15] ), .B(
        \mult_20/CARRYB[9][15] ), .CI(\mult_20/SUMB[9][16] ), .CO(
        \mult_20/CARRYB[10][15] ), .S(\mult_20/SUMB[10][15] ) );
  FA_X1 \mult_20/S2_10_14  ( .A(\mult_20/ab[10][14] ), .B(
        \mult_20/CARRYB[9][14] ), .CI(\mult_20/SUMB[9][15] ), .CO(
        \mult_20/CARRYB[10][14] ), .S(\mult_20/SUMB[10][14] ) );
  FA_X1 \mult_20/S2_10_13  ( .A(\mult_20/ab[10][13] ), .B(
        \mult_20/CARRYB[9][13] ), .CI(\mult_20/SUMB[9][14] ), .CO(
        \mult_20/CARRYB[10][13] ), .S(\mult_20/SUMB[10][13] ) );
  FA_X1 \mult_20/S2_10_12  ( .A(\mult_20/ab[10][12] ), .B(
        \mult_20/CARRYB[9][12] ), .CI(\mult_20/SUMB[9][13] ), .CO(
        \mult_20/CARRYB[10][12] ), .S(\mult_20/SUMB[10][12] ) );
  FA_X1 \mult_20/S2_10_11  ( .A(\mult_20/ab[10][11] ), .B(
        \mult_20/CARRYB[9][11] ), .CI(\mult_20/SUMB[9][12] ), .CO(
        \mult_20/CARRYB[10][11] ), .S(\mult_20/SUMB[10][11] ) );
  FA_X1 \mult_20/S2_10_10  ( .A(\mult_20/ab[10][10] ), .B(
        \mult_20/CARRYB[9][10] ), .CI(\mult_20/SUMB[9][11] ), .CO(
        \mult_20/CARRYB[10][10] ), .S(\mult_20/SUMB[10][10] ) );
  FA_X1 \mult_20/S2_10_9  ( .A(\mult_20/ab[10][9] ), .B(\mult_20/CARRYB[9][9] ), .CI(\mult_20/SUMB[9][10] ), .CO(\mult_20/CARRYB[10][9] ), .S(
        \mult_20/SUMB[10][9] ) );
  FA_X1 \mult_20/S2_10_8  ( .A(\mult_20/ab[10][8] ), .B(\mult_20/CARRYB[9][8] ), .CI(\mult_20/SUMB[9][9] ), .CO(\mult_20/CARRYB[10][8] ), .S(
        \mult_20/SUMB[10][8] ) );
  FA_X1 \mult_20/S2_10_7  ( .A(\mult_20/ab[10][7] ), .B(\mult_20/CARRYB[9][7] ), .CI(\mult_20/SUMB[9][8] ), .CO(\mult_20/CARRYB[10][7] ), .S(
        \mult_20/SUMB[10][7] ) );
  FA_X1 \mult_20/S2_10_6  ( .A(\mult_20/ab[10][6] ), .B(\mult_20/CARRYB[9][6] ), .CI(\mult_20/SUMB[9][7] ), .CO(\mult_20/CARRYB[10][6] ), .S(
        \mult_20/SUMB[10][6] ) );
  FA_X1 \mult_20/S2_10_5  ( .A(\mult_20/ab[10][5] ), .B(\mult_20/CARRYB[9][5] ), .CI(\mult_20/SUMB[9][6] ), .CO(\mult_20/CARRYB[10][5] ), .S(
        \mult_20/SUMB[10][5] ) );
  FA_X1 \mult_20/S2_10_4  ( .A(\mult_20/ab[10][4] ), .B(\mult_20/CARRYB[9][4] ), .CI(\mult_20/SUMB[9][5] ), .CO(\mult_20/CARRYB[10][4] ), .S(
        \mult_20/SUMB[10][4] ) );
  FA_X1 \mult_20/S2_10_3  ( .A(\mult_20/ab[10][3] ), .B(\mult_20/CARRYB[9][3] ), .CI(\mult_20/SUMB[9][4] ), .CO(\mult_20/CARRYB[10][3] ), .S(
        \mult_20/SUMB[10][3] ) );
  FA_X1 \mult_20/S2_10_2  ( .A(\mult_20/ab[10][2] ), .B(\mult_20/CARRYB[9][2] ), .CI(\mult_20/SUMB[9][3] ), .CO(\mult_20/CARRYB[10][2] ), .S(
        \mult_20/SUMB[10][2] ) );
  FA_X1 \mult_20/S2_10_1  ( .A(\mult_20/ab[10][1] ), .B(\mult_20/CARRYB[9][1] ), .CI(\mult_20/SUMB[9][2] ), .CO(\mult_20/CARRYB[10][1] ), .S(
        \mult_20/SUMB[10][1] ) );
  FA_X1 \mult_20/S1_10_0  ( .A(\mult_20/ab[10][0] ), .B(\mult_20/CARRYB[9][0] ), .CI(\mult_20/SUMB[9][1] ), .CO(\mult_20/CARRYB[10][0] ), .S(N74) );
  FA_X1 \mult_20/S3_11_30  ( .A(\mult_20/ab[11][30] ), .B(
        \mult_20/CARRYB[10][30] ), .CI(\mult_20/ab[10][31] ), .CO(
        \mult_20/CARRYB[11][30] ), .S(\mult_20/SUMB[11][30] ) );
  FA_X1 \mult_20/S2_11_29  ( .A(\mult_20/ab[11][29] ), .B(
        \mult_20/CARRYB[10][29] ), .CI(\mult_20/SUMB[10][30] ), .CO(
        \mult_20/CARRYB[11][29] ), .S(\mult_20/SUMB[11][29] ) );
  FA_X1 \mult_20/S2_11_28  ( .A(\mult_20/ab[11][28] ), .B(
        \mult_20/CARRYB[10][28] ), .CI(\mult_20/SUMB[10][29] ), .CO(
        \mult_20/CARRYB[11][28] ), .S(\mult_20/SUMB[11][28] ) );
  FA_X1 \mult_20/S2_11_27  ( .A(\mult_20/ab[11][27] ), .B(
        \mult_20/CARRYB[10][27] ), .CI(\mult_20/SUMB[10][28] ), .CO(
        \mult_20/CARRYB[11][27] ), .S(\mult_20/SUMB[11][27] ) );
  FA_X1 \mult_20/S2_11_26  ( .A(\mult_20/ab[11][26] ), .B(
        \mult_20/CARRYB[10][26] ), .CI(\mult_20/SUMB[10][27] ), .CO(
        \mult_20/CARRYB[11][26] ), .S(\mult_20/SUMB[11][26] ) );
  FA_X1 \mult_20/S2_11_25  ( .A(\mult_20/ab[11][25] ), .B(
        \mult_20/CARRYB[10][25] ), .CI(\mult_20/SUMB[10][26] ), .CO(
        \mult_20/CARRYB[11][25] ), .S(\mult_20/SUMB[11][25] ) );
  FA_X1 \mult_20/S2_11_24  ( .A(\mult_20/ab[11][24] ), .B(
        \mult_20/CARRYB[10][24] ), .CI(\mult_20/SUMB[10][25] ), .CO(
        \mult_20/CARRYB[11][24] ), .S(\mult_20/SUMB[11][24] ) );
  FA_X1 \mult_20/S2_11_23  ( .A(\mult_20/ab[11][23] ), .B(
        \mult_20/CARRYB[10][23] ), .CI(\mult_20/SUMB[10][24] ), .CO(
        \mult_20/CARRYB[11][23] ), .S(\mult_20/SUMB[11][23] ) );
  FA_X1 \mult_20/S2_11_22  ( .A(\mult_20/ab[11][22] ), .B(
        \mult_20/CARRYB[10][22] ), .CI(\mult_20/SUMB[10][23] ), .CO(
        \mult_20/CARRYB[11][22] ), .S(\mult_20/SUMB[11][22] ) );
  FA_X1 \mult_20/S2_11_21  ( .A(\mult_20/ab[11][21] ), .B(
        \mult_20/CARRYB[10][21] ), .CI(\mult_20/SUMB[10][22] ), .CO(
        \mult_20/CARRYB[11][21] ), .S(\mult_20/SUMB[11][21] ) );
  FA_X1 \mult_20/S2_11_20  ( .A(\mult_20/ab[11][20] ), .B(
        \mult_20/CARRYB[10][20] ), .CI(\mult_20/SUMB[10][21] ), .CO(
        \mult_20/CARRYB[11][20] ), .S(\mult_20/SUMB[11][20] ) );
  FA_X1 \mult_20/S2_11_19  ( .A(\mult_20/ab[11][19] ), .B(
        \mult_20/CARRYB[10][19] ), .CI(\mult_20/SUMB[10][20] ), .CO(
        \mult_20/CARRYB[11][19] ), .S(\mult_20/SUMB[11][19] ) );
  FA_X1 \mult_20/S2_11_18  ( .A(\mult_20/ab[11][18] ), .B(
        \mult_20/CARRYB[10][18] ), .CI(\mult_20/SUMB[10][19] ), .CO(
        \mult_20/CARRYB[11][18] ), .S(\mult_20/SUMB[11][18] ) );
  FA_X1 \mult_20/S2_11_17  ( .A(\mult_20/ab[11][17] ), .B(
        \mult_20/CARRYB[10][17] ), .CI(\mult_20/SUMB[10][18] ), .CO(
        \mult_20/CARRYB[11][17] ), .S(\mult_20/SUMB[11][17] ) );
  FA_X1 \mult_20/S2_11_16  ( .A(\mult_20/ab[11][16] ), .B(
        \mult_20/CARRYB[10][16] ), .CI(\mult_20/SUMB[10][17] ), .CO(
        \mult_20/CARRYB[11][16] ), .S(\mult_20/SUMB[11][16] ) );
  FA_X1 \mult_20/S2_11_15  ( .A(\mult_20/ab[11][15] ), .B(
        \mult_20/CARRYB[10][15] ), .CI(\mult_20/SUMB[10][16] ), .CO(
        \mult_20/CARRYB[11][15] ), .S(\mult_20/SUMB[11][15] ) );
  FA_X1 \mult_20/S2_11_14  ( .A(\mult_20/ab[11][14] ), .B(
        \mult_20/CARRYB[10][14] ), .CI(\mult_20/SUMB[10][15] ), .CO(
        \mult_20/CARRYB[11][14] ), .S(\mult_20/SUMB[11][14] ) );
  FA_X1 \mult_20/S2_11_13  ( .A(\mult_20/ab[11][13] ), .B(
        \mult_20/CARRYB[10][13] ), .CI(\mult_20/SUMB[10][14] ), .CO(
        \mult_20/CARRYB[11][13] ), .S(\mult_20/SUMB[11][13] ) );
  FA_X1 \mult_20/S2_11_12  ( .A(\mult_20/ab[11][12] ), .B(
        \mult_20/CARRYB[10][12] ), .CI(\mult_20/SUMB[10][13] ), .CO(
        \mult_20/CARRYB[11][12] ), .S(\mult_20/SUMB[11][12] ) );
  FA_X1 \mult_20/S2_11_11  ( .A(\mult_20/ab[11][11] ), .B(
        \mult_20/CARRYB[10][11] ), .CI(\mult_20/SUMB[10][12] ), .CO(
        \mult_20/CARRYB[11][11] ), .S(\mult_20/SUMB[11][11] ) );
  FA_X1 \mult_20/S2_11_10  ( .A(\mult_20/ab[11][10] ), .B(
        \mult_20/CARRYB[10][10] ), .CI(\mult_20/SUMB[10][11] ), .CO(
        \mult_20/CARRYB[11][10] ), .S(\mult_20/SUMB[11][10] ) );
  FA_X1 \mult_20/S2_11_9  ( .A(\mult_20/ab[11][9] ), .B(
        \mult_20/CARRYB[10][9] ), .CI(\mult_20/SUMB[10][10] ), .CO(
        \mult_20/CARRYB[11][9] ), .S(\mult_20/SUMB[11][9] ) );
  FA_X1 \mult_20/S2_11_8  ( .A(\mult_20/ab[11][8] ), .B(
        \mult_20/CARRYB[10][8] ), .CI(\mult_20/SUMB[10][9] ), .CO(
        \mult_20/CARRYB[11][8] ), .S(\mult_20/SUMB[11][8] ) );
  FA_X1 \mult_20/S2_11_7  ( .A(\mult_20/ab[11][7] ), .B(
        \mult_20/CARRYB[10][7] ), .CI(\mult_20/SUMB[10][8] ), .CO(
        \mult_20/CARRYB[11][7] ), .S(\mult_20/SUMB[11][7] ) );
  FA_X1 \mult_20/S2_11_6  ( .A(\mult_20/ab[11][6] ), .B(
        \mult_20/CARRYB[10][6] ), .CI(\mult_20/SUMB[10][7] ), .CO(
        \mult_20/CARRYB[11][6] ), .S(\mult_20/SUMB[11][6] ) );
  FA_X1 \mult_20/S2_11_5  ( .A(\mult_20/ab[11][5] ), .B(
        \mult_20/CARRYB[10][5] ), .CI(\mult_20/SUMB[10][6] ), .CO(
        \mult_20/CARRYB[11][5] ), .S(\mult_20/SUMB[11][5] ) );
  FA_X1 \mult_20/S2_11_4  ( .A(\mult_20/ab[11][4] ), .B(
        \mult_20/CARRYB[10][4] ), .CI(\mult_20/SUMB[10][5] ), .CO(
        \mult_20/CARRYB[11][4] ), .S(\mult_20/SUMB[11][4] ) );
  FA_X1 \mult_20/S2_11_3  ( .A(\mult_20/ab[11][3] ), .B(
        \mult_20/CARRYB[10][3] ), .CI(\mult_20/SUMB[10][4] ), .CO(
        \mult_20/CARRYB[11][3] ), .S(\mult_20/SUMB[11][3] ) );
  FA_X1 \mult_20/S2_11_2  ( .A(\mult_20/ab[11][2] ), .B(
        \mult_20/CARRYB[10][2] ), .CI(\mult_20/SUMB[10][3] ), .CO(
        \mult_20/CARRYB[11][2] ), .S(\mult_20/SUMB[11][2] ) );
  FA_X1 \mult_20/S2_11_1  ( .A(\mult_20/ab[11][1] ), .B(
        \mult_20/CARRYB[10][1] ), .CI(\mult_20/SUMB[10][2] ), .CO(
        \mult_20/CARRYB[11][1] ), .S(\mult_20/SUMB[11][1] ) );
  FA_X1 \mult_20/S1_11_0  ( .A(\mult_20/ab[11][0] ), .B(
        \mult_20/CARRYB[10][0] ), .CI(\mult_20/SUMB[10][1] ), .CO(
        \mult_20/CARRYB[11][0] ), .S(N75) );
  FA_X1 \mult_20/S3_12_30  ( .A(\mult_20/ab[12][30] ), .B(
        \mult_20/CARRYB[11][30] ), .CI(\mult_20/ab[11][31] ), .CO(
        \mult_20/CARRYB[12][30] ), .S(\mult_20/SUMB[12][30] ) );
  FA_X1 \mult_20/S2_12_29  ( .A(\mult_20/ab[12][29] ), .B(
        \mult_20/CARRYB[11][29] ), .CI(\mult_20/SUMB[11][30] ), .CO(
        \mult_20/CARRYB[12][29] ), .S(\mult_20/SUMB[12][29] ) );
  FA_X1 \mult_20/S2_12_28  ( .A(\mult_20/ab[12][28] ), .B(
        \mult_20/CARRYB[11][28] ), .CI(\mult_20/SUMB[11][29] ), .CO(
        \mult_20/CARRYB[12][28] ), .S(\mult_20/SUMB[12][28] ) );
  FA_X1 \mult_20/S2_12_27  ( .A(\mult_20/ab[12][27] ), .B(
        \mult_20/CARRYB[11][27] ), .CI(\mult_20/SUMB[11][28] ), .CO(
        \mult_20/CARRYB[12][27] ), .S(\mult_20/SUMB[12][27] ) );
  FA_X1 \mult_20/S2_12_26  ( .A(\mult_20/ab[12][26] ), .B(
        \mult_20/CARRYB[11][26] ), .CI(\mult_20/SUMB[11][27] ), .CO(
        \mult_20/CARRYB[12][26] ), .S(\mult_20/SUMB[12][26] ) );
  FA_X1 \mult_20/S2_12_25  ( .A(\mult_20/ab[12][25] ), .B(
        \mult_20/CARRYB[11][25] ), .CI(\mult_20/SUMB[11][26] ), .CO(
        \mult_20/CARRYB[12][25] ), .S(\mult_20/SUMB[12][25] ) );
  FA_X1 \mult_20/S2_12_24  ( .A(\mult_20/ab[12][24] ), .B(
        \mult_20/CARRYB[11][24] ), .CI(\mult_20/SUMB[11][25] ), .CO(
        \mult_20/CARRYB[12][24] ), .S(\mult_20/SUMB[12][24] ) );
  FA_X1 \mult_20/S2_12_23  ( .A(\mult_20/ab[12][23] ), .B(
        \mult_20/CARRYB[11][23] ), .CI(\mult_20/SUMB[11][24] ), .CO(
        \mult_20/CARRYB[12][23] ), .S(\mult_20/SUMB[12][23] ) );
  FA_X1 \mult_20/S2_12_22  ( .A(\mult_20/ab[12][22] ), .B(
        \mult_20/CARRYB[11][22] ), .CI(\mult_20/SUMB[11][23] ), .CO(
        \mult_20/CARRYB[12][22] ), .S(\mult_20/SUMB[12][22] ) );
  FA_X1 \mult_20/S2_12_21  ( .A(\mult_20/ab[12][21] ), .B(
        \mult_20/CARRYB[11][21] ), .CI(\mult_20/SUMB[11][22] ), .CO(
        \mult_20/CARRYB[12][21] ), .S(\mult_20/SUMB[12][21] ) );
  FA_X1 \mult_20/S2_12_20  ( .A(\mult_20/ab[12][20] ), .B(
        \mult_20/CARRYB[11][20] ), .CI(\mult_20/SUMB[11][21] ), .CO(
        \mult_20/CARRYB[12][20] ), .S(\mult_20/SUMB[12][20] ) );
  FA_X1 \mult_20/S2_12_19  ( .A(\mult_20/ab[12][19] ), .B(
        \mult_20/CARRYB[11][19] ), .CI(\mult_20/SUMB[11][20] ), .CO(
        \mult_20/CARRYB[12][19] ), .S(\mult_20/SUMB[12][19] ) );
  FA_X1 \mult_20/S2_12_18  ( .A(\mult_20/ab[12][18] ), .B(
        \mult_20/CARRYB[11][18] ), .CI(\mult_20/SUMB[11][19] ), .CO(
        \mult_20/CARRYB[12][18] ), .S(\mult_20/SUMB[12][18] ) );
  FA_X1 \mult_20/S2_12_17  ( .A(\mult_20/ab[12][17] ), .B(
        \mult_20/CARRYB[11][17] ), .CI(\mult_20/SUMB[11][18] ), .CO(
        \mult_20/CARRYB[12][17] ), .S(\mult_20/SUMB[12][17] ) );
  FA_X1 \mult_20/S2_12_16  ( .A(\mult_20/ab[12][16] ), .B(
        \mult_20/CARRYB[11][16] ), .CI(\mult_20/SUMB[11][17] ), .CO(
        \mult_20/CARRYB[12][16] ), .S(\mult_20/SUMB[12][16] ) );
  FA_X1 \mult_20/S2_12_15  ( .A(\mult_20/ab[12][15] ), .B(
        \mult_20/CARRYB[11][15] ), .CI(\mult_20/SUMB[11][16] ), .CO(
        \mult_20/CARRYB[12][15] ), .S(\mult_20/SUMB[12][15] ) );
  FA_X1 \mult_20/S2_12_14  ( .A(\mult_20/ab[12][14] ), .B(
        \mult_20/CARRYB[11][14] ), .CI(\mult_20/SUMB[11][15] ), .CO(
        \mult_20/CARRYB[12][14] ), .S(\mult_20/SUMB[12][14] ) );
  FA_X1 \mult_20/S2_12_13  ( .A(\mult_20/ab[12][13] ), .B(
        \mult_20/CARRYB[11][13] ), .CI(\mult_20/SUMB[11][14] ), .CO(
        \mult_20/CARRYB[12][13] ), .S(\mult_20/SUMB[12][13] ) );
  FA_X1 \mult_20/S2_12_12  ( .A(\mult_20/ab[12][12] ), .B(
        \mult_20/CARRYB[11][12] ), .CI(\mult_20/SUMB[11][13] ), .CO(
        \mult_20/CARRYB[12][12] ), .S(\mult_20/SUMB[12][12] ) );
  FA_X1 \mult_20/S2_12_11  ( .A(\mult_20/ab[12][11] ), .B(
        \mult_20/CARRYB[11][11] ), .CI(\mult_20/SUMB[11][12] ), .CO(
        \mult_20/CARRYB[12][11] ), .S(\mult_20/SUMB[12][11] ) );
  FA_X1 \mult_20/S2_12_10  ( .A(\mult_20/ab[12][10] ), .B(
        \mult_20/CARRYB[11][10] ), .CI(\mult_20/SUMB[11][11] ), .CO(
        \mult_20/CARRYB[12][10] ), .S(\mult_20/SUMB[12][10] ) );
  FA_X1 \mult_20/S2_12_9  ( .A(\mult_20/ab[12][9] ), .B(
        \mult_20/CARRYB[11][9] ), .CI(\mult_20/SUMB[11][10] ), .CO(
        \mult_20/CARRYB[12][9] ), .S(\mult_20/SUMB[12][9] ) );
  FA_X1 \mult_20/S2_12_8  ( .A(\mult_20/ab[12][8] ), .B(
        \mult_20/CARRYB[11][8] ), .CI(\mult_20/SUMB[11][9] ), .CO(
        \mult_20/CARRYB[12][8] ), .S(\mult_20/SUMB[12][8] ) );
  FA_X1 \mult_20/S2_12_7  ( .A(\mult_20/ab[12][7] ), .B(
        \mult_20/CARRYB[11][7] ), .CI(\mult_20/SUMB[11][8] ), .CO(
        \mult_20/CARRYB[12][7] ), .S(\mult_20/SUMB[12][7] ) );
  FA_X1 \mult_20/S2_12_6  ( .A(\mult_20/ab[12][6] ), .B(
        \mult_20/CARRYB[11][6] ), .CI(\mult_20/SUMB[11][7] ), .CO(
        \mult_20/CARRYB[12][6] ), .S(\mult_20/SUMB[12][6] ) );
  FA_X1 \mult_20/S2_12_5  ( .A(\mult_20/ab[12][5] ), .B(
        \mult_20/CARRYB[11][5] ), .CI(\mult_20/SUMB[11][6] ), .CO(
        \mult_20/CARRYB[12][5] ), .S(\mult_20/SUMB[12][5] ) );
  FA_X1 \mult_20/S2_12_4  ( .A(\mult_20/ab[12][4] ), .B(
        \mult_20/CARRYB[11][4] ), .CI(\mult_20/SUMB[11][5] ), .CO(
        \mult_20/CARRYB[12][4] ), .S(\mult_20/SUMB[12][4] ) );
  FA_X1 \mult_20/S2_12_3  ( .A(\mult_20/ab[12][3] ), .B(
        \mult_20/CARRYB[11][3] ), .CI(\mult_20/SUMB[11][4] ), .CO(
        \mult_20/CARRYB[12][3] ), .S(\mult_20/SUMB[12][3] ) );
  FA_X1 \mult_20/S2_12_2  ( .A(\mult_20/ab[12][2] ), .B(
        \mult_20/CARRYB[11][2] ), .CI(\mult_20/SUMB[11][3] ), .CO(
        \mult_20/CARRYB[12][2] ), .S(\mult_20/SUMB[12][2] ) );
  FA_X1 \mult_20/S2_12_1  ( .A(\mult_20/ab[12][1] ), .B(
        \mult_20/CARRYB[11][1] ), .CI(\mult_20/SUMB[11][2] ), .CO(
        \mult_20/CARRYB[12][1] ), .S(\mult_20/SUMB[12][1] ) );
  FA_X1 \mult_20/S1_12_0  ( .A(\mult_20/ab[12][0] ), .B(
        \mult_20/CARRYB[11][0] ), .CI(\mult_20/SUMB[11][1] ), .CO(
        \mult_20/CARRYB[12][0] ), .S(N76) );
  FA_X1 \mult_20/S3_13_30  ( .A(\mult_20/ab[13][30] ), .B(
        \mult_20/CARRYB[12][30] ), .CI(\mult_20/ab[12][31] ), .CO(
        \mult_20/CARRYB[13][30] ), .S(\mult_20/SUMB[13][30] ) );
  FA_X1 \mult_20/S2_13_29  ( .A(\mult_20/ab[13][29] ), .B(
        \mult_20/CARRYB[12][29] ), .CI(\mult_20/SUMB[12][30] ), .CO(
        \mult_20/CARRYB[13][29] ), .S(\mult_20/SUMB[13][29] ) );
  FA_X1 \mult_20/S2_13_28  ( .A(\mult_20/ab[13][28] ), .B(
        \mult_20/CARRYB[12][28] ), .CI(\mult_20/SUMB[12][29] ), .CO(
        \mult_20/CARRYB[13][28] ), .S(\mult_20/SUMB[13][28] ) );
  FA_X1 \mult_20/S2_13_27  ( .A(\mult_20/ab[13][27] ), .B(
        \mult_20/CARRYB[12][27] ), .CI(\mult_20/SUMB[12][28] ), .CO(
        \mult_20/CARRYB[13][27] ), .S(\mult_20/SUMB[13][27] ) );
  FA_X1 \mult_20/S2_13_26  ( .A(\mult_20/ab[13][26] ), .B(
        \mult_20/CARRYB[12][26] ), .CI(\mult_20/SUMB[12][27] ), .CO(
        \mult_20/CARRYB[13][26] ), .S(\mult_20/SUMB[13][26] ) );
  FA_X1 \mult_20/S2_13_25  ( .A(\mult_20/ab[13][25] ), .B(
        \mult_20/CARRYB[12][25] ), .CI(\mult_20/SUMB[12][26] ), .CO(
        \mult_20/CARRYB[13][25] ), .S(\mult_20/SUMB[13][25] ) );
  FA_X1 \mult_20/S2_13_24  ( .A(\mult_20/ab[13][24] ), .B(
        \mult_20/CARRYB[12][24] ), .CI(\mult_20/SUMB[12][25] ), .CO(
        \mult_20/CARRYB[13][24] ), .S(\mult_20/SUMB[13][24] ) );
  FA_X1 \mult_20/S2_13_23  ( .A(\mult_20/ab[13][23] ), .B(
        \mult_20/CARRYB[12][23] ), .CI(\mult_20/SUMB[12][24] ), .CO(
        \mult_20/CARRYB[13][23] ), .S(\mult_20/SUMB[13][23] ) );
  FA_X1 \mult_20/S2_13_22  ( .A(\mult_20/ab[13][22] ), .B(
        \mult_20/CARRYB[12][22] ), .CI(\mult_20/SUMB[12][23] ), .CO(
        \mult_20/CARRYB[13][22] ), .S(\mult_20/SUMB[13][22] ) );
  FA_X1 \mult_20/S2_13_21  ( .A(\mult_20/ab[13][21] ), .B(
        \mult_20/CARRYB[12][21] ), .CI(\mult_20/SUMB[12][22] ), .CO(
        \mult_20/CARRYB[13][21] ), .S(\mult_20/SUMB[13][21] ) );
  FA_X1 \mult_20/S2_13_20  ( .A(\mult_20/ab[13][20] ), .B(
        \mult_20/CARRYB[12][20] ), .CI(\mult_20/SUMB[12][21] ), .CO(
        \mult_20/CARRYB[13][20] ), .S(\mult_20/SUMB[13][20] ) );
  FA_X1 \mult_20/S2_13_19  ( .A(\mult_20/ab[13][19] ), .B(
        \mult_20/CARRYB[12][19] ), .CI(\mult_20/SUMB[12][20] ), .CO(
        \mult_20/CARRYB[13][19] ), .S(\mult_20/SUMB[13][19] ) );
  FA_X1 \mult_20/S2_13_18  ( .A(\mult_20/ab[13][18] ), .B(
        \mult_20/CARRYB[12][18] ), .CI(\mult_20/SUMB[12][19] ), .CO(
        \mult_20/CARRYB[13][18] ), .S(\mult_20/SUMB[13][18] ) );
  FA_X1 \mult_20/S2_13_17  ( .A(\mult_20/ab[13][17] ), .B(
        \mult_20/CARRYB[12][17] ), .CI(\mult_20/SUMB[12][18] ), .CO(
        \mult_20/CARRYB[13][17] ), .S(\mult_20/SUMB[13][17] ) );
  FA_X1 \mult_20/S2_13_16  ( .A(\mult_20/ab[13][16] ), .B(
        \mult_20/CARRYB[12][16] ), .CI(\mult_20/SUMB[12][17] ), .CO(
        \mult_20/CARRYB[13][16] ), .S(\mult_20/SUMB[13][16] ) );
  FA_X1 \mult_20/S2_13_15  ( .A(\mult_20/ab[13][15] ), .B(
        \mult_20/CARRYB[12][15] ), .CI(\mult_20/SUMB[12][16] ), .CO(
        \mult_20/CARRYB[13][15] ), .S(\mult_20/SUMB[13][15] ) );
  FA_X1 \mult_20/S2_13_14  ( .A(\mult_20/ab[13][14] ), .B(
        \mult_20/CARRYB[12][14] ), .CI(\mult_20/SUMB[12][15] ), .CO(
        \mult_20/CARRYB[13][14] ), .S(\mult_20/SUMB[13][14] ) );
  FA_X1 \mult_20/S2_13_13  ( .A(\mult_20/ab[13][13] ), .B(
        \mult_20/CARRYB[12][13] ), .CI(\mult_20/SUMB[12][14] ), .CO(
        \mult_20/CARRYB[13][13] ), .S(\mult_20/SUMB[13][13] ) );
  FA_X1 \mult_20/S2_13_12  ( .A(\mult_20/ab[13][12] ), .B(
        \mult_20/CARRYB[12][12] ), .CI(\mult_20/SUMB[12][13] ), .CO(
        \mult_20/CARRYB[13][12] ), .S(\mult_20/SUMB[13][12] ) );
  FA_X1 \mult_20/S2_13_11  ( .A(\mult_20/ab[13][11] ), .B(
        \mult_20/CARRYB[12][11] ), .CI(\mult_20/SUMB[12][12] ), .CO(
        \mult_20/CARRYB[13][11] ), .S(\mult_20/SUMB[13][11] ) );
  FA_X1 \mult_20/S2_13_10  ( .A(\mult_20/ab[13][10] ), .B(
        \mult_20/CARRYB[12][10] ), .CI(\mult_20/SUMB[12][11] ), .CO(
        \mult_20/CARRYB[13][10] ), .S(\mult_20/SUMB[13][10] ) );
  FA_X1 \mult_20/S2_13_9  ( .A(\mult_20/ab[13][9] ), .B(
        \mult_20/CARRYB[12][9] ), .CI(\mult_20/SUMB[12][10] ), .CO(
        \mult_20/CARRYB[13][9] ), .S(\mult_20/SUMB[13][9] ) );
  FA_X1 \mult_20/S2_13_8  ( .A(\mult_20/ab[13][8] ), .B(
        \mult_20/CARRYB[12][8] ), .CI(\mult_20/SUMB[12][9] ), .CO(
        \mult_20/CARRYB[13][8] ), .S(\mult_20/SUMB[13][8] ) );
  FA_X1 \mult_20/S2_13_7  ( .A(\mult_20/ab[13][7] ), .B(
        \mult_20/CARRYB[12][7] ), .CI(\mult_20/SUMB[12][8] ), .CO(
        \mult_20/CARRYB[13][7] ), .S(\mult_20/SUMB[13][7] ) );
  FA_X1 \mult_20/S2_13_6  ( .A(\mult_20/ab[13][6] ), .B(
        \mult_20/CARRYB[12][6] ), .CI(\mult_20/SUMB[12][7] ), .CO(
        \mult_20/CARRYB[13][6] ), .S(\mult_20/SUMB[13][6] ) );
  FA_X1 \mult_20/S2_13_5  ( .A(\mult_20/ab[13][5] ), .B(
        \mult_20/CARRYB[12][5] ), .CI(\mult_20/SUMB[12][6] ), .CO(
        \mult_20/CARRYB[13][5] ), .S(\mult_20/SUMB[13][5] ) );
  FA_X1 \mult_20/S2_13_4  ( .A(\mult_20/ab[13][4] ), .B(
        \mult_20/CARRYB[12][4] ), .CI(\mult_20/SUMB[12][5] ), .CO(
        \mult_20/CARRYB[13][4] ), .S(\mult_20/SUMB[13][4] ) );
  FA_X1 \mult_20/S2_13_3  ( .A(\mult_20/ab[13][3] ), .B(
        \mult_20/CARRYB[12][3] ), .CI(\mult_20/SUMB[12][4] ), .CO(
        \mult_20/CARRYB[13][3] ), .S(\mult_20/SUMB[13][3] ) );
  FA_X1 \mult_20/S2_13_2  ( .A(\mult_20/ab[13][2] ), .B(
        \mult_20/CARRYB[12][2] ), .CI(\mult_20/SUMB[12][3] ), .CO(
        \mult_20/CARRYB[13][2] ), .S(\mult_20/SUMB[13][2] ) );
  FA_X1 \mult_20/S2_13_1  ( .A(\mult_20/ab[13][1] ), .B(
        \mult_20/CARRYB[12][1] ), .CI(\mult_20/SUMB[12][2] ), .CO(
        \mult_20/CARRYB[13][1] ), .S(\mult_20/SUMB[13][1] ) );
  FA_X1 \mult_20/S1_13_0  ( .A(\mult_20/ab[13][0] ), .B(
        \mult_20/CARRYB[12][0] ), .CI(\mult_20/SUMB[12][1] ), .CO(
        \mult_20/CARRYB[13][0] ), .S(N77) );
  FA_X1 \mult_20/S3_14_30  ( .A(\mult_20/ab[14][30] ), .B(
        \mult_20/CARRYB[13][30] ), .CI(\mult_20/ab[13][31] ), .CO(
        \mult_20/CARRYB[14][30] ), .S(\mult_20/SUMB[14][30] ) );
  FA_X1 \mult_20/S2_14_29  ( .A(\mult_20/ab[14][29] ), .B(
        \mult_20/CARRYB[13][29] ), .CI(\mult_20/SUMB[13][30] ), .CO(
        \mult_20/CARRYB[14][29] ), .S(\mult_20/SUMB[14][29] ) );
  FA_X1 \mult_20/S2_14_28  ( .A(\mult_20/ab[14][28] ), .B(
        \mult_20/CARRYB[13][28] ), .CI(\mult_20/SUMB[13][29] ), .CO(
        \mult_20/CARRYB[14][28] ), .S(\mult_20/SUMB[14][28] ) );
  FA_X1 \mult_20/S2_14_27  ( .A(\mult_20/ab[14][27] ), .B(
        \mult_20/CARRYB[13][27] ), .CI(\mult_20/SUMB[13][28] ), .CO(
        \mult_20/CARRYB[14][27] ), .S(\mult_20/SUMB[14][27] ) );
  FA_X1 \mult_20/S2_14_26  ( .A(\mult_20/ab[14][26] ), .B(
        \mult_20/CARRYB[13][26] ), .CI(\mult_20/SUMB[13][27] ), .CO(
        \mult_20/CARRYB[14][26] ), .S(\mult_20/SUMB[14][26] ) );
  FA_X1 \mult_20/S2_14_25  ( .A(\mult_20/ab[14][25] ), .B(
        \mult_20/CARRYB[13][25] ), .CI(\mult_20/SUMB[13][26] ), .CO(
        \mult_20/CARRYB[14][25] ), .S(\mult_20/SUMB[14][25] ) );
  FA_X1 \mult_20/S2_14_24  ( .A(\mult_20/ab[14][24] ), .B(
        \mult_20/CARRYB[13][24] ), .CI(\mult_20/SUMB[13][25] ), .CO(
        \mult_20/CARRYB[14][24] ), .S(\mult_20/SUMB[14][24] ) );
  FA_X1 \mult_20/S2_14_23  ( .A(\mult_20/ab[14][23] ), .B(
        \mult_20/CARRYB[13][23] ), .CI(\mult_20/SUMB[13][24] ), .CO(
        \mult_20/CARRYB[14][23] ), .S(\mult_20/SUMB[14][23] ) );
  FA_X1 \mult_20/S2_14_22  ( .A(\mult_20/ab[14][22] ), .B(
        \mult_20/CARRYB[13][22] ), .CI(\mult_20/SUMB[13][23] ), .CO(
        \mult_20/CARRYB[14][22] ), .S(\mult_20/SUMB[14][22] ) );
  FA_X1 \mult_20/S2_14_21  ( .A(\mult_20/ab[14][21] ), .B(
        \mult_20/CARRYB[13][21] ), .CI(\mult_20/SUMB[13][22] ), .CO(
        \mult_20/CARRYB[14][21] ), .S(\mult_20/SUMB[14][21] ) );
  FA_X1 \mult_20/S2_14_20  ( .A(\mult_20/ab[14][20] ), .B(
        \mult_20/CARRYB[13][20] ), .CI(\mult_20/SUMB[13][21] ), .CO(
        \mult_20/CARRYB[14][20] ), .S(\mult_20/SUMB[14][20] ) );
  FA_X1 \mult_20/S2_14_19  ( .A(\mult_20/ab[14][19] ), .B(
        \mult_20/CARRYB[13][19] ), .CI(\mult_20/SUMB[13][20] ), .CO(
        \mult_20/CARRYB[14][19] ), .S(\mult_20/SUMB[14][19] ) );
  FA_X1 \mult_20/S2_14_18  ( .A(\mult_20/ab[14][18] ), .B(
        \mult_20/CARRYB[13][18] ), .CI(\mult_20/SUMB[13][19] ), .CO(
        \mult_20/CARRYB[14][18] ), .S(\mult_20/SUMB[14][18] ) );
  FA_X1 \mult_20/S2_14_17  ( .A(\mult_20/ab[14][17] ), .B(
        \mult_20/CARRYB[13][17] ), .CI(\mult_20/SUMB[13][18] ), .CO(
        \mult_20/CARRYB[14][17] ), .S(\mult_20/SUMB[14][17] ) );
  FA_X1 \mult_20/S2_14_16  ( .A(\mult_20/ab[14][16] ), .B(
        \mult_20/CARRYB[13][16] ), .CI(\mult_20/SUMB[13][17] ), .CO(
        \mult_20/CARRYB[14][16] ), .S(\mult_20/SUMB[14][16] ) );
  FA_X1 \mult_20/S2_14_15  ( .A(\mult_20/ab[14][15] ), .B(
        \mult_20/CARRYB[13][15] ), .CI(\mult_20/SUMB[13][16] ), .CO(
        \mult_20/CARRYB[14][15] ), .S(\mult_20/SUMB[14][15] ) );
  FA_X1 \mult_20/S2_14_14  ( .A(\mult_20/ab[14][14] ), .B(
        \mult_20/CARRYB[13][14] ), .CI(\mult_20/SUMB[13][15] ), .CO(
        \mult_20/CARRYB[14][14] ), .S(\mult_20/SUMB[14][14] ) );
  FA_X1 \mult_20/S2_14_13  ( .A(\mult_20/ab[14][13] ), .B(
        \mult_20/CARRYB[13][13] ), .CI(\mult_20/SUMB[13][14] ), .CO(
        \mult_20/CARRYB[14][13] ), .S(\mult_20/SUMB[14][13] ) );
  FA_X1 \mult_20/S2_14_12  ( .A(\mult_20/ab[14][12] ), .B(
        \mult_20/CARRYB[13][12] ), .CI(\mult_20/SUMB[13][13] ), .CO(
        \mult_20/CARRYB[14][12] ), .S(\mult_20/SUMB[14][12] ) );
  FA_X1 \mult_20/S2_14_11  ( .A(\mult_20/ab[14][11] ), .B(
        \mult_20/CARRYB[13][11] ), .CI(\mult_20/SUMB[13][12] ), .CO(
        \mult_20/CARRYB[14][11] ), .S(\mult_20/SUMB[14][11] ) );
  FA_X1 \mult_20/S2_14_10  ( .A(\mult_20/ab[14][10] ), .B(
        \mult_20/CARRYB[13][10] ), .CI(\mult_20/SUMB[13][11] ), .CO(
        \mult_20/CARRYB[14][10] ), .S(\mult_20/SUMB[14][10] ) );
  FA_X1 \mult_20/S2_14_9  ( .A(\mult_20/ab[14][9] ), .B(
        \mult_20/CARRYB[13][9] ), .CI(\mult_20/SUMB[13][10] ), .CO(
        \mult_20/CARRYB[14][9] ), .S(\mult_20/SUMB[14][9] ) );
  FA_X1 \mult_20/S2_14_8  ( .A(\mult_20/ab[14][8] ), .B(
        \mult_20/CARRYB[13][8] ), .CI(\mult_20/SUMB[13][9] ), .CO(
        \mult_20/CARRYB[14][8] ), .S(\mult_20/SUMB[14][8] ) );
  FA_X1 \mult_20/S2_14_7  ( .A(\mult_20/ab[14][7] ), .B(
        \mult_20/CARRYB[13][7] ), .CI(\mult_20/SUMB[13][8] ), .CO(
        \mult_20/CARRYB[14][7] ), .S(\mult_20/SUMB[14][7] ) );
  FA_X1 \mult_20/S2_14_6  ( .A(\mult_20/ab[14][6] ), .B(
        \mult_20/CARRYB[13][6] ), .CI(\mult_20/SUMB[13][7] ), .CO(
        \mult_20/CARRYB[14][6] ), .S(\mult_20/SUMB[14][6] ) );
  FA_X1 \mult_20/S2_14_5  ( .A(\mult_20/ab[14][5] ), .B(
        \mult_20/CARRYB[13][5] ), .CI(\mult_20/SUMB[13][6] ), .CO(
        \mult_20/CARRYB[14][5] ), .S(\mult_20/SUMB[14][5] ) );
  FA_X1 \mult_20/S2_14_4  ( .A(\mult_20/ab[14][4] ), .B(
        \mult_20/CARRYB[13][4] ), .CI(\mult_20/SUMB[13][5] ), .CO(
        \mult_20/CARRYB[14][4] ), .S(\mult_20/SUMB[14][4] ) );
  FA_X1 \mult_20/S2_14_3  ( .A(\mult_20/ab[14][3] ), .B(
        \mult_20/CARRYB[13][3] ), .CI(\mult_20/SUMB[13][4] ), .CO(
        \mult_20/CARRYB[14][3] ), .S(\mult_20/SUMB[14][3] ) );
  FA_X1 \mult_20/S2_14_2  ( .A(\mult_20/ab[14][2] ), .B(
        \mult_20/CARRYB[13][2] ), .CI(\mult_20/SUMB[13][3] ), .CO(
        \mult_20/CARRYB[14][2] ), .S(\mult_20/SUMB[14][2] ) );
  FA_X1 \mult_20/S2_14_1  ( .A(\mult_20/ab[14][1] ), .B(
        \mult_20/CARRYB[13][1] ), .CI(\mult_20/SUMB[13][2] ), .CO(
        \mult_20/CARRYB[14][1] ), .S(\mult_20/SUMB[14][1] ) );
  FA_X1 \mult_20/S1_14_0  ( .A(\mult_20/ab[14][0] ), .B(
        \mult_20/CARRYB[13][0] ), .CI(\mult_20/SUMB[13][1] ), .CO(
        \mult_20/CARRYB[14][0] ), .S(N78) );
  FA_X1 \mult_20/S3_15_30  ( .A(\mult_20/ab[15][30] ), .B(
        \mult_20/CARRYB[14][30] ), .CI(\mult_20/ab[14][31] ), .CO(
        \mult_20/CARRYB[15][30] ), .S(\mult_20/SUMB[15][30] ) );
  FA_X1 \mult_20/S2_15_29  ( .A(\mult_20/ab[15][29] ), .B(
        \mult_20/CARRYB[14][29] ), .CI(\mult_20/SUMB[14][30] ), .CO(
        \mult_20/CARRYB[15][29] ), .S(\mult_20/SUMB[15][29] ) );
  FA_X1 \mult_20/S2_15_28  ( .A(\mult_20/ab[15][28] ), .B(
        \mult_20/CARRYB[14][28] ), .CI(\mult_20/SUMB[14][29] ), .CO(
        \mult_20/CARRYB[15][28] ), .S(\mult_20/SUMB[15][28] ) );
  FA_X1 \mult_20/S2_15_27  ( .A(\mult_20/ab[15][27] ), .B(
        \mult_20/CARRYB[14][27] ), .CI(\mult_20/SUMB[14][28] ), .CO(
        \mult_20/CARRYB[15][27] ), .S(\mult_20/SUMB[15][27] ) );
  FA_X1 \mult_20/S2_15_26  ( .A(\mult_20/ab[15][26] ), .B(
        \mult_20/CARRYB[14][26] ), .CI(\mult_20/SUMB[14][27] ), .CO(
        \mult_20/CARRYB[15][26] ), .S(\mult_20/SUMB[15][26] ) );
  FA_X1 \mult_20/S2_15_25  ( .A(\mult_20/ab[15][25] ), .B(
        \mult_20/CARRYB[14][25] ), .CI(\mult_20/SUMB[14][26] ), .CO(
        \mult_20/CARRYB[15][25] ), .S(\mult_20/SUMB[15][25] ) );
  FA_X1 \mult_20/S2_15_24  ( .A(\mult_20/ab[15][24] ), .B(
        \mult_20/CARRYB[14][24] ), .CI(\mult_20/SUMB[14][25] ), .CO(
        \mult_20/CARRYB[15][24] ), .S(\mult_20/SUMB[15][24] ) );
  FA_X1 \mult_20/S2_15_23  ( .A(\mult_20/ab[15][23] ), .B(
        \mult_20/CARRYB[14][23] ), .CI(\mult_20/SUMB[14][24] ), .CO(
        \mult_20/CARRYB[15][23] ), .S(\mult_20/SUMB[15][23] ) );
  FA_X1 \mult_20/S2_15_22  ( .A(\mult_20/ab[15][22] ), .B(
        \mult_20/CARRYB[14][22] ), .CI(\mult_20/SUMB[14][23] ), .CO(
        \mult_20/CARRYB[15][22] ), .S(\mult_20/SUMB[15][22] ) );
  FA_X1 \mult_20/S2_15_21  ( .A(\mult_20/ab[15][21] ), .B(
        \mult_20/CARRYB[14][21] ), .CI(\mult_20/SUMB[14][22] ), .CO(
        \mult_20/CARRYB[15][21] ), .S(\mult_20/SUMB[15][21] ) );
  FA_X1 \mult_20/S2_15_20  ( .A(\mult_20/ab[15][20] ), .B(
        \mult_20/CARRYB[14][20] ), .CI(\mult_20/SUMB[14][21] ), .CO(
        \mult_20/CARRYB[15][20] ), .S(\mult_20/SUMB[15][20] ) );
  FA_X1 \mult_20/S2_15_19  ( .A(\mult_20/ab[15][19] ), .B(
        \mult_20/CARRYB[14][19] ), .CI(\mult_20/SUMB[14][20] ), .CO(
        \mult_20/CARRYB[15][19] ), .S(\mult_20/SUMB[15][19] ) );
  FA_X1 \mult_20/S2_15_18  ( .A(\mult_20/ab[15][18] ), .B(
        \mult_20/CARRYB[14][18] ), .CI(\mult_20/SUMB[14][19] ), .CO(
        \mult_20/CARRYB[15][18] ), .S(\mult_20/SUMB[15][18] ) );
  FA_X1 \mult_20/S2_15_17  ( .A(\mult_20/ab[15][17] ), .B(
        \mult_20/CARRYB[14][17] ), .CI(\mult_20/SUMB[14][18] ), .CO(
        \mult_20/CARRYB[15][17] ), .S(\mult_20/SUMB[15][17] ) );
  FA_X1 \mult_20/S2_15_16  ( .A(\mult_20/ab[15][16] ), .B(
        \mult_20/CARRYB[14][16] ), .CI(\mult_20/SUMB[14][17] ), .CO(
        \mult_20/CARRYB[15][16] ), .S(\mult_20/SUMB[15][16] ) );
  FA_X1 \mult_20/S2_15_15  ( .A(\mult_20/ab[15][15] ), .B(
        \mult_20/CARRYB[14][15] ), .CI(\mult_20/SUMB[14][16] ), .CO(
        \mult_20/CARRYB[15][15] ), .S(\mult_20/SUMB[15][15] ) );
  FA_X1 \mult_20/S2_15_14  ( .A(\mult_20/ab[15][14] ), .B(
        \mult_20/CARRYB[14][14] ), .CI(\mult_20/SUMB[14][15] ), .CO(
        \mult_20/CARRYB[15][14] ), .S(\mult_20/SUMB[15][14] ) );
  FA_X1 \mult_20/S2_15_13  ( .A(\mult_20/ab[15][13] ), .B(
        \mult_20/CARRYB[14][13] ), .CI(\mult_20/SUMB[14][14] ), .CO(
        \mult_20/CARRYB[15][13] ), .S(\mult_20/SUMB[15][13] ) );
  FA_X1 \mult_20/S2_15_12  ( .A(\mult_20/ab[15][12] ), .B(
        \mult_20/CARRYB[14][12] ), .CI(\mult_20/SUMB[14][13] ), .CO(
        \mult_20/CARRYB[15][12] ), .S(\mult_20/SUMB[15][12] ) );
  FA_X1 \mult_20/S2_15_11  ( .A(\mult_20/ab[15][11] ), .B(
        \mult_20/CARRYB[14][11] ), .CI(\mult_20/SUMB[14][12] ), .CO(
        \mult_20/CARRYB[15][11] ), .S(\mult_20/SUMB[15][11] ) );
  FA_X1 \mult_20/S2_15_10  ( .A(\mult_20/ab[15][10] ), .B(
        \mult_20/CARRYB[14][10] ), .CI(\mult_20/SUMB[14][11] ), .CO(
        \mult_20/CARRYB[15][10] ), .S(\mult_20/SUMB[15][10] ) );
  FA_X1 \mult_20/S2_15_9  ( .A(\mult_20/ab[15][9] ), .B(
        \mult_20/CARRYB[14][9] ), .CI(\mult_20/SUMB[14][10] ), .CO(
        \mult_20/CARRYB[15][9] ), .S(\mult_20/SUMB[15][9] ) );
  FA_X1 \mult_20/S2_15_8  ( .A(\mult_20/ab[15][8] ), .B(
        \mult_20/CARRYB[14][8] ), .CI(\mult_20/SUMB[14][9] ), .CO(
        \mult_20/CARRYB[15][8] ), .S(\mult_20/SUMB[15][8] ) );
  FA_X1 \mult_20/S2_15_7  ( .A(\mult_20/ab[15][7] ), .B(
        \mult_20/CARRYB[14][7] ), .CI(\mult_20/SUMB[14][8] ), .CO(
        \mult_20/CARRYB[15][7] ), .S(\mult_20/SUMB[15][7] ) );
  FA_X1 \mult_20/S2_15_6  ( .A(\mult_20/ab[15][6] ), .B(
        \mult_20/CARRYB[14][6] ), .CI(\mult_20/SUMB[14][7] ), .CO(
        \mult_20/CARRYB[15][6] ), .S(\mult_20/SUMB[15][6] ) );
  FA_X1 \mult_20/S2_15_5  ( .A(\mult_20/ab[15][5] ), .B(
        \mult_20/CARRYB[14][5] ), .CI(\mult_20/SUMB[14][6] ), .CO(
        \mult_20/CARRYB[15][5] ), .S(\mult_20/SUMB[15][5] ) );
  FA_X1 \mult_20/S2_15_4  ( .A(\mult_20/ab[15][4] ), .B(
        \mult_20/CARRYB[14][4] ), .CI(\mult_20/SUMB[14][5] ), .CO(
        \mult_20/CARRYB[15][4] ), .S(\mult_20/SUMB[15][4] ) );
  FA_X1 \mult_20/S2_15_3  ( .A(\mult_20/ab[15][3] ), .B(
        \mult_20/CARRYB[14][3] ), .CI(\mult_20/SUMB[14][4] ), .CO(
        \mult_20/CARRYB[15][3] ), .S(\mult_20/SUMB[15][3] ) );
  FA_X1 \mult_20/S2_15_2  ( .A(\mult_20/ab[15][2] ), .B(
        \mult_20/CARRYB[14][2] ), .CI(\mult_20/SUMB[14][3] ), .CO(
        \mult_20/CARRYB[15][2] ), .S(\mult_20/SUMB[15][2] ) );
  FA_X1 \mult_20/S2_15_1  ( .A(\mult_20/ab[15][1] ), .B(
        \mult_20/CARRYB[14][1] ), .CI(\mult_20/SUMB[14][2] ), .CO(
        \mult_20/CARRYB[15][1] ), .S(\mult_20/SUMB[15][1] ) );
  FA_X1 \mult_20/S1_15_0  ( .A(\mult_20/ab[15][0] ), .B(
        \mult_20/CARRYB[14][0] ), .CI(\mult_20/SUMB[14][1] ), .CO(
        \mult_20/CARRYB[15][0] ), .S(N79) );
  FA_X1 \mult_20/S3_16_30  ( .A(\mult_20/ab[16][30] ), .B(
        \mult_20/CARRYB[15][30] ), .CI(\mult_20/ab[15][31] ), .CO(
        \mult_20/CARRYB[16][30] ), .S(\mult_20/SUMB[16][30] ) );
  FA_X1 \mult_20/S2_16_29  ( .A(\mult_20/ab[16][29] ), .B(
        \mult_20/CARRYB[15][29] ), .CI(\mult_20/SUMB[15][30] ), .CO(
        \mult_20/CARRYB[16][29] ), .S(\mult_20/SUMB[16][29] ) );
  FA_X1 \mult_20/S2_16_28  ( .A(\mult_20/ab[16][28] ), .B(
        \mult_20/CARRYB[15][28] ), .CI(\mult_20/SUMB[15][29] ), .CO(
        \mult_20/CARRYB[16][28] ), .S(\mult_20/SUMB[16][28] ) );
  FA_X1 \mult_20/S2_16_27  ( .A(\mult_20/ab[16][27] ), .B(
        \mult_20/CARRYB[15][27] ), .CI(\mult_20/SUMB[15][28] ), .CO(
        \mult_20/CARRYB[16][27] ), .S(\mult_20/SUMB[16][27] ) );
  FA_X1 \mult_20/S2_16_26  ( .A(\mult_20/ab[16][26] ), .B(
        \mult_20/CARRYB[15][26] ), .CI(\mult_20/SUMB[15][27] ), .CO(
        \mult_20/CARRYB[16][26] ), .S(\mult_20/SUMB[16][26] ) );
  FA_X1 \mult_20/S2_16_25  ( .A(\mult_20/ab[16][25] ), .B(
        \mult_20/CARRYB[15][25] ), .CI(\mult_20/SUMB[15][26] ), .CO(
        \mult_20/CARRYB[16][25] ), .S(\mult_20/SUMB[16][25] ) );
  FA_X1 \mult_20/S2_16_24  ( .A(\mult_20/ab[16][24] ), .B(
        \mult_20/CARRYB[15][24] ), .CI(\mult_20/SUMB[15][25] ), .CO(
        \mult_20/CARRYB[16][24] ), .S(\mult_20/SUMB[16][24] ) );
  FA_X1 \mult_20/S2_16_23  ( .A(\mult_20/ab[16][23] ), .B(
        \mult_20/CARRYB[15][23] ), .CI(\mult_20/SUMB[15][24] ), .CO(
        \mult_20/CARRYB[16][23] ), .S(\mult_20/SUMB[16][23] ) );
  FA_X1 \mult_20/S2_16_22  ( .A(\mult_20/ab[16][22] ), .B(
        \mult_20/CARRYB[15][22] ), .CI(\mult_20/SUMB[15][23] ), .CO(
        \mult_20/CARRYB[16][22] ), .S(\mult_20/SUMB[16][22] ) );
  FA_X1 \mult_20/S2_16_21  ( .A(\mult_20/ab[16][21] ), .B(
        \mult_20/CARRYB[15][21] ), .CI(\mult_20/SUMB[15][22] ), .CO(
        \mult_20/CARRYB[16][21] ), .S(\mult_20/SUMB[16][21] ) );
  FA_X1 \mult_20/S2_16_20  ( .A(\mult_20/ab[16][20] ), .B(
        \mult_20/CARRYB[15][20] ), .CI(\mult_20/SUMB[15][21] ), .CO(
        \mult_20/CARRYB[16][20] ), .S(\mult_20/SUMB[16][20] ) );
  FA_X1 \mult_20/S2_16_19  ( .A(\mult_20/ab[16][19] ), .B(
        \mult_20/CARRYB[15][19] ), .CI(\mult_20/SUMB[15][20] ), .CO(
        \mult_20/CARRYB[16][19] ), .S(\mult_20/SUMB[16][19] ) );
  FA_X1 \mult_20/S2_16_18  ( .A(\mult_20/ab[16][18] ), .B(
        \mult_20/CARRYB[15][18] ), .CI(\mult_20/SUMB[15][19] ), .CO(
        \mult_20/CARRYB[16][18] ), .S(\mult_20/SUMB[16][18] ) );
  FA_X1 \mult_20/S2_16_17  ( .A(\mult_20/ab[16][17] ), .B(
        \mult_20/CARRYB[15][17] ), .CI(\mult_20/SUMB[15][18] ), .CO(
        \mult_20/CARRYB[16][17] ), .S(\mult_20/SUMB[16][17] ) );
  FA_X1 \mult_20/S2_16_16  ( .A(\mult_20/ab[16][16] ), .B(
        \mult_20/CARRYB[15][16] ), .CI(\mult_20/SUMB[15][17] ), .CO(
        \mult_20/CARRYB[16][16] ), .S(\mult_20/SUMB[16][16] ) );
  FA_X1 \mult_20/S2_16_15  ( .A(\mult_20/ab[16][15] ), .B(
        \mult_20/CARRYB[15][15] ), .CI(\mult_20/SUMB[15][16] ), .CO(
        \mult_20/CARRYB[16][15] ), .S(\mult_20/SUMB[16][15] ) );
  FA_X1 \mult_20/S2_16_14  ( .A(\mult_20/ab[16][14] ), .B(
        \mult_20/CARRYB[15][14] ), .CI(\mult_20/SUMB[15][15] ), .CO(
        \mult_20/CARRYB[16][14] ), .S(\mult_20/SUMB[16][14] ) );
  FA_X1 \mult_20/S2_16_13  ( .A(\mult_20/ab[16][13] ), .B(
        \mult_20/CARRYB[15][13] ), .CI(\mult_20/SUMB[15][14] ), .CO(
        \mult_20/CARRYB[16][13] ), .S(\mult_20/SUMB[16][13] ) );
  FA_X1 \mult_20/S2_16_12  ( .A(\mult_20/ab[16][12] ), .B(
        \mult_20/CARRYB[15][12] ), .CI(\mult_20/SUMB[15][13] ), .CO(
        \mult_20/CARRYB[16][12] ), .S(\mult_20/SUMB[16][12] ) );
  FA_X1 \mult_20/S2_16_11  ( .A(\mult_20/ab[16][11] ), .B(
        \mult_20/CARRYB[15][11] ), .CI(\mult_20/SUMB[15][12] ), .CO(
        \mult_20/CARRYB[16][11] ), .S(\mult_20/SUMB[16][11] ) );
  FA_X1 \mult_20/S2_16_10  ( .A(\mult_20/ab[16][10] ), .B(
        \mult_20/CARRYB[15][10] ), .CI(\mult_20/SUMB[15][11] ), .CO(
        \mult_20/CARRYB[16][10] ), .S(\mult_20/SUMB[16][10] ) );
  FA_X1 \mult_20/S2_16_9  ( .A(\mult_20/ab[16][9] ), .B(
        \mult_20/CARRYB[15][9] ), .CI(\mult_20/SUMB[15][10] ), .CO(
        \mult_20/CARRYB[16][9] ), .S(\mult_20/SUMB[16][9] ) );
  FA_X1 \mult_20/S2_16_8  ( .A(\mult_20/ab[16][8] ), .B(
        \mult_20/CARRYB[15][8] ), .CI(\mult_20/SUMB[15][9] ), .CO(
        \mult_20/CARRYB[16][8] ), .S(\mult_20/SUMB[16][8] ) );
  FA_X1 \mult_20/S2_16_7  ( .A(\mult_20/ab[16][7] ), .B(
        \mult_20/CARRYB[15][7] ), .CI(\mult_20/SUMB[15][8] ), .CO(
        \mult_20/CARRYB[16][7] ), .S(\mult_20/SUMB[16][7] ) );
  FA_X1 \mult_20/S2_16_6  ( .A(\mult_20/ab[16][6] ), .B(
        \mult_20/CARRYB[15][6] ), .CI(\mult_20/SUMB[15][7] ), .CO(
        \mult_20/CARRYB[16][6] ), .S(\mult_20/SUMB[16][6] ) );
  FA_X1 \mult_20/S2_16_5  ( .A(\mult_20/ab[16][5] ), .B(
        \mult_20/CARRYB[15][5] ), .CI(\mult_20/SUMB[15][6] ), .CO(
        \mult_20/CARRYB[16][5] ), .S(\mult_20/SUMB[16][5] ) );
  FA_X1 \mult_20/S2_16_4  ( .A(\mult_20/ab[16][4] ), .B(
        \mult_20/CARRYB[15][4] ), .CI(\mult_20/SUMB[15][5] ), .CO(
        \mult_20/CARRYB[16][4] ), .S(\mult_20/SUMB[16][4] ) );
  FA_X1 \mult_20/S2_16_3  ( .A(\mult_20/ab[16][3] ), .B(
        \mult_20/CARRYB[15][3] ), .CI(\mult_20/SUMB[15][4] ), .CO(
        \mult_20/CARRYB[16][3] ), .S(\mult_20/SUMB[16][3] ) );
  FA_X1 \mult_20/S2_16_2  ( .A(\mult_20/ab[16][2] ), .B(
        \mult_20/CARRYB[15][2] ), .CI(\mult_20/SUMB[15][3] ), .CO(
        \mult_20/CARRYB[16][2] ), .S(\mult_20/SUMB[16][2] ) );
  FA_X1 \mult_20/S2_16_1  ( .A(\mult_20/ab[16][1] ), .B(
        \mult_20/CARRYB[15][1] ), .CI(\mult_20/SUMB[15][2] ), .CO(
        \mult_20/CARRYB[16][1] ), .S(\mult_20/SUMB[16][1] ) );
  FA_X1 \mult_20/S1_16_0  ( .A(\mult_20/ab[16][0] ), .B(
        \mult_20/CARRYB[15][0] ), .CI(\mult_20/SUMB[15][1] ), .CO(
        \mult_20/CARRYB[16][0] ), .S(N80) );
  FA_X1 \mult_20/S3_17_30  ( .A(\mult_20/ab[17][30] ), .B(
        \mult_20/CARRYB[16][30] ), .CI(\mult_20/ab[16][31] ), .CO(
        \mult_20/CARRYB[17][30] ), .S(\mult_20/SUMB[17][30] ) );
  FA_X1 \mult_20/S2_17_29  ( .A(\mult_20/ab[17][29] ), .B(
        \mult_20/CARRYB[16][29] ), .CI(\mult_20/SUMB[16][30] ), .CO(
        \mult_20/CARRYB[17][29] ), .S(\mult_20/SUMB[17][29] ) );
  FA_X1 \mult_20/S2_17_28  ( .A(\mult_20/ab[17][28] ), .B(
        \mult_20/CARRYB[16][28] ), .CI(\mult_20/SUMB[16][29] ), .CO(
        \mult_20/CARRYB[17][28] ), .S(\mult_20/SUMB[17][28] ) );
  FA_X1 \mult_20/S2_17_27  ( .A(\mult_20/ab[17][27] ), .B(
        \mult_20/CARRYB[16][27] ), .CI(\mult_20/SUMB[16][28] ), .CO(
        \mult_20/CARRYB[17][27] ), .S(\mult_20/SUMB[17][27] ) );
  FA_X1 \mult_20/S2_17_26  ( .A(\mult_20/ab[17][26] ), .B(
        \mult_20/CARRYB[16][26] ), .CI(\mult_20/SUMB[16][27] ), .CO(
        \mult_20/CARRYB[17][26] ), .S(\mult_20/SUMB[17][26] ) );
  FA_X1 \mult_20/S2_17_25  ( .A(\mult_20/ab[17][25] ), .B(
        \mult_20/CARRYB[16][25] ), .CI(\mult_20/SUMB[16][26] ), .CO(
        \mult_20/CARRYB[17][25] ), .S(\mult_20/SUMB[17][25] ) );
  FA_X1 \mult_20/S2_17_24  ( .A(\mult_20/ab[17][24] ), .B(
        \mult_20/CARRYB[16][24] ), .CI(\mult_20/SUMB[16][25] ), .CO(
        \mult_20/CARRYB[17][24] ), .S(\mult_20/SUMB[17][24] ) );
  FA_X1 \mult_20/S2_17_23  ( .A(\mult_20/ab[17][23] ), .B(
        \mult_20/CARRYB[16][23] ), .CI(\mult_20/SUMB[16][24] ), .CO(
        \mult_20/CARRYB[17][23] ), .S(\mult_20/SUMB[17][23] ) );
  FA_X1 \mult_20/S2_17_22  ( .A(\mult_20/ab[17][22] ), .B(
        \mult_20/CARRYB[16][22] ), .CI(\mult_20/SUMB[16][23] ), .CO(
        \mult_20/CARRYB[17][22] ), .S(\mult_20/SUMB[17][22] ) );
  FA_X1 \mult_20/S2_17_21  ( .A(\mult_20/ab[17][21] ), .B(
        \mult_20/CARRYB[16][21] ), .CI(\mult_20/SUMB[16][22] ), .CO(
        \mult_20/CARRYB[17][21] ), .S(\mult_20/SUMB[17][21] ) );
  FA_X1 \mult_20/S2_17_20  ( .A(\mult_20/ab[17][20] ), .B(
        \mult_20/CARRYB[16][20] ), .CI(\mult_20/SUMB[16][21] ), .CO(
        \mult_20/CARRYB[17][20] ), .S(\mult_20/SUMB[17][20] ) );
  FA_X1 \mult_20/S2_17_19  ( .A(\mult_20/ab[17][19] ), .B(
        \mult_20/CARRYB[16][19] ), .CI(\mult_20/SUMB[16][20] ), .CO(
        \mult_20/CARRYB[17][19] ), .S(\mult_20/SUMB[17][19] ) );
  FA_X1 \mult_20/S2_17_18  ( .A(\mult_20/ab[17][18] ), .B(
        \mult_20/CARRYB[16][18] ), .CI(\mult_20/SUMB[16][19] ), .CO(
        \mult_20/CARRYB[17][18] ), .S(\mult_20/SUMB[17][18] ) );
  FA_X1 \mult_20/S2_17_17  ( .A(\mult_20/ab[17][17] ), .B(
        \mult_20/CARRYB[16][17] ), .CI(\mult_20/SUMB[16][18] ), .CO(
        \mult_20/CARRYB[17][17] ), .S(\mult_20/SUMB[17][17] ) );
  FA_X1 \mult_20/S2_17_16  ( .A(\mult_20/ab[17][16] ), .B(
        \mult_20/CARRYB[16][16] ), .CI(\mult_20/SUMB[16][17] ), .CO(
        \mult_20/CARRYB[17][16] ), .S(\mult_20/SUMB[17][16] ) );
  FA_X1 \mult_20/S2_17_15  ( .A(\mult_20/ab[17][15] ), .B(
        \mult_20/CARRYB[16][15] ), .CI(\mult_20/SUMB[16][16] ), .CO(
        \mult_20/CARRYB[17][15] ), .S(\mult_20/SUMB[17][15] ) );
  FA_X1 \mult_20/S2_17_14  ( .A(\mult_20/ab[17][14] ), .B(
        \mult_20/CARRYB[16][14] ), .CI(\mult_20/SUMB[16][15] ), .CO(
        \mult_20/CARRYB[17][14] ), .S(\mult_20/SUMB[17][14] ) );
  FA_X1 \mult_20/S2_17_13  ( .A(\mult_20/ab[17][13] ), .B(
        \mult_20/CARRYB[16][13] ), .CI(\mult_20/SUMB[16][14] ), .CO(
        \mult_20/CARRYB[17][13] ), .S(\mult_20/SUMB[17][13] ) );
  FA_X1 \mult_20/S2_17_12  ( .A(\mult_20/ab[17][12] ), .B(
        \mult_20/CARRYB[16][12] ), .CI(\mult_20/SUMB[16][13] ), .CO(
        \mult_20/CARRYB[17][12] ), .S(\mult_20/SUMB[17][12] ) );
  FA_X1 \mult_20/S2_17_11  ( .A(\mult_20/ab[17][11] ), .B(
        \mult_20/CARRYB[16][11] ), .CI(\mult_20/SUMB[16][12] ), .CO(
        \mult_20/CARRYB[17][11] ), .S(\mult_20/SUMB[17][11] ) );
  FA_X1 \mult_20/S2_17_10  ( .A(\mult_20/ab[17][10] ), .B(
        \mult_20/CARRYB[16][10] ), .CI(\mult_20/SUMB[16][11] ), .CO(
        \mult_20/CARRYB[17][10] ), .S(\mult_20/SUMB[17][10] ) );
  FA_X1 \mult_20/S2_17_9  ( .A(\mult_20/ab[17][9] ), .B(
        \mult_20/CARRYB[16][9] ), .CI(\mult_20/SUMB[16][10] ), .CO(
        \mult_20/CARRYB[17][9] ), .S(\mult_20/SUMB[17][9] ) );
  FA_X1 \mult_20/S2_17_8  ( .A(\mult_20/ab[17][8] ), .B(
        \mult_20/CARRYB[16][8] ), .CI(\mult_20/SUMB[16][9] ), .CO(
        \mult_20/CARRYB[17][8] ), .S(\mult_20/SUMB[17][8] ) );
  FA_X1 \mult_20/S2_17_7  ( .A(\mult_20/ab[17][7] ), .B(
        \mult_20/CARRYB[16][7] ), .CI(\mult_20/SUMB[16][8] ), .CO(
        \mult_20/CARRYB[17][7] ), .S(\mult_20/SUMB[17][7] ) );
  FA_X1 \mult_20/S2_17_6  ( .A(\mult_20/ab[17][6] ), .B(
        \mult_20/CARRYB[16][6] ), .CI(\mult_20/SUMB[16][7] ), .CO(
        \mult_20/CARRYB[17][6] ), .S(\mult_20/SUMB[17][6] ) );
  FA_X1 \mult_20/S2_17_5  ( .A(\mult_20/ab[17][5] ), .B(
        \mult_20/CARRYB[16][5] ), .CI(\mult_20/SUMB[16][6] ), .CO(
        \mult_20/CARRYB[17][5] ), .S(\mult_20/SUMB[17][5] ) );
  FA_X1 \mult_20/S2_17_4  ( .A(\mult_20/ab[17][4] ), .B(
        \mult_20/CARRYB[16][4] ), .CI(\mult_20/SUMB[16][5] ), .CO(
        \mult_20/CARRYB[17][4] ), .S(\mult_20/SUMB[17][4] ) );
  FA_X1 \mult_20/S2_17_3  ( .A(\mult_20/ab[17][3] ), .B(
        \mult_20/CARRYB[16][3] ), .CI(\mult_20/SUMB[16][4] ), .CO(
        \mult_20/CARRYB[17][3] ), .S(\mult_20/SUMB[17][3] ) );
  FA_X1 \mult_20/S2_17_2  ( .A(\mult_20/ab[17][2] ), .B(
        \mult_20/CARRYB[16][2] ), .CI(\mult_20/SUMB[16][3] ), .CO(
        \mult_20/CARRYB[17][2] ), .S(\mult_20/SUMB[17][2] ) );
  FA_X1 \mult_20/S2_17_1  ( .A(\mult_20/ab[17][1] ), .B(
        \mult_20/CARRYB[16][1] ), .CI(\mult_20/SUMB[16][2] ), .CO(
        \mult_20/CARRYB[17][1] ), .S(\mult_20/SUMB[17][1] ) );
  FA_X1 \mult_20/S1_17_0  ( .A(\mult_20/ab[17][0] ), .B(
        \mult_20/CARRYB[16][0] ), .CI(\mult_20/SUMB[16][1] ), .CO(
        \mult_20/CARRYB[17][0] ), .S(N81) );
  FA_X1 \mult_20/S3_18_30  ( .A(\mult_20/ab[18][30] ), .B(
        \mult_20/CARRYB[17][30] ), .CI(\mult_20/ab[17][31] ), .CO(
        \mult_20/CARRYB[18][30] ), .S(\mult_20/SUMB[18][30] ) );
  FA_X1 \mult_20/S2_18_29  ( .A(\mult_20/ab[18][29] ), .B(
        \mult_20/CARRYB[17][29] ), .CI(\mult_20/SUMB[17][30] ), .CO(
        \mult_20/CARRYB[18][29] ), .S(\mult_20/SUMB[18][29] ) );
  FA_X1 \mult_20/S2_18_28  ( .A(\mult_20/ab[18][28] ), .B(
        \mult_20/CARRYB[17][28] ), .CI(\mult_20/SUMB[17][29] ), .CO(
        \mult_20/CARRYB[18][28] ), .S(\mult_20/SUMB[18][28] ) );
  FA_X1 \mult_20/S2_18_27  ( .A(\mult_20/ab[18][27] ), .B(
        \mult_20/CARRYB[17][27] ), .CI(\mult_20/SUMB[17][28] ), .CO(
        \mult_20/CARRYB[18][27] ), .S(\mult_20/SUMB[18][27] ) );
  FA_X1 \mult_20/S2_18_26  ( .A(\mult_20/ab[18][26] ), .B(
        \mult_20/CARRYB[17][26] ), .CI(\mult_20/SUMB[17][27] ), .CO(
        \mult_20/CARRYB[18][26] ), .S(\mult_20/SUMB[18][26] ) );
  FA_X1 \mult_20/S2_18_25  ( .A(\mult_20/ab[18][25] ), .B(
        \mult_20/CARRYB[17][25] ), .CI(\mult_20/SUMB[17][26] ), .CO(
        \mult_20/CARRYB[18][25] ), .S(\mult_20/SUMB[18][25] ) );
  FA_X1 \mult_20/S2_18_24  ( .A(\mult_20/ab[18][24] ), .B(
        \mult_20/CARRYB[17][24] ), .CI(\mult_20/SUMB[17][25] ), .CO(
        \mult_20/CARRYB[18][24] ), .S(\mult_20/SUMB[18][24] ) );
  FA_X1 \mult_20/S2_18_23  ( .A(\mult_20/ab[18][23] ), .B(
        \mult_20/CARRYB[17][23] ), .CI(\mult_20/SUMB[17][24] ), .CO(
        \mult_20/CARRYB[18][23] ), .S(\mult_20/SUMB[18][23] ) );
  FA_X1 \mult_20/S2_18_22  ( .A(\mult_20/ab[18][22] ), .B(
        \mult_20/CARRYB[17][22] ), .CI(\mult_20/SUMB[17][23] ), .CO(
        \mult_20/CARRYB[18][22] ), .S(\mult_20/SUMB[18][22] ) );
  FA_X1 \mult_20/S2_18_21  ( .A(\mult_20/ab[18][21] ), .B(
        \mult_20/CARRYB[17][21] ), .CI(\mult_20/SUMB[17][22] ), .CO(
        \mult_20/CARRYB[18][21] ), .S(\mult_20/SUMB[18][21] ) );
  FA_X1 \mult_20/S2_18_20  ( .A(\mult_20/ab[18][20] ), .B(
        \mult_20/CARRYB[17][20] ), .CI(\mult_20/SUMB[17][21] ), .CO(
        \mult_20/CARRYB[18][20] ), .S(\mult_20/SUMB[18][20] ) );
  FA_X1 \mult_20/S2_18_19  ( .A(\mult_20/ab[18][19] ), .B(
        \mult_20/CARRYB[17][19] ), .CI(\mult_20/SUMB[17][20] ), .CO(
        \mult_20/CARRYB[18][19] ), .S(\mult_20/SUMB[18][19] ) );
  FA_X1 \mult_20/S2_18_18  ( .A(\mult_20/ab[18][18] ), .B(
        \mult_20/CARRYB[17][18] ), .CI(\mult_20/SUMB[17][19] ), .CO(
        \mult_20/CARRYB[18][18] ), .S(\mult_20/SUMB[18][18] ) );
  FA_X1 \mult_20/S2_18_17  ( .A(\mult_20/ab[18][17] ), .B(
        \mult_20/CARRYB[17][17] ), .CI(\mult_20/SUMB[17][18] ), .CO(
        \mult_20/CARRYB[18][17] ), .S(\mult_20/SUMB[18][17] ) );
  FA_X1 \mult_20/S2_18_16  ( .A(\mult_20/ab[18][16] ), .B(
        \mult_20/CARRYB[17][16] ), .CI(\mult_20/SUMB[17][17] ), .CO(
        \mult_20/CARRYB[18][16] ), .S(\mult_20/SUMB[18][16] ) );
  FA_X1 \mult_20/S2_18_15  ( .A(\mult_20/ab[18][15] ), .B(
        \mult_20/CARRYB[17][15] ), .CI(\mult_20/SUMB[17][16] ), .CO(
        \mult_20/CARRYB[18][15] ), .S(\mult_20/SUMB[18][15] ) );
  FA_X1 \mult_20/S2_18_14  ( .A(\mult_20/ab[18][14] ), .B(
        \mult_20/CARRYB[17][14] ), .CI(\mult_20/SUMB[17][15] ), .CO(
        \mult_20/CARRYB[18][14] ), .S(\mult_20/SUMB[18][14] ) );
  FA_X1 \mult_20/S2_18_13  ( .A(\mult_20/ab[18][13] ), .B(
        \mult_20/CARRYB[17][13] ), .CI(\mult_20/SUMB[17][14] ), .CO(
        \mult_20/CARRYB[18][13] ), .S(\mult_20/SUMB[18][13] ) );
  FA_X1 \mult_20/S2_18_12  ( .A(\mult_20/ab[18][12] ), .B(
        \mult_20/CARRYB[17][12] ), .CI(\mult_20/SUMB[17][13] ), .CO(
        \mult_20/CARRYB[18][12] ), .S(\mult_20/SUMB[18][12] ) );
  FA_X1 \mult_20/S2_18_11  ( .A(\mult_20/ab[18][11] ), .B(
        \mult_20/CARRYB[17][11] ), .CI(\mult_20/SUMB[17][12] ), .CO(
        \mult_20/CARRYB[18][11] ), .S(\mult_20/SUMB[18][11] ) );
  FA_X1 \mult_20/S2_18_10  ( .A(\mult_20/ab[18][10] ), .B(
        \mult_20/CARRYB[17][10] ), .CI(\mult_20/SUMB[17][11] ), .CO(
        \mult_20/CARRYB[18][10] ), .S(\mult_20/SUMB[18][10] ) );
  FA_X1 \mult_20/S2_18_9  ( .A(\mult_20/ab[18][9] ), .B(
        \mult_20/CARRYB[17][9] ), .CI(\mult_20/SUMB[17][10] ), .CO(
        \mult_20/CARRYB[18][9] ), .S(\mult_20/SUMB[18][9] ) );
  FA_X1 \mult_20/S2_18_8  ( .A(\mult_20/ab[18][8] ), .B(
        \mult_20/CARRYB[17][8] ), .CI(\mult_20/SUMB[17][9] ), .CO(
        \mult_20/CARRYB[18][8] ), .S(\mult_20/SUMB[18][8] ) );
  FA_X1 \mult_20/S2_18_7  ( .A(\mult_20/ab[18][7] ), .B(
        \mult_20/CARRYB[17][7] ), .CI(\mult_20/SUMB[17][8] ), .CO(
        \mult_20/CARRYB[18][7] ), .S(\mult_20/SUMB[18][7] ) );
  FA_X1 \mult_20/S2_18_6  ( .A(\mult_20/ab[18][6] ), .B(
        \mult_20/CARRYB[17][6] ), .CI(\mult_20/SUMB[17][7] ), .CO(
        \mult_20/CARRYB[18][6] ), .S(\mult_20/SUMB[18][6] ) );
  FA_X1 \mult_20/S2_18_5  ( .A(\mult_20/ab[18][5] ), .B(
        \mult_20/CARRYB[17][5] ), .CI(\mult_20/SUMB[17][6] ), .CO(
        \mult_20/CARRYB[18][5] ), .S(\mult_20/SUMB[18][5] ) );
  FA_X1 \mult_20/S2_18_4  ( .A(\mult_20/ab[18][4] ), .B(
        \mult_20/CARRYB[17][4] ), .CI(\mult_20/SUMB[17][5] ), .CO(
        \mult_20/CARRYB[18][4] ), .S(\mult_20/SUMB[18][4] ) );
  FA_X1 \mult_20/S2_18_3  ( .A(\mult_20/ab[18][3] ), .B(
        \mult_20/CARRYB[17][3] ), .CI(\mult_20/SUMB[17][4] ), .CO(
        \mult_20/CARRYB[18][3] ), .S(\mult_20/SUMB[18][3] ) );
  FA_X1 \mult_20/S2_18_2  ( .A(\mult_20/ab[18][2] ), .B(
        \mult_20/CARRYB[17][2] ), .CI(\mult_20/SUMB[17][3] ), .CO(
        \mult_20/CARRYB[18][2] ), .S(\mult_20/SUMB[18][2] ) );
  FA_X1 \mult_20/S2_18_1  ( .A(\mult_20/ab[18][1] ), .B(
        \mult_20/CARRYB[17][1] ), .CI(\mult_20/SUMB[17][2] ), .CO(
        \mult_20/CARRYB[18][1] ), .S(\mult_20/SUMB[18][1] ) );
  FA_X1 \mult_20/S1_18_0  ( .A(\mult_20/ab[18][0] ), .B(
        \mult_20/CARRYB[17][0] ), .CI(\mult_20/SUMB[17][1] ), .CO(
        \mult_20/CARRYB[18][0] ), .S(N82) );
  FA_X1 \mult_20/S3_19_30  ( .A(\mult_20/ab[19][30] ), .B(
        \mult_20/CARRYB[18][30] ), .CI(\mult_20/ab[18][31] ), .CO(
        \mult_20/CARRYB[19][30] ), .S(\mult_20/SUMB[19][30] ) );
  FA_X1 \mult_20/S2_19_29  ( .A(\mult_20/ab[19][29] ), .B(
        \mult_20/CARRYB[18][29] ), .CI(\mult_20/SUMB[18][30] ), .CO(
        \mult_20/CARRYB[19][29] ), .S(\mult_20/SUMB[19][29] ) );
  FA_X1 \mult_20/S2_19_28  ( .A(\mult_20/ab[19][28] ), .B(
        \mult_20/CARRYB[18][28] ), .CI(\mult_20/SUMB[18][29] ), .CO(
        \mult_20/CARRYB[19][28] ), .S(\mult_20/SUMB[19][28] ) );
  FA_X1 \mult_20/S2_19_27  ( .A(\mult_20/ab[19][27] ), .B(
        \mult_20/CARRYB[18][27] ), .CI(\mult_20/SUMB[18][28] ), .CO(
        \mult_20/CARRYB[19][27] ), .S(\mult_20/SUMB[19][27] ) );
  FA_X1 \mult_20/S2_19_26  ( .A(\mult_20/ab[19][26] ), .B(
        \mult_20/CARRYB[18][26] ), .CI(\mult_20/SUMB[18][27] ), .CO(
        \mult_20/CARRYB[19][26] ), .S(\mult_20/SUMB[19][26] ) );
  FA_X1 \mult_20/S2_19_25  ( .A(\mult_20/ab[19][25] ), .B(
        \mult_20/CARRYB[18][25] ), .CI(\mult_20/SUMB[18][26] ), .CO(
        \mult_20/CARRYB[19][25] ), .S(\mult_20/SUMB[19][25] ) );
  FA_X1 \mult_20/S2_19_24  ( .A(\mult_20/ab[19][24] ), .B(
        \mult_20/CARRYB[18][24] ), .CI(\mult_20/SUMB[18][25] ), .CO(
        \mult_20/CARRYB[19][24] ), .S(\mult_20/SUMB[19][24] ) );
  FA_X1 \mult_20/S2_19_23  ( .A(\mult_20/ab[19][23] ), .B(
        \mult_20/CARRYB[18][23] ), .CI(\mult_20/SUMB[18][24] ), .CO(
        \mult_20/CARRYB[19][23] ), .S(\mult_20/SUMB[19][23] ) );
  FA_X1 \mult_20/S2_19_22  ( .A(\mult_20/ab[19][22] ), .B(
        \mult_20/CARRYB[18][22] ), .CI(\mult_20/SUMB[18][23] ), .CO(
        \mult_20/CARRYB[19][22] ), .S(\mult_20/SUMB[19][22] ) );
  FA_X1 \mult_20/S2_19_21  ( .A(\mult_20/ab[19][21] ), .B(
        \mult_20/CARRYB[18][21] ), .CI(\mult_20/SUMB[18][22] ), .CO(
        \mult_20/CARRYB[19][21] ), .S(\mult_20/SUMB[19][21] ) );
  FA_X1 \mult_20/S2_19_20  ( .A(\mult_20/ab[19][20] ), .B(
        \mult_20/CARRYB[18][20] ), .CI(\mult_20/SUMB[18][21] ), .CO(
        \mult_20/CARRYB[19][20] ), .S(\mult_20/SUMB[19][20] ) );
  FA_X1 \mult_20/S2_19_19  ( .A(\mult_20/ab[19][19] ), .B(
        \mult_20/CARRYB[18][19] ), .CI(\mult_20/SUMB[18][20] ), .CO(
        \mult_20/CARRYB[19][19] ), .S(\mult_20/SUMB[19][19] ) );
  FA_X1 \mult_20/S2_19_18  ( .A(\mult_20/ab[19][18] ), .B(
        \mult_20/CARRYB[18][18] ), .CI(\mult_20/SUMB[18][19] ), .CO(
        \mult_20/CARRYB[19][18] ), .S(\mult_20/SUMB[19][18] ) );
  FA_X1 \mult_20/S2_19_17  ( .A(\mult_20/ab[19][17] ), .B(
        \mult_20/CARRYB[18][17] ), .CI(\mult_20/SUMB[18][18] ), .CO(
        \mult_20/CARRYB[19][17] ), .S(\mult_20/SUMB[19][17] ) );
  FA_X1 \mult_20/S2_19_16  ( .A(\mult_20/ab[19][16] ), .B(
        \mult_20/CARRYB[18][16] ), .CI(\mult_20/SUMB[18][17] ), .CO(
        \mult_20/CARRYB[19][16] ), .S(\mult_20/SUMB[19][16] ) );
  FA_X1 \mult_20/S2_19_15  ( .A(\mult_20/ab[19][15] ), .B(
        \mult_20/CARRYB[18][15] ), .CI(\mult_20/SUMB[18][16] ), .CO(
        \mult_20/CARRYB[19][15] ), .S(\mult_20/SUMB[19][15] ) );
  FA_X1 \mult_20/S2_19_14  ( .A(\mult_20/ab[19][14] ), .B(
        \mult_20/CARRYB[18][14] ), .CI(\mult_20/SUMB[18][15] ), .CO(
        \mult_20/CARRYB[19][14] ), .S(\mult_20/SUMB[19][14] ) );
  FA_X1 \mult_20/S2_19_13  ( .A(\mult_20/ab[19][13] ), .B(
        \mult_20/CARRYB[18][13] ), .CI(\mult_20/SUMB[18][14] ), .CO(
        \mult_20/CARRYB[19][13] ), .S(\mult_20/SUMB[19][13] ) );
  FA_X1 \mult_20/S2_19_12  ( .A(\mult_20/ab[19][12] ), .B(
        \mult_20/CARRYB[18][12] ), .CI(\mult_20/SUMB[18][13] ), .CO(
        \mult_20/CARRYB[19][12] ), .S(\mult_20/SUMB[19][12] ) );
  FA_X1 \mult_20/S2_19_11  ( .A(\mult_20/ab[19][11] ), .B(
        \mult_20/CARRYB[18][11] ), .CI(\mult_20/SUMB[18][12] ), .CO(
        \mult_20/CARRYB[19][11] ), .S(\mult_20/SUMB[19][11] ) );
  FA_X1 \mult_20/S2_19_10  ( .A(\mult_20/ab[19][10] ), .B(
        \mult_20/CARRYB[18][10] ), .CI(\mult_20/SUMB[18][11] ), .CO(
        \mult_20/CARRYB[19][10] ), .S(\mult_20/SUMB[19][10] ) );
  FA_X1 \mult_20/S2_19_9  ( .A(\mult_20/ab[19][9] ), .B(
        \mult_20/CARRYB[18][9] ), .CI(\mult_20/SUMB[18][10] ), .CO(
        \mult_20/CARRYB[19][9] ), .S(\mult_20/SUMB[19][9] ) );
  FA_X1 \mult_20/S2_19_8  ( .A(\mult_20/ab[19][8] ), .B(
        \mult_20/CARRYB[18][8] ), .CI(\mult_20/SUMB[18][9] ), .CO(
        \mult_20/CARRYB[19][8] ), .S(\mult_20/SUMB[19][8] ) );
  FA_X1 \mult_20/S2_19_7  ( .A(\mult_20/ab[19][7] ), .B(
        \mult_20/CARRYB[18][7] ), .CI(\mult_20/SUMB[18][8] ), .CO(
        \mult_20/CARRYB[19][7] ), .S(\mult_20/SUMB[19][7] ) );
  FA_X1 \mult_20/S2_19_6  ( .A(\mult_20/ab[19][6] ), .B(
        \mult_20/CARRYB[18][6] ), .CI(\mult_20/SUMB[18][7] ), .CO(
        \mult_20/CARRYB[19][6] ), .S(\mult_20/SUMB[19][6] ) );
  FA_X1 \mult_20/S2_19_5  ( .A(\mult_20/ab[19][5] ), .B(
        \mult_20/CARRYB[18][5] ), .CI(\mult_20/SUMB[18][6] ), .CO(
        \mult_20/CARRYB[19][5] ), .S(\mult_20/SUMB[19][5] ) );
  FA_X1 \mult_20/S2_19_4  ( .A(\mult_20/ab[19][4] ), .B(
        \mult_20/CARRYB[18][4] ), .CI(\mult_20/SUMB[18][5] ), .CO(
        \mult_20/CARRYB[19][4] ), .S(\mult_20/SUMB[19][4] ) );
  FA_X1 \mult_20/S2_19_3  ( .A(\mult_20/ab[19][3] ), .B(
        \mult_20/CARRYB[18][3] ), .CI(\mult_20/SUMB[18][4] ), .CO(
        \mult_20/CARRYB[19][3] ), .S(\mult_20/SUMB[19][3] ) );
  FA_X1 \mult_20/S2_19_2  ( .A(\mult_20/ab[19][2] ), .B(
        \mult_20/CARRYB[18][2] ), .CI(\mult_20/SUMB[18][3] ), .CO(
        \mult_20/CARRYB[19][2] ), .S(\mult_20/SUMB[19][2] ) );
  FA_X1 \mult_20/S2_19_1  ( .A(\mult_20/ab[19][1] ), .B(
        \mult_20/CARRYB[18][1] ), .CI(\mult_20/SUMB[18][2] ), .CO(
        \mult_20/CARRYB[19][1] ), .S(\mult_20/SUMB[19][1] ) );
  FA_X1 \mult_20/S1_19_0  ( .A(\mult_20/ab[19][0] ), .B(
        \mult_20/CARRYB[18][0] ), .CI(\mult_20/SUMB[18][1] ), .CO(
        \mult_20/CARRYB[19][0] ), .S(N83) );
  FA_X1 \mult_20/S3_20_30  ( .A(\mult_20/ab[20][30] ), .B(
        \mult_20/CARRYB[19][30] ), .CI(\mult_20/ab[19][31] ), .CO(
        \mult_20/CARRYB[20][30] ), .S(\mult_20/SUMB[20][30] ) );
  FA_X1 \mult_20/S2_20_29  ( .A(\mult_20/ab[20][29] ), .B(
        \mult_20/CARRYB[19][29] ), .CI(\mult_20/SUMB[19][30] ), .CO(
        \mult_20/CARRYB[20][29] ), .S(\mult_20/SUMB[20][29] ) );
  FA_X1 \mult_20/S2_20_28  ( .A(\mult_20/ab[20][28] ), .B(
        \mult_20/CARRYB[19][28] ), .CI(\mult_20/SUMB[19][29] ), .CO(
        \mult_20/CARRYB[20][28] ), .S(\mult_20/SUMB[20][28] ) );
  FA_X1 \mult_20/S2_20_27  ( .A(\mult_20/ab[20][27] ), .B(
        \mult_20/CARRYB[19][27] ), .CI(\mult_20/SUMB[19][28] ), .CO(
        \mult_20/CARRYB[20][27] ), .S(\mult_20/SUMB[20][27] ) );
  FA_X1 \mult_20/S2_20_26  ( .A(\mult_20/ab[20][26] ), .B(
        \mult_20/CARRYB[19][26] ), .CI(\mult_20/SUMB[19][27] ), .CO(
        \mult_20/CARRYB[20][26] ), .S(\mult_20/SUMB[20][26] ) );
  FA_X1 \mult_20/S2_20_25  ( .A(\mult_20/ab[20][25] ), .B(
        \mult_20/CARRYB[19][25] ), .CI(\mult_20/SUMB[19][26] ), .CO(
        \mult_20/CARRYB[20][25] ), .S(\mult_20/SUMB[20][25] ) );
  FA_X1 \mult_20/S2_20_24  ( .A(\mult_20/ab[20][24] ), .B(
        \mult_20/CARRYB[19][24] ), .CI(\mult_20/SUMB[19][25] ), .CO(
        \mult_20/CARRYB[20][24] ), .S(\mult_20/SUMB[20][24] ) );
  FA_X1 \mult_20/S2_20_23  ( .A(\mult_20/ab[20][23] ), .B(
        \mult_20/CARRYB[19][23] ), .CI(\mult_20/SUMB[19][24] ), .CO(
        \mult_20/CARRYB[20][23] ), .S(\mult_20/SUMB[20][23] ) );
  FA_X1 \mult_20/S2_20_22  ( .A(\mult_20/ab[20][22] ), .B(
        \mult_20/CARRYB[19][22] ), .CI(\mult_20/SUMB[19][23] ), .CO(
        \mult_20/CARRYB[20][22] ), .S(\mult_20/SUMB[20][22] ) );
  FA_X1 \mult_20/S2_20_21  ( .A(\mult_20/ab[20][21] ), .B(
        \mult_20/CARRYB[19][21] ), .CI(\mult_20/SUMB[19][22] ), .CO(
        \mult_20/CARRYB[20][21] ), .S(\mult_20/SUMB[20][21] ) );
  FA_X1 \mult_20/S2_20_20  ( .A(\mult_20/ab[20][20] ), .B(
        \mult_20/CARRYB[19][20] ), .CI(\mult_20/SUMB[19][21] ), .CO(
        \mult_20/CARRYB[20][20] ), .S(\mult_20/SUMB[20][20] ) );
  FA_X1 \mult_20/S2_20_19  ( .A(\mult_20/ab[20][19] ), .B(
        \mult_20/CARRYB[19][19] ), .CI(\mult_20/SUMB[19][20] ), .CO(
        \mult_20/CARRYB[20][19] ), .S(\mult_20/SUMB[20][19] ) );
  FA_X1 \mult_20/S2_20_18  ( .A(\mult_20/ab[20][18] ), .B(
        \mult_20/CARRYB[19][18] ), .CI(\mult_20/SUMB[19][19] ), .CO(
        \mult_20/CARRYB[20][18] ), .S(\mult_20/SUMB[20][18] ) );
  FA_X1 \mult_20/S2_20_17  ( .A(\mult_20/ab[20][17] ), .B(
        \mult_20/CARRYB[19][17] ), .CI(\mult_20/SUMB[19][18] ), .CO(
        \mult_20/CARRYB[20][17] ), .S(\mult_20/SUMB[20][17] ) );
  FA_X1 \mult_20/S2_20_16  ( .A(\mult_20/ab[20][16] ), .B(
        \mult_20/CARRYB[19][16] ), .CI(\mult_20/SUMB[19][17] ), .CO(
        \mult_20/CARRYB[20][16] ), .S(\mult_20/SUMB[20][16] ) );
  FA_X1 \mult_20/S2_20_15  ( .A(\mult_20/ab[20][15] ), .B(
        \mult_20/CARRYB[19][15] ), .CI(\mult_20/SUMB[19][16] ), .CO(
        \mult_20/CARRYB[20][15] ), .S(\mult_20/SUMB[20][15] ) );
  FA_X1 \mult_20/S2_20_14  ( .A(\mult_20/ab[20][14] ), .B(
        \mult_20/CARRYB[19][14] ), .CI(\mult_20/SUMB[19][15] ), .CO(
        \mult_20/CARRYB[20][14] ), .S(\mult_20/SUMB[20][14] ) );
  FA_X1 \mult_20/S2_20_13  ( .A(\mult_20/ab[20][13] ), .B(
        \mult_20/CARRYB[19][13] ), .CI(\mult_20/SUMB[19][14] ), .CO(
        \mult_20/CARRYB[20][13] ), .S(\mult_20/SUMB[20][13] ) );
  FA_X1 \mult_20/S2_20_12  ( .A(\mult_20/ab[20][12] ), .B(
        \mult_20/CARRYB[19][12] ), .CI(\mult_20/SUMB[19][13] ), .CO(
        \mult_20/CARRYB[20][12] ), .S(\mult_20/SUMB[20][12] ) );
  FA_X1 \mult_20/S2_20_11  ( .A(\mult_20/ab[20][11] ), .B(
        \mult_20/CARRYB[19][11] ), .CI(\mult_20/SUMB[19][12] ), .CO(
        \mult_20/CARRYB[20][11] ), .S(\mult_20/SUMB[20][11] ) );
  FA_X1 \mult_20/S2_20_10  ( .A(\mult_20/ab[20][10] ), .B(
        \mult_20/CARRYB[19][10] ), .CI(\mult_20/SUMB[19][11] ), .CO(
        \mult_20/CARRYB[20][10] ), .S(\mult_20/SUMB[20][10] ) );
  FA_X1 \mult_20/S2_20_9  ( .A(\mult_20/ab[20][9] ), .B(
        \mult_20/CARRYB[19][9] ), .CI(\mult_20/SUMB[19][10] ), .CO(
        \mult_20/CARRYB[20][9] ), .S(\mult_20/SUMB[20][9] ) );
  FA_X1 \mult_20/S2_20_8  ( .A(\mult_20/ab[20][8] ), .B(
        \mult_20/CARRYB[19][8] ), .CI(\mult_20/SUMB[19][9] ), .CO(
        \mult_20/CARRYB[20][8] ), .S(\mult_20/SUMB[20][8] ) );
  FA_X1 \mult_20/S2_20_7  ( .A(\mult_20/ab[20][7] ), .B(
        \mult_20/CARRYB[19][7] ), .CI(\mult_20/SUMB[19][8] ), .CO(
        \mult_20/CARRYB[20][7] ), .S(\mult_20/SUMB[20][7] ) );
  FA_X1 \mult_20/S2_20_6  ( .A(\mult_20/ab[20][6] ), .B(
        \mult_20/CARRYB[19][6] ), .CI(\mult_20/SUMB[19][7] ), .CO(
        \mult_20/CARRYB[20][6] ), .S(\mult_20/SUMB[20][6] ) );
  FA_X1 \mult_20/S2_20_5  ( .A(\mult_20/ab[20][5] ), .B(
        \mult_20/CARRYB[19][5] ), .CI(\mult_20/SUMB[19][6] ), .CO(
        \mult_20/CARRYB[20][5] ), .S(\mult_20/SUMB[20][5] ) );
  FA_X1 \mult_20/S2_20_4  ( .A(\mult_20/ab[20][4] ), .B(
        \mult_20/CARRYB[19][4] ), .CI(\mult_20/SUMB[19][5] ), .CO(
        \mult_20/CARRYB[20][4] ), .S(\mult_20/SUMB[20][4] ) );
  FA_X1 \mult_20/S2_20_3  ( .A(\mult_20/ab[20][3] ), .B(
        \mult_20/CARRYB[19][3] ), .CI(\mult_20/SUMB[19][4] ), .CO(
        \mult_20/CARRYB[20][3] ), .S(\mult_20/SUMB[20][3] ) );
  FA_X1 \mult_20/S2_20_2  ( .A(\mult_20/ab[20][2] ), .B(
        \mult_20/CARRYB[19][2] ), .CI(\mult_20/SUMB[19][3] ), .CO(
        \mult_20/CARRYB[20][2] ), .S(\mult_20/SUMB[20][2] ) );
  FA_X1 \mult_20/S2_20_1  ( .A(\mult_20/ab[20][1] ), .B(
        \mult_20/CARRYB[19][1] ), .CI(\mult_20/SUMB[19][2] ), .CO(
        \mult_20/CARRYB[20][1] ), .S(\mult_20/SUMB[20][1] ) );
  FA_X1 \mult_20/S1_20_0  ( .A(\mult_20/ab[20][0] ), .B(
        \mult_20/CARRYB[19][0] ), .CI(\mult_20/SUMB[19][1] ), .CO(
        \mult_20/CARRYB[20][0] ), .S(N84) );
  FA_X1 \mult_20/S3_21_30  ( .A(\mult_20/ab[21][30] ), .B(
        \mult_20/CARRYB[20][30] ), .CI(\mult_20/ab[20][31] ), .CO(
        \mult_20/CARRYB[21][30] ), .S(\mult_20/SUMB[21][30] ) );
  FA_X1 \mult_20/S2_21_29  ( .A(\mult_20/ab[21][29] ), .B(
        \mult_20/CARRYB[20][29] ), .CI(\mult_20/SUMB[20][30] ), .CO(
        \mult_20/CARRYB[21][29] ), .S(\mult_20/SUMB[21][29] ) );
  FA_X1 \mult_20/S2_21_28  ( .A(\mult_20/ab[21][28] ), .B(
        \mult_20/CARRYB[20][28] ), .CI(\mult_20/SUMB[20][29] ), .CO(
        \mult_20/CARRYB[21][28] ), .S(\mult_20/SUMB[21][28] ) );
  FA_X1 \mult_20/S2_21_27  ( .A(\mult_20/ab[21][27] ), .B(
        \mult_20/CARRYB[20][27] ), .CI(\mult_20/SUMB[20][28] ), .CO(
        \mult_20/CARRYB[21][27] ), .S(\mult_20/SUMB[21][27] ) );
  FA_X1 \mult_20/S2_21_26  ( .A(\mult_20/ab[21][26] ), .B(
        \mult_20/CARRYB[20][26] ), .CI(\mult_20/SUMB[20][27] ), .CO(
        \mult_20/CARRYB[21][26] ), .S(\mult_20/SUMB[21][26] ) );
  FA_X1 \mult_20/S2_21_25  ( .A(\mult_20/ab[21][25] ), .B(
        \mult_20/CARRYB[20][25] ), .CI(\mult_20/SUMB[20][26] ), .CO(
        \mult_20/CARRYB[21][25] ), .S(\mult_20/SUMB[21][25] ) );
  FA_X1 \mult_20/S2_21_24  ( .A(\mult_20/ab[21][24] ), .B(
        \mult_20/CARRYB[20][24] ), .CI(\mult_20/SUMB[20][25] ), .CO(
        \mult_20/CARRYB[21][24] ), .S(\mult_20/SUMB[21][24] ) );
  FA_X1 \mult_20/S2_21_23  ( .A(\mult_20/ab[21][23] ), .B(
        \mult_20/CARRYB[20][23] ), .CI(\mult_20/SUMB[20][24] ), .CO(
        \mult_20/CARRYB[21][23] ), .S(\mult_20/SUMB[21][23] ) );
  FA_X1 \mult_20/S2_21_22  ( .A(\mult_20/ab[21][22] ), .B(
        \mult_20/CARRYB[20][22] ), .CI(\mult_20/SUMB[20][23] ), .CO(
        \mult_20/CARRYB[21][22] ), .S(\mult_20/SUMB[21][22] ) );
  FA_X1 \mult_20/S2_21_21  ( .A(\mult_20/ab[21][21] ), .B(
        \mult_20/CARRYB[20][21] ), .CI(\mult_20/SUMB[20][22] ), .CO(
        \mult_20/CARRYB[21][21] ), .S(\mult_20/SUMB[21][21] ) );
  FA_X1 \mult_20/S2_21_20  ( .A(\mult_20/ab[21][20] ), .B(
        \mult_20/CARRYB[20][20] ), .CI(\mult_20/SUMB[20][21] ), .CO(
        \mult_20/CARRYB[21][20] ), .S(\mult_20/SUMB[21][20] ) );
  FA_X1 \mult_20/S2_21_19  ( .A(\mult_20/ab[21][19] ), .B(
        \mult_20/CARRYB[20][19] ), .CI(\mult_20/SUMB[20][20] ), .CO(
        \mult_20/CARRYB[21][19] ), .S(\mult_20/SUMB[21][19] ) );
  FA_X1 \mult_20/S2_21_18  ( .A(\mult_20/ab[21][18] ), .B(
        \mult_20/CARRYB[20][18] ), .CI(\mult_20/SUMB[20][19] ), .CO(
        \mult_20/CARRYB[21][18] ), .S(\mult_20/SUMB[21][18] ) );
  FA_X1 \mult_20/S2_21_17  ( .A(\mult_20/ab[21][17] ), .B(
        \mult_20/CARRYB[20][17] ), .CI(\mult_20/SUMB[20][18] ), .CO(
        \mult_20/CARRYB[21][17] ), .S(\mult_20/SUMB[21][17] ) );
  FA_X1 \mult_20/S2_21_16  ( .A(\mult_20/ab[21][16] ), .B(
        \mult_20/CARRYB[20][16] ), .CI(\mult_20/SUMB[20][17] ), .CO(
        \mult_20/CARRYB[21][16] ), .S(\mult_20/SUMB[21][16] ) );
  FA_X1 \mult_20/S2_21_15  ( .A(\mult_20/ab[21][15] ), .B(
        \mult_20/CARRYB[20][15] ), .CI(\mult_20/SUMB[20][16] ), .CO(
        \mult_20/CARRYB[21][15] ), .S(\mult_20/SUMB[21][15] ) );
  FA_X1 \mult_20/S2_21_14  ( .A(\mult_20/ab[21][14] ), .B(
        \mult_20/CARRYB[20][14] ), .CI(\mult_20/SUMB[20][15] ), .CO(
        \mult_20/CARRYB[21][14] ), .S(\mult_20/SUMB[21][14] ) );
  FA_X1 \mult_20/S2_21_13  ( .A(\mult_20/ab[21][13] ), .B(
        \mult_20/CARRYB[20][13] ), .CI(\mult_20/SUMB[20][14] ), .CO(
        \mult_20/CARRYB[21][13] ), .S(\mult_20/SUMB[21][13] ) );
  FA_X1 \mult_20/S2_21_12  ( .A(\mult_20/ab[21][12] ), .B(
        \mult_20/CARRYB[20][12] ), .CI(\mult_20/SUMB[20][13] ), .CO(
        \mult_20/CARRYB[21][12] ), .S(\mult_20/SUMB[21][12] ) );
  FA_X1 \mult_20/S2_21_11  ( .A(\mult_20/ab[21][11] ), .B(
        \mult_20/CARRYB[20][11] ), .CI(\mult_20/SUMB[20][12] ), .CO(
        \mult_20/CARRYB[21][11] ), .S(\mult_20/SUMB[21][11] ) );
  FA_X1 \mult_20/S2_21_10  ( .A(\mult_20/ab[21][10] ), .B(
        \mult_20/CARRYB[20][10] ), .CI(\mult_20/SUMB[20][11] ), .CO(
        \mult_20/CARRYB[21][10] ), .S(\mult_20/SUMB[21][10] ) );
  FA_X1 \mult_20/S2_21_9  ( .A(\mult_20/ab[21][9] ), .B(
        \mult_20/CARRYB[20][9] ), .CI(\mult_20/SUMB[20][10] ), .CO(
        \mult_20/CARRYB[21][9] ), .S(\mult_20/SUMB[21][9] ) );
  FA_X1 \mult_20/S2_21_8  ( .A(\mult_20/ab[21][8] ), .B(
        \mult_20/CARRYB[20][8] ), .CI(\mult_20/SUMB[20][9] ), .CO(
        \mult_20/CARRYB[21][8] ), .S(\mult_20/SUMB[21][8] ) );
  FA_X1 \mult_20/S2_21_7  ( .A(\mult_20/ab[21][7] ), .B(
        \mult_20/CARRYB[20][7] ), .CI(\mult_20/SUMB[20][8] ), .CO(
        \mult_20/CARRYB[21][7] ), .S(\mult_20/SUMB[21][7] ) );
  FA_X1 \mult_20/S2_21_6  ( .A(\mult_20/ab[21][6] ), .B(
        \mult_20/CARRYB[20][6] ), .CI(\mult_20/SUMB[20][7] ), .CO(
        \mult_20/CARRYB[21][6] ), .S(\mult_20/SUMB[21][6] ) );
  FA_X1 \mult_20/S2_21_5  ( .A(\mult_20/ab[21][5] ), .B(
        \mult_20/CARRYB[20][5] ), .CI(\mult_20/SUMB[20][6] ), .CO(
        \mult_20/CARRYB[21][5] ), .S(\mult_20/SUMB[21][5] ) );
  FA_X1 \mult_20/S2_21_4  ( .A(\mult_20/ab[21][4] ), .B(
        \mult_20/CARRYB[20][4] ), .CI(\mult_20/SUMB[20][5] ), .CO(
        \mult_20/CARRYB[21][4] ), .S(\mult_20/SUMB[21][4] ) );
  FA_X1 \mult_20/S2_21_3  ( .A(\mult_20/ab[21][3] ), .B(
        \mult_20/CARRYB[20][3] ), .CI(\mult_20/SUMB[20][4] ), .CO(
        \mult_20/CARRYB[21][3] ), .S(\mult_20/SUMB[21][3] ) );
  FA_X1 \mult_20/S2_21_2  ( .A(\mult_20/ab[21][2] ), .B(
        \mult_20/CARRYB[20][2] ), .CI(\mult_20/SUMB[20][3] ), .CO(
        \mult_20/CARRYB[21][2] ), .S(\mult_20/SUMB[21][2] ) );
  FA_X1 \mult_20/S2_21_1  ( .A(\mult_20/ab[21][1] ), .B(
        \mult_20/CARRYB[20][1] ), .CI(\mult_20/SUMB[20][2] ), .CO(
        \mult_20/CARRYB[21][1] ), .S(\mult_20/SUMB[21][1] ) );
  FA_X1 \mult_20/S1_21_0  ( .A(\mult_20/ab[21][0] ), .B(
        \mult_20/CARRYB[20][0] ), .CI(\mult_20/SUMB[20][1] ), .CO(
        \mult_20/CARRYB[21][0] ), .S(N85) );
  FA_X1 \mult_20/S3_22_30  ( .A(\mult_20/ab[22][30] ), .B(
        \mult_20/CARRYB[21][30] ), .CI(\mult_20/ab[21][31] ), .CO(
        \mult_20/CARRYB[22][30] ), .S(\mult_20/SUMB[22][30] ) );
  FA_X1 \mult_20/S2_22_29  ( .A(\mult_20/ab[22][29] ), .B(
        \mult_20/CARRYB[21][29] ), .CI(\mult_20/SUMB[21][30] ), .CO(
        \mult_20/CARRYB[22][29] ), .S(\mult_20/SUMB[22][29] ) );
  FA_X1 \mult_20/S2_22_28  ( .A(\mult_20/ab[22][28] ), .B(
        \mult_20/CARRYB[21][28] ), .CI(\mult_20/SUMB[21][29] ), .CO(
        \mult_20/CARRYB[22][28] ), .S(\mult_20/SUMB[22][28] ) );
  FA_X1 \mult_20/S2_22_27  ( .A(\mult_20/ab[22][27] ), .B(
        \mult_20/CARRYB[21][27] ), .CI(\mult_20/SUMB[21][28] ), .CO(
        \mult_20/CARRYB[22][27] ), .S(\mult_20/SUMB[22][27] ) );
  FA_X1 \mult_20/S2_22_26  ( .A(\mult_20/ab[22][26] ), .B(
        \mult_20/CARRYB[21][26] ), .CI(\mult_20/SUMB[21][27] ), .CO(
        \mult_20/CARRYB[22][26] ), .S(\mult_20/SUMB[22][26] ) );
  FA_X1 \mult_20/S2_22_25  ( .A(\mult_20/ab[22][25] ), .B(
        \mult_20/CARRYB[21][25] ), .CI(\mult_20/SUMB[21][26] ), .CO(
        \mult_20/CARRYB[22][25] ), .S(\mult_20/SUMB[22][25] ) );
  FA_X1 \mult_20/S2_22_24  ( .A(\mult_20/ab[22][24] ), .B(
        \mult_20/CARRYB[21][24] ), .CI(\mult_20/SUMB[21][25] ), .CO(
        \mult_20/CARRYB[22][24] ), .S(\mult_20/SUMB[22][24] ) );
  FA_X1 \mult_20/S2_22_23  ( .A(\mult_20/ab[22][23] ), .B(
        \mult_20/CARRYB[21][23] ), .CI(\mult_20/SUMB[21][24] ), .CO(
        \mult_20/CARRYB[22][23] ), .S(\mult_20/SUMB[22][23] ) );
  FA_X1 \mult_20/S2_22_22  ( .A(\mult_20/ab[22][22] ), .B(
        \mult_20/CARRYB[21][22] ), .CI(\mult_20/SUMB[21][23] ), .CO(
        \mult_20/CARRYB[22][22] ), .S(\mult_20/SUMB[22][22] ) );
  FA_X1 \mult_20/S2_22_21  ( .A(\mult_20/ab[22][21] ), .B(
        \mult_20/CARRYB[21][21] ), .CI(\mult_20/SUMB[21][22] ), .CO(
        \mult_20/CARRYB[22][21] ), .S(\mult_20/SUMB[22][21] ) );
  FA_X1 \mult_20/S2_22_20  ( .A(\mult_20/ab[22][20] ), .B(
        \mult_20/CARRYB[21][20] ), .CI(\mult_20/SUMB[21][21] ), .CO(
        \mult_20/CARRYB[22][20] ), .S(\mult_20/SUMB[22][20] ) );
  FA_X1 \mult_20/S2_22_19  ( .A(\mult_20/ab[22][19] ), .B(
        \mult_20/CARRYB[21][19] ), .CI(\mult_20/SUMB[21][20] ), .CO(
        \mult_20/CARRYB[22][19] ), .S(\mult_20/SUMB[22][19] ) );
  FA_X1 \mult_20/S2_22_18  ( .A(\mult_20/ab[22][18] ), .B(
        \mult_20/CARRYB[21][18] ), .CI(\mult_20/SUMB[21][19] ), .CO(
        \mult_20/CARRYB[22][18] ), .S(\mult_20/SUMB[22][18] ) );
  FA_X1 \mult_20/S2_22_17  ( .A(\mult_20/ab[22][17] ), .B(
        \mult_20/CARRYB[21][17] ), .CI(\mult_20/SUMB[21][18] ), .CO(
        \mult_20/CARRYB[22][17] ), .S(\mult_20/SUMB[22][17] ) );
  FA_X1 \mult_20/S2_22_16  ( .A(\mult_20/ab[22][16] ), .B(
        \mult_20/CARRYB[21][16] ), .CI(\mult_20/SUMB[21][17] ), .CO(
        \mult_20/CARRYB[22][16] ), .S(\mult_20/SUMB[22][16] ) );
  FA_X1 \mult_20/S2_22_15  ( .A(\mult_20/ab[22][15] ), .B(
        \mult_20/CARRYB[21][15] ), .CI(\mult_20/SUMB[21][16] ), .CO(
        \mult_20/CARRYB[22][15] ), .S(\mult_20/SUMB[22][15] ) );
  FA_X1 \mult_20/S2_22_14  ( .A(\mult_20/ab[22][14] ), .B(
        \mult_20/CARRYB[21][14] ), .CI(\mult_20/SUMB[21][15] ), .CO(
        \mult_20/CARRYB[22][14] ), .S(\mult_20/SUMB[22][14] ) );
  FA_X1 \mult_20/S2_22_13  ( .A(\mult_20/ab[22][13] ), .B(
        \mult_20/CARRYB[21][13] ), .CI(\mult_20/SUMB[21][14] ), .CO(
        \mult_20/CARRYB[22][13] ), .S(\mult_20/SUMB[22][13] ) );
  FA_X1 \mult_20/S2_22_12  ( .A(\mult_20/ab[22][12] ), .B(
        \mult_20/CARRYB[21][12] ), .CI(\mult_20/SUMB[21][13] ), .CO(
        \mult_20/CARRYB[22][12] ), .S(\mult_20/SUMB[22][12] ) );
  FA_X1 \mult_20/S2_22_11  ( .A(\mult_20/ab[22][11] ), .B(
        \mult_20/CARRYB[21][11] ), .CI(\mult_20/SUMB[21][12] ), .CO(
        \mult_20/CARRYB[22][11] ), .S(\mult_20/SUMB[22][11] ) );
  FA_X1 \mult_20/S2_22_10  ( .A(\mult_20/ab[22][10] ), .B(
        \mult_20/CARRYB[21][10] ), .CI(\mult_20/SUMB[21][11] ), .CO(
        \mult_20/CARRYB[22][10] ), .S(\mult_20/SUMB[22][10] ) );
  FA_X1 \mult_20/S2_22_9  ( .A(\mult_20/ab[22][9] ), .B(
        \mult_20/CARRYB[21][9] ), .CI(\mult_20/SUMB[21][10] ), .CO(
        \mult_20/CARRYB[22][9] ), .S(\mult_20/SUMB[22][9] ) );
  FA_X1 \mult_20/S2_22_8  ( .A(\mult_20/ab[22][8] ), .B(
        \mult_20/CARRYB[21][8] ), .CI(\mult_20/SUMB[21][9] ), .CO(
        \mult_20/CARRYB[22][8] ), .S(\mult_20/SUMB[22][8] ) );
  FA_X1 \mult_20/S2_22_7  ( .A(\mult_20/ab[22][7] ), .B(
        \mult_20/CARRYB[21][7] ), .CI(\mult_20/SUMB[21][8] ), .CO(
        \mult_20/CARRYB[22][7] ), .S(\mult_20/SUMB[22][7] ) );
  FA_X1 \mult_20/S2_22_6  ( .A(\mult_20/ab[22][6] ), .B(
        \mult_20/CARRYB[21][6] ), .CI(\mult_20/SUMB[21][7] ), .CO(
        \mult_20/CARRYB[22][6] ), .S(\mult_20/SUMB[22][6] ) );
  FA_X1 \mult_20/S2_22_5  ( .A(\mult_20/ab[22][5] ), .B(
        \mult_20/CARRYB[21][5] ), .CI(\mult_20/SUMB[21][6] ), .CO(
        \mult_20/CARRYB[22][5] ), .S(\mult_20/SUMB[22][5] ) );
  FA_X1 \mult_20/S2_22_4  ( .A(\mult_20/ab[22][4] ), .B(
        \mult_20/CARRYB[21][4] ), .CI(\mult_20/SUMB[21][5] ), .CO(
        \mult_20/CARRYB[22][4] ), .S(\mult_20/SUMB[22][4] ) );
  FA_X1 \mult_20/S2_22_3  ( .A(\mult_20/ab[22][3] ), .B(
        \mult_20/CARRYB[21][3] ), .CI(\mult_20/SUMB[21][4] ), .CO(
        \mult_20/CARRYB[22][3] ), .S(\mult_20/SUMB[22][3] ) );
  FA_X1 \mult_20/S2_22_2  ( .A(\mult_20/ab[22][2] ), .B(
        \mult_20/CARRYB[21][2] ), .CI(\mult_20/SUMB[21][3] ), .CO(
        \mult_20/CARRYB[22][2] ), .S(\mult_20/SUMB[22][2] ) );
  FA_X1 \mult_20/S2_22_1  ( .A(\mult_20/ab[22][1] ), .B(
        \mult_20/CARRYB[21][1] ), .CI(\mult_20/SUMB[21][2] ), .CO(
        \mult_20/CARRYB[22][1] ), .S(\mult_20/SUMB[22][1] ) );
  FA_X1 \mult_20/S1_22_0  ( .A(\mult_20/ab[22][0] ), .B(
        \mult_20/CARRYB[21][0] ), .CI(\mult_20/SUMB[21][1] ), .CO(
        \mult_20/CARRYB[22][0] ), .S(N86) );
  FA_X1 \mult_20/S3_23_30  ( .A(\mult_20/ab[23][30] ), .B(
        \mult_20/CARRYB[22][30] ), .CI(\mult_20/ab[22][31] ), .CO(
        \mult_20/CARRYB[23][30] ), .S(\mult_20/SUMB[23][30] ) );
  FA_X1 \mult_20/S2_23_29  ( .A(\mult_20/ab[23][29] ), .B(
        \mult_20/CARRYB[22][29] ), .CI(\mult_20/SUMB[22][30] ), .CO(
        \mult_20/CARRYB[23][29] ), .S(\mult_20/SUMB[23][29] ) );
  FA_X1 \mult_20/S2_23_28  ( .A(\mult_20/ab[23][28] ), .B(
        \mult_20/CARRYB[22][28] ), .CI(\mult_20/SUMB[22][29] ), .CO(
        \mult_20/CARRYB[23][28] ), .S(\mult_20/SUMB[23][28] ) );
  FA_X1 \mult_20/S2_23_27  ( .A(\mult_20/ab[23][27] ), .B(
        \mult_20/CARRYB[22][27] ), .CI(\mult_20/SUMB[22][28] ), .CO(
        \mult_20/CARRYB[23][27] ), .S(\mult_20/SUMB[23][27] ) );
  FA_X1 \mult_20/S2_23_26  ( .A(\mult_20/ab[23][26] ), .B(
        \mult_20/CARRYB[22][26] ), .CI(\mult_20/SUMB[22][27] ), .CO(
        \mult_20/CARRYB[23][26] ), .S(\mult_20/SUMB[23][26] ) );
  FA_X1 \mult_20/S2_23_25  ( .A(\mult_20/ab[23][25] ), .B(
        \mult_20/CARRYB[22][25] ), .CI(\mult_20/SUMB[22][26] ), .CO(
        \mult_20/CARRYB[23][25] ), .S(\mult_20/SUMB[23][25] ) );
  FA_X1 \mult_20/S2_23_24  ( .A(\mult_20/ab[23][24] ), .B(
        \mult_20/CARRYB[22][24] ), .CI(\mult_20/SUMB[22][25] ), .CO(
        \mult_20/CARRYB[23][24] ), .S(\mult_20/SUMB[23][24] ) );
  FA_X1 \mult_20/S2_23_23  ( .A(\mult_20/ab[23][23] ), .B(
        \mult_20/CARRYB[22][23] ), .CI(\mult_20/SUMB[22][24] ), .CO(
        \mult_20/CARRYB[23][23] ), .S(\mult_20/SUMB[23][23] ) );
  FA_X1 \mult_20/S2_23_22  ( .A(\mult_20/ab[23][22] ), .B(
        \mult_20/CARRYB[22][22] ), .CI(\mult_20/SUMB[22][23] ), .CO(
        \mult_20/CARRYB[23][22] ), .S(\mult_20/SUMB[23][22] ) );
  FA_X1 \mult_20/S2_23_21  ( .A(\mult_20/ab[23][21] ), .B(
        \mult_20/CARRYB[22][21] ), .CI(\mult_20/SUMB[22][22] ), .CO(
        \mult_20/CARRYB[23][21] ), .S(\mult_20/SUMB[23][21] ) );
  FA_X1 \mult_20/S2_23_20  ( .A(\mult_20/ab[23][20] ), .B(
        \mult_20/CARRYB[22][20] ), .CI(\mult_20/SUMB[22][21] ), .CO(
        \mult_20/CARRYB[23][20] ), .S(\mult_20/SUMB[23][20] ) );
  FA_X1 \mult_20/S2_23_19  ( .A(\mult_20/ab[23][19] ), .B(
        \mult_20/CARRYB[22][19] ), .CI(\mult_20/SUMB[22][20] ), .CO(
        \mult_20/CARRYB[23][19] ), .S(\mult_20/SUMB[23][19] ) );
  FA_X1 \mult_20/S2_23_18  ( .A(\mult_20/ab[23][18] ), .B(
        \mult_20/CARRYB[22][18] ), .CI(\mult_20/SUMB[22][19] ), .CO(
        \mult_20/CARRYB[23][18] ), .S(\mult_20/SUMB[23][18] ) );
  FA_X1 \mult_20/S2_23_17  ( .A(\mult_20/ab[23][17] ), .B(
        \mult_20/CARRYB[22][17] ), .CI(\mult_20/SUMB[22][18] ), .CO(
        \mult_20/CARRYB[23][17] ), .S(\mult_20/SUMB[23][17] ) );
  FA_X1 \mult_20/S2_23_16  ( .A(\mult_20/ab[23][16] ), .B(
        \mult_20/CARRYB[22][16] ), .CI(\mult_20/SUMB[22][17] ), .CO(
        \mult_20/CARRYB[23][16] ), .S(\mult_20/SUMB[23][16] ) );
  FA_X1 \mult_20/S2_23_15  ( .A(\mult_20/ab[23][15] ), .B(
        \mult_20/CARRYB[22][15] ), .CI(\mult_20/SUMB[22][16] ), .CO(
        \mult_20/CARRYB[23][15] ), .S(\mult_20/SUMB[23][15] ) );
  FA_X1 \mult_20/S2_23_14  ( .A(\mult_20/ab[23][14] ), .B(
        \mult_20/CARRYB[22][14] ), .CI(\mult_20/SUMB[22][15] ), .CO(
        \mult_20/CARRYB[23][14] ), .S(\mult_20/SUMB[23][14] ) );
  FA_X1 \mult_20/S2_23_13  ( .A(\mult_20/ab[23][13] ), .B(
        \mult_20/CARRYB[22][13] ), .CI(\mult_20/SUMB[22][14] ), .CO(
        \mult_20/CARRYB[23][13] ), .S(\mult_20/SUMB[23][13] ) );
  FA_X1 \mult_20/S2_23_12  ( .A(\mult_20/ab[23][12] ), .B(
        \mult_20/CARRYB[22][12] ), .CI(\mult_20/SUMB[22][13] ), .CO(
        \mult_20/CARRYB[23][12] ), .S(\mult_20/SUMB[23][12] ) );
  FA_X1 \mult_20/S2_23_11  ( .A(\mult_20/ab[23][11] ), .B(
        \mult_20/CARRYB[22][11] ), .CI(\mult_20/SUMB[22][12] ), .CO(
        \mult_20/CARRYB[23][11] ), .S(\mult_20/SUMB[23][11] ) );
  FA_X1 \mult_20/S2_23_10  ( .A(\mult_20/ab[23][10] ), .B(
        \mult_20/CARRYB[22][10] ), .CI(\mult_20/SUMB[22][11] ), .CO(
        \mult_20/CARRYB[23][10] ), .S(\mult_20/SUMB[23][10] ) );
  FA_X1 \mult_20/S2_23_9  ( .A(\mult_20/ab[23][9] ), .B(
        \mult_20/CARRYB[22][9] ), .CI(\mult_20/SUMB[22][10] ), .CO(
        \mult_20/CARRYB[23][9] ), .S(\mult_20/SUMB[23][9] ) );
  FA_X1 \mult_20/S2_23_8  ( .A(\mult_20/ab[23][8] ), .B(
        \mult_20/CARRYB[22][8] ), .CI(\mult_20/SUMB[22][9] ), .CO(
        \mult_20/CARRYB[23][8] ), .S(\mult_20/SUMB[23][8] ) );
  FA_X1 \mult_20/S2_23_7  ( .A(\mult_20/ab[23][7] ), .B(
        \mult_20/CARRYB[22][7] ), .CI(\mult_20/SUMB[22][8] ), .CO(
        \mult_20/CARRYB[23][7] ), .S(\mult_20/SUMB[23][7] ) );
  FA_X1 \mult_20/S2_23_6  ( .A(\mult_20/ab[23][6] ), .B(
        \mult_20/CARRYB[22][6] ), .CI(\mult_20/SUMB[22][7] ), .CO(
        \mult_20/CARRYB[23][6] ), .S(\mult_20/SUMB[23][6] ) );
  FA_X1 \mult_20/S2_23_5  ( .A(\mult_20/ab[23][5] ), .B(
        \mult_20/CARRYB[22][5] ), .CI(\mult_20/SUMB[22][6] ), .CO(
        \mult_20/CARRYB[23][5] ), .S(\mult_20/SUMB[23][5] ) );
  FA_X1 \mult_20/S2_23_4  ( .A(\mult_20/ab[23][4] ), .B(
        \mult_20/CARRYB[22][4] ), .CI(\mult_20/SUMB[22][5] ), .CO(
        \mult_20/CARRYB[23][4] ), .S(\mult_20/SUMB[23][4] ) );
  FA_X1 \mult_20/S2_23_3  ( .A(\mult_20/ab[23][3] ), .B(
        \mult_20/CARRYB[22][3] ), .CI(\mult_20/SUMB[22][4] ), .CO(
        \mult_20/CARRYB[23][3] ), .S(\mult_20/SUMB[23][3] ) );
  FA_X1 \mult_20/S2_23_2  ( .A(\mult_20/ab[23][2] ), .B(
        \mult_20/CARRYB[22][2] ), .CI(\mult_20/SUMB[22][3] ), .CO(
        \mult_20/CARRYB[23][2] ), .S(\mult_20/SUMB[23][2] ) );
  FA_X1 \mult_20/S2_23_1  ( .A(\mult_20/ab[23][1] ), .B(
        \mult_20/CARRYB[22][1] ), .CI(\mult_20/SUMB[22][2] ), .CO(
        \mult_20/CARRYB[23][1] ), .S(\mult_20/SUMB[23][1] ) );
  FA_X1 \mult_20/S1_23_0  ( .A(\mult_20/ab[23][0] ), .B(
        \mult_20/CARRYB[22][0] ), .CI(\mult_20/SUMB[22][1] ), .CO(
        \mult_20/CARRYB[23][0] ), .S(N87) );
  FA_X1 \mult_20/S3_24_30  ( .A(\mult_20/ab[24][30] ), .B(
        \mult_20/CARRYB[23][30] ), .CI(\mult_20/ab[23][31] ), .CO(
        \mult_20/CARRYB[24][30] ), .S(\mult_20/SUMB[24][30] ) );
  FA_X1 \mult_20/S2_24_29  ( .A(\mult_20/ab[24][29] ), .B(
        \mult_20/CARRYB[23][29] ), .CI(\mult_20/SUMB[23][30] ), .CO(
        \mult_20/CARRYB[24][29] ), .S(\mult_20/SUMB[24][29] ) );
  FA_X1 \mult_20/S2_24_28  ( .A(\mult_20/ab[24][28] ), .B(
        \mult_20/CARRYB[23][28] ), .CI(\mult_20/SUMB[23][29] ), .CO(
        \mult_20/CARRYB[24][28] ), .S(\mult_20/SUMB[24][28] ) );
  FA_X1 \mult_20/S2_24_27  ( .A(\mult_20/ab[24][27] ), .B(
        \mult_20/CARRYB[23][27] ), .CI(\mult_20/SUMB[23][28] ), .CO(
        \mult_20/CARRYB[24][27] ), .S(\mult_20/SUMB[24][27] ) );
  FA_X1 \mult_20/S2_24_26  ( .A(\mult_20/ab[24][26] ), .B(
        \mult_20/CARRYB[23][26] ), .CI(\mult_20/SUMB[23][27] ), .CO(
        \mult_20/CARRYB[24][26] ), .S(\mult_20/SUMB[24][26] ) );
  FA_X1 \mult_20/S2_24_25  ( .A(\mult_20/ab[24][25] ), .B(
        \mult_20/CARRYB[23][25] ), .CI(\mult_20/SUMB[23][26] ), .CO(
        \mult_20/CARRYB[24][25] ), .S(\mult_20/SUMB[24][25] ) );
  FA_X1 \mult_20/S2_24_24  ( .A(\mult_20/ab[24][24] ), .B(
        \mult_20/CARRYB[23][24] ), .CI(\mult_20/SUMB[23][25] ), .CO(
        \mult_20/CARRYB[24][24] ), .S(\mult_20/SUMB[24][24] ) );
  FA_X1 \mult_20/S2_24_23  ( .A(\mult_20/ab[24][23] ), .B(
        \mult_20/CARRYB[23][23] ), .CI(\mult_20/SUMB[23][24] ), .CO(
        \mult_20/CARRYB[24][23] ), .S(\mult_20/SUMB[24][23] ) );
  FA_X1 \mult_20/S2_24_22  ( .A(\mult_20/ab[24][22] ), .B(
        \mult_20/CARRYB[23][22] ), .CI(\mult_20/SUMB[23][23] ), .CO(
        \mult_20/CARRYB[24][22] ), .S(\mult_20/SUMB[24][22] ) );
  FA_X1 \mult_20/S2_24_21  ( .A(\mult_20/ab[24][21] ), .B(
        \mult_20/CARRYB[23][21] ), .CI(\mult_20/SUMB[23][22] ), .CO(
        \mult_20/CARRYB[24][21] ), .S(\mult_20/SUMB[24][21] ) );
  FA_X1 \mult_20/S2_24_20  ( .A(\mult_20/ab[24][20] ), .B(
        \mult_20/CARRYB[23][20] ), .CI(\mult_20/SUMB[23][21] ), .CO(
        \mult_20/CARRYB[24][20] ), .S(\mult_20/SUMB[24][20] ) );
  FA_X1 \mult_20/S2_24_19  ( .A(\mult_20/ab[24][19] ), .B(
        \mult_20/CARRYB[23][19] ), .CI(\mult_20/SUMB[23][20] ), .CO(
        \mult_20/CARRYB[24][19] ), .S(\mult_20/SUMB[24][19] ) );
  FA_X1 \mult_20/S2_24_18  ( .A(\mult_20/ab[24][18] ), .B(
        \mult_20/CARRYB[23][18] ), .CI(\mult_20/SUMB[23][19] ), .CO(
        \mult_20/CARRYB[24][18] ), .S(\mult_20/SUMB[24][18] ) );
  FA_X1 \mult_20/S2_24_17  ( .A(\mult_20/ab[24][17] ), .B(
        \mult_20/CARRYB[23][17] ), .CI(\mult_20/SUMB[23][18] ), .CO(
        \mult_20/CARRYB[24][17] ), .S(\mult_20/SUMB[24][17] ) );
  FA_X1 \mult_20/S2_24_16  ( .A(\mult_20/ab[24][16] ), .B(
        \mult_20/CARRYB[23][16] ), .CI(\mult_20/SUMB[23][17] ), .CO(
        \mult_20/CARRYB[24][16] ), .S(\mult_20/SUMB[24][16] ) );
  FA_X1 \mult_20/S2_24_15  ( .A(\mult_20/ab[24][15] ), .B(
        \mult_20/CARRYB[23][15] ), .CI(\mult_20/SUMB[23][16] ), .CO(
        \mult_20/CARRYB[24][15] ), .S(\mult_20/SUMB[24][15] ) );
  FA_X1 \mult_20/S2_24_14  ( .A(\mult_20/ab[24][14] ), .B(
        \mult_20/CARRYB[23][14] ), .CI(\mult_20/SUMB[23][15] ), .CO(
        \mult_20/CARRYB[24][14] ), .S(\mult_20/SUMB[24][14] ) );
  FA_X1 \mult_20/S2_24_13  ( .A(\mult_20/ab[24][13] ), .B(
        \mult_20/CARRYB[23][13] ), .CI(\mult_20/SUMB[23][14] ), .CO(
        \mult_20/CARRYB[24][13] ), .S(\mult_20/SUMB[24][13] ) );
  FA_X1 \mult_20/S2_24_12  ( .A(\mult_20/ab[24][12] ), .B(
        \mult_20/CARRYB[23][12] ), .CI(\mult_20/SUMB[23][13] ), .CO(
        \mult_20/CARRYB[24][12] ), .S(\mult_20/SUMB[24][12] ) );
  FA_X1 \mult_20/S2_24_11  ( .A(\mult_20/ab[24][11] ), .B(
        \mult_20/CARRYB[23][11] ), .CI(\mult_20/SUMB[23][12] ), .CO(
        \mult_20/CARRYB[24][11] ), .S(\mult_20/SUMB[24][11] ) );
  FA_X1 \mult_20/S2_24_10  ( .A(\mult_20/ab[24][10] ), .B(
        \mult_20/CARRYB[23][10] ), .CI(\mult_20/SUMB[23][11] ), .CO(
        \mult_20/CARRYB[24][10] ), .S(\mult_20/SUMB[24][10] ) );
  FA_X1 \mult_20/S2_24_9  ( .A(\mult_20/ab[24][9] ), .B(
        \mult_20/CARRYB[23][9] ), .CI(\mult_20/SUMB[23][10] ), .CO(
        \mult_20/CARRYB[24][9] ), .S(\mult_20/SUMB[24][9] ) );
  FA_X1 \mult_20/S2_24_8  ( .A(\mult_20/ab[24][8] ), .B(
        \mult_20/CARRYB[23][8] ), .CI(\mult_20/SUMB[23][9] ), .CO(
        \mult_20/CARRYB[24][8] ), .S(\mult_20/SUMB[24][8] ) );
  FA_X1 \mult_20/S2_24_7  ( .A(\mult_20/ab[24][7] ), .B(
        \mult_20/CARRYB[23][7] ), .CI(\mult_20/SUMB[23][8] ), .CO(
        \mult_20/CARRYB[24][7] ), .S(\mult_20/SUMB[24][7] ) );
  FA_X1 \mult_20/S2_24_6  ( .A(\mult_20/ab[24][6] ), .B(
        \mult_20/CARRYB[23][6] ), .CI(\mult_20/SUMB[23][7] ), .CO(
        \mult_20/CARRYB[24][6] ), .S(\mult_20/SUMB[24][6] ) );
  FA_X1 \mult_20/S2_24_5  ( .A(\mult_20/ab[24][5] ), .B(
        \mult_20/CARRYB[23][5] ), .CI(\mult_20/SUMB[23][6] ), .CO(
        \mult_20/CARRYB[24][5] ), .S(\mult_20/SUMB[24][5] ) );
  FA_X1 \mult_20/S2_24_4  ( .A(\mult_20/ab[24][4] ), .B(
        \mult_20/CARRYB[23][4] ), .CI(\mult_20/SUMB[23][5] ), .CO(
        \mult_20/CARRYB[24][4] ), .S(\mult_20/SUMB[24][4] ) );
  FA_X1 \mult_20/S2_24_3  ( .A(\mult_20/ab[24][3] ), .B(
        \mult_20/CARRYB[23][3] ), .CI(\mult_20/SUMB[23][4] ), .CO(
        \mult_20/CARRYB[24][3] ), .S(\mult_20/SUMB[24][3] ) );
  FA_X1 \mult_20/S2_24_2  ( .A(\mult_20/ab[24][2] ), .B(
        \mult_20/CARRYB[23][2] ), .CI(\mult_20/SUMB[23][3] ), .CO(
        \mult_20/CARRYB[24][2] ), .S(\mult_20/SUMB[24][2] ) );
  FA_X1 \mult_20/S2_24_1  ( .A(\mult_20/ab[24][1] ), .B(
        \mult_20/CARRYB[23][1] ), .CI(\mult_20/SUMB[23][2] ), .CO(
        \mult_20/CARRYB[24][1] ), .S(\mult_20/SUMB[24][1] ) );
  FA_X1 \mult_20/S1_24_0  ( .A(\mult_20/ab[24][0] ), .B(
        \mult_20/CARRYB[23][0] ), .CI(\mult_20/SUMB[23][1] ), .CO(
        \mult_20/CARRYB[24][0] ), .S(N88) );
  FA_X1 \mult_20/S3_25_30  ( .A(\mult_20/ab[25][30] ), .B(
        \mult_20/CARRYB[24][30] ), .CI(\mult_20/ab[24][31] ), .CO(
        \mult_20/CARRYB[25][30] ), .S(\mult_20/SUMB[25][30] ) );
  FA_X1 \mult_20/S2_25_29  ( .A(\mult_20/ab[25][29] ), .B(
        \mult_20/CARRYB[24][29] ), .CI(\mult_20/SUMB[24][30] ), .CO(
        \mult_20/CARRYB[25][29] ), .S(\mult_20/SUMB[25][29] ) );
  FA_X1 \mult_20/S2_25_28  ( .A(\mult_20/ab[25][28] ), .B(
        \mult_20/CARRYB[24][28] ), .CI(\mult_20/SUMB[24][29] ), .CO(
        \mult_20/CARRYB[25][28] ), .S(\mult_20/SUMB[25][28] ) );
  FA_X1 \mult_20/S2_25_27  ( .A(\mult_20/ab[25][27] ), .B(
        \mult_20/CARRYB[24][27] ), .CI(\mult_20/SUMB[24][28] ), .CO(
        \mult_20/CARRYB[25][27] ), .S(\mult_20/SUMB[25][27] ) );
  FA_X1 \mult_20/S2_25_26  ( .A(\mult_20/ab[25][26] ), .B(
        \mult_20/CARRYB[24][26] ), .CI(\mult_20/SUMB[24][27] ), .CO(
        \mult_20/CARRYB[25][26] ), .S(\mult_20/SUMB[25][26] ) );
  FA_X1 \mult_20/S2_25_25  ( .A(\mult_20/ab[25][25] ), .B(
        \mult_20/CARRYB[24][25] ), .CI(\mult_20/SUMB[24][26] ), .CO(
        \mult_20/CARRYB[25][25] ), .S(\mult_20/SUMB[25][25] ) );
  FA_X1 \mult_20/S2_25_24  ( .A(\mult_20/ab[25][24] ), .B(
        \mult_20/CARRYB[24][24] ), .CI(\mult_20/SUMB[24][25] ), .CO(
        \mult_20/CARRYB[25][24] ), .S(\mult_20/SUMB[25][24] ) );
  FA_X1 \mult_20/S2_25_23  ( .A(\mult_20/ab[25][23] ), .B(
        \mult_20/CARRYB[24][23] ), .CI(\mult_20/SUMB[24][24] ), .CO(
        \mult_20/CARRYB[25][23] ), .S(\mult_20/SUMB[25][23] ) );
  FA_X1 \mult_20/S2_25_22  ( .A(\mult_20/ab[25][22] ), .B(
        \mult_20/CARRYB[24][22] ), .CI(\mult_20/SUMB[24][23] ), .CO(
        \mult_20/CARRYB[25][22] ), .S(\mult_20/SUMB[25][22] ) );
  FA_X1 \mult_20/S2_25_21  ( .A(\mult_20/ab[25][21] ), .B(
        \mult_20/CARRYB[24][21] ), .CI(\mult_20/SUMB[24][22] ), .CO(
        \mult_20/CARRYB[25][21] ), .S(\mult_20/SUMB[25][21] ) );
  FA_X1 \mult_20/S2_25_20  ( .A(\mult_20/ab[25][20] ), .B(
        \mult_20/CARRYB[24][20] ), .CI(\mult_20/SUMB[24][21] ), .CO(
        \mult_20/CARRYB[25][20] ), .S(\mult_20/SUMB[25][20] ) );
  FA_X1 \mult_20/S2_25_19  ( .A(\mult_20/ab[25][19] ), .B(
        \mult_20/CARRYB[24][19] ), .CI(\mult_20/SUMB[24][20] ), .CO(
        \mult_20/CARRYB[25][19] ), .S(\mult_20/SUMB[25][19] ) );
  FA_X1 \mult_20/S2_25_18  ( .A(\mult_20/ab[25][18] ), .B(
        \mult_20/CARRYB[24][18] ), .CI(\mult_20/SUMB[24][19] ), .CO(
        \mult_20/CARRYB[25][18] ), .S(\mult_20/SUMB[25][18] ) );
  FA_X1 \mult_20/S2_25_17  ( .A(\mult_20/ab[25][17] ), .B(
        \mult_20/CARRYB[24][17] ), .CI(\mult_20/SUMB[24][18] ), .CO(
        \mult_20/CARRYB[25][17] ), .S(\mult_20/SUMB[25][17] ) );
  FA_X1 \mult_20/S2_25_16  ( .A(\mult_20/ab[25][16] ), .B(
        \mult_20/CARRYB[24][16] ), .CI(\mult_20/SUMB[24][17] ), .CO(
        \mult_20/CARRYB[25][16] ), .S(\mult_20/SUMB[25][16] ) );
  FA_X1 \mult_20/S2_25_15  ( .A(\mult_20/ab[25][15] ), .B(
        \mult_20/CARRYB[24][15] ), .CI(\mult_20/SUMB[24][16] ), .CO(
        \mult_20/CARRYB[25][15] ), .S(\mult_20/SUMB[25][15] ) );
  FA_X1 \mult_20/S2_25_14  ( .A(\mult_20/ab[25][14] ), .B(
        \mult_20/CARRYB[24][14] ), .CI(\mult_20/SUMB[24][15] ), .CO(
        \mult_20/CARRYB[25][14] ), .S(\mult_20/SUMB[25][14] ) );
  FA_X1 \mult_20/S2_25_13  ( .A(\mult_20/ab[25][13] ), .B(
        \mult_20/CARRYB[24][13] ), .CI(\mult_20/SUMB[24][14] ), .CO(
        \mult_20/CARRYB[25][13] ), .S(\mult_20/SUMB[25][13] ) );
  FA_X1 \mult_20/S2_25_12  ( .A(\mult_20/ab[25][12] ), .B(
        \mult_20/CARRYB[24][12] ), .CI(\mult_20/SUMB[24][13] ), .CO(
        \mult_20/CARRYB[25][12] ), .S(\mult_20/SUMB[25][12] ) );
  FA_X1 \mult_20/S2_25_11  ( .A(\mult_20/ab[25][11] ), .B(
        \mult_20/CARRYB[24][11] ), .CI(\mult_20/SUMB[24][12] ), .CO(
        \mult_20/CARRYB[25][11] ), .S(\mult_20/SUMB[25][11] ) );
  FA_X1 \mult_20/S2_25_10  ( .A(\mult_20/ab[25][10] ), .B(
        \mult_20/CARRYB[24][10] ), .CI(\mult_20/SUMB[24][11] ), .CO(
        \mult_20/CARRYB[25][10] ), .S(\mult_20/SUMB[25][10] ) );
  FA_X1 \mult_20/S2_25_9  ( .A(\mult_20/ab[25][9] ), .B(
        \mult_20/CARRYB[24][9] ), .CI(\mult_20/SUMB[24][10] ), .CO(
        \mult_20/CARRYB[25][9] ), .S(\mult_20/SUMB[25][9] ) );
  FA_X1 \mult_20/S2_25_8  ( .A(\mult_20/ab[25][8] ), .B(
        \mult_20/CARRYB[24][8] ), .CI(\mult_20/SUMB[24][9] ), .CO(
        \mult_20/CARRYB[25][8] ), .S(\mult_20/SUMB[25][8] ) );
  FA_X1 \mult_20/S2_25_7  ( .A(\mult_20/ab[25][7] ), .B(
        \mult_20/CARRYB[24][7] ), .CI(\mult_20/SUMB[24][8] ), .CO(
        \mult_20/CARRYB[25][7] ), .S(\mult_20/SUMB[25][7] ) );
  FA_X1 \mult_20/S2_25_6  ( .A(\mult_20/ab[25][6] ), .B(
        \mult_20/CARRYB[24][6] ), .CI(\mult_20/SUMB[24][7] ), .CO(
        \mult_20/CARRYB[25][6] ), .S(\mult_20/SUMB[25][6] ) );
  FA_X1 \mult_20/S2_25_5  ( .A(\mult_20/ab[25][5] ), .B(
        \mult_20/CARRYB[24][5] ), .CI(\mult_20/SUMB[24][6] ), .CO(
        \mult_20/CARRYB[25][5] ), .S(\mult_20/SUMB[25][5] ) );
  FA_X1 \mult_20/S2_25_4  ( .A(\mult_20/ab[25][4] ), .B(
        \mult_20/CARRYB[24][4] ), .CI(\mult_20/SUMB[24][5] ), .CO(
        \mult_20/CARRYB[25][4] ), .S(\mult_20/SUMB[25][4] ) );
  FA_X1 \mult_20/S2_25_3  ( .A(\mult_20/ab[25][3] ), .B(
        \mult_20/CARRYB[24][3] ), .CI(\mult_20/SUMB[24][4] ), .CO(
        \mult_20/CARRYB[25][3] ), .S(\mult_20/SUMB[25][3] ) );
  FA_X1 \mult_20/S2_25_2  ( .A(\mult_20/ab[25][2] ), .B(
        \mult_20/CARRYB[24][2] ), .CI(\mult_20/SUMB[24][3] ), .CO(
        \mult_20/CARRYB[25][2] ), .S(\mult_20/SUMB[25][2] ) );
  FA_X1 \mult_20/S2_25_1  ( .A(\mult_20/ab[25][1] ), .B(
        \mult_20/CARRYB[24][1] ), .CI(\mult_20/SUMB[24][2] ), .CO(
        \mult_20/CARRYB[25][1] ), .S(\mult_20/SUMB[25][1] ) );
  FA_X1 \mult_20/S1_25_0  ( .A(\mult_20/ab[25][0] ), .B(
        \mult_20/CARRYB[24][0] ), .CI(\mult_20/SUMB[24][1] ), .CO(
        \mult_20/CARRYB[25][0] ), .S(N89) );
  FA_X1 \mult_20/S3_26_30  ( .A(\mult_20/ab[26][30] ), .B(
        \mult_20/CARRYB[25][30] ), .CI(\mult_20/ab[25][31] ), .CO(
        \mult_20/CARRYB[26][30] ), .S(\mult_20/SUMB[26][30] ) );
  FA_X1 \mult_20/S2_26_29  ( .A(\mult_20/ab[26][29] ), .B(
        \mult_20/CARRYB[25][29] ), .CI(\mult_20/SUMB[25][30] ), .CO(
        \mult_20/CARRYB[26][29] ), .S(\mult_20/SUMB[26][29] ) );
  FA_X1 \mult_20/S2_26_28  ( .A(\mult_20/ab[26][28] ), .B(
        \mult_20/CARRYB[25][28] ), .CI(\mult_20/SUMB[25][29] ), .CO(
        \mult_20/CARRYB[26][28] ), .S(\mult_20/SUMB[26][28] ) );
  FA_X1 \mult_20/S2_26_27  ( .A(\mult_20/ab[26][27] ), .B(
        \mult_20/CARRYB[25][27] ), .CI(\mult_20/SUMB[25][28] ), .CO(
        \mult_20/CARRYB[26][27] ), .S(\mult_20/SUMB[26][27] ) );
  FA_X1 \mult_20/S2_26_26  ( .A(\mult_20/ab[26][26] ), .B(
        \mult_20/CARRYB[25][26] ), .CI(\mult_20/SUMB[25][27] ), .CO(
        \mult_20/CARRYB[26][26] ), .S(\mult_20/SUMB[26][26] ) );
  FA_X1 \mult_20/S2_26_25  ( .A(\mult_20/ab[26][25] ), .B(
        \mult_20/CARRYB[25][25] ), .CI(\mult_20/SUMB[25][26] ), .CO(
        \mult_20/CARRYB[26][25] ), .S(\mult_20/SUMB[26][25] ) );
  FA_X1 \mult_20/S2_26_24  ( .A(\mult_20/ab[26][24] ), .B(
        \mult_20/CARRYB[25][24] ), .CI(\mult_20/SUMB[25][25] ), .CO(
        \mult_20/CARRYB[26][24] ), .S(\mult_20/SUMB[26][24] ) );
  FA_X1 \mult_20/S2_26_23  ( .A(\mult_20/ab[26][23] ), .B(
        \mult_20/CARRYB[25][23] ), .CI(\mult_20/SUMB[25][24] ), .CO(
        \mult_20/CARRYB[26][23] ), .S(\mult_20/SUMB[26][23] ) );
  FA_X1 \mult_20/S2_26_22  ( .A(\mult_20/ab[26][22] ), .B(
        \mult_20/CARRYB[25][22] ), .CI(\mult_20/SUMB[25][23] ), .CO(
        \mult_20/CARRYB[26][22] ), .S(\mult_20/SUMB[26][22] ) );
  FA_X1 \mult_20/S2_26_21  ( .A(\mult_20/ab[26][21] ), .B(
        \mult_20/CARRYB[25][21] ), .CI(\mult_20/SUMB[25][22] ), .CO(
        \mult_20/CARRYB[26][21] ), .S(\mult_20/SUMB[26][21] ) );
  FA_X1 \mult_20/S2_26_20  ( .A(\mult_20/ab[26][20] ), .B(
        \mult_20/CARRYB[25][20] ), .CI(\mult_20/SUMB[25][21] ), .CO(
        \mult_20/CARRYB[26][20] ), .S(\mult_20/SUMB[26][20] ) );
  FA_X1 \mult_20/S2_26_19  ( .A(\mult_20/ab[26][19] ), .B(
        \mult_20/CARRYB[25][19] ), .CI(\mult_20/SUMB[25][20] ), .CO(
        \mult_20/CARRYB[26][19] ), .S(\mult_20/SUMB[26][19] ) );
  FA_X1 \mult_20/S2_26_18  ( .A(\mult_20/ab[26][18] ), .B(
        \mult_20/CARRYB[25][18] ), .CI(\mult_20/SUMB[25][19] ), .CO(
        \mult_20/CARRYB[26][18] ), .S(\mult_20/SUMB[26][18] ) );
  FA_X1 \mult_20/S2_26_17  ( .A(\mult_20/ab[26][17] ), .B(
        \mult_20/CARRYB[25][17] ), .CI(\mult_20/SUMB[25][18] ), .CO(
        \mult_20/CARRYB[26][17] ), .S(\mult_20/SUMB[26][17] ) );
  FA_X1 \mult_20/S2_26_16  ( .A(\mult_20/ab[26][16] ), .B(
        \mult_20/CARRYB[25][16] ), .CI(\mult_20/SUMB[25][17] ), .CO(
        \mult_20/CARRYB[26][16] ), .S(\mult_20/SUMB[26][16] ) );
  FA_X1 \mult_20/S2_26_15  ( .A(\mult_20/ab[26][15] ), .B(
        \mult_20/CARRYB[25][15] ), .CI(\mult_20/SUMB[25][16] ), .CO(
        \mult_20/CARRYB[26][15] ), .S(\mult_20/SUMB[26][15] ) );
  FA_X1 \mult_20/S2_26_14  ( .A(\mult_20/ab[26][14] ), .B(
        \mult_20/CARRYB[25][14] ), .CI(\mult_20/SUMB[25][15] ), .CO(
        \mult_20/CARRYB[26][14] ), .S(\mult_20/SUMB[26][14] ) );
  FA_X1 \mult_20/S2_26_13  ( .A(\mult_20/ab[26][13] ), .B(
        \mult_20/CARRYB[25][13] ), .CI(\mult_20/SUMB[25][14] ), .CO(
        \mult_20/CARRYB[26][13] ), .S(\mult_20/SUMB[26][13] ) );
  FA_X1 \mult_20/S2_26_12  ( .A(\mult_20/ab[26][12] ), .B(
        \mult_20/CARRYB[25][12] ), .CI(\mult_20/SUMB[25][13] ), .CO(
        \mult_20/CARRYB[26][12] ), .S(\mult_20/SUMB[26][12] ) );
  FA_X1 \mult_20/S2_26_11  ( .A(\mult_20/ab[26][11] ), .B(
        \mult_20/CARRYB[25][11] ), .CI(\mult_20/SUMB[25][12] ), .CO(
        \mult_20/CARRYB[26][11] ), .S(\mult_20/SUMB[26][11] ) );
  FA_X1 \mult_20/S2_26_10  ( .A(\mult_20/ab[26][10] ), .B(
        \mult_20/CARRYB[25][10] ), .CI(\mult_20/SUMB[25][11] ), .CO(
        \mult_20/CARRYB[26][10] ), .S(\mult_20/SUMB[26][10] ) );
  FA_X1 \mult_20/S2_26_9  ( .A(\mult_20/ab[26][9] ), .B(
        \mult_20/CARRYB[25][9] ), .CI(\mult_20/SUMB[25][10] ), .CO(
        \mult_20/CARRYB[26][9] ), .S(\mult_20/SUMB[26][9] ) );
  FA_X1 \mult_20/S2_26_8  ( .A(\mult_20/ab[26][8] ), .B(
        \mult_20/CARRYB[25][8] ), .CI(\mult_20/SUMB[25][9] ), .CO(
        \mult_20/CARRYB[26][8] ), .S(\mult_20/SUMB[26][8] ) );
  FA_X1 \mult_20/S2_26_7  ( .A(\mult_20/ab[26][7] ), .B(
        \mult_20/CARRYB[25][7] ), .CI(\mult_20/SUMB[25][8] ), .CO(
        \mult_20/CARRYB[26][7] ), .S(\mult_20/SUMB[26][7] ) );
  FA_X1 \mult_20/S2_26_6  ( .A(\mult_20/ab[26][6] ), .B(
        \mult_20/CARRYB[25][6] ), .CI(\mult_20/SUMB[25][7] ), .CO(
        \mult_20/CARRYB[26][6] ), .S(\mult_20/SUMB[26][6] ) );
  FA_X1 \mult_20/S2_26_5  ( .A(\mult_20/ab[26][5] ), .B(
        \mult_20/CARRYB[25][5] ), .CI(\mult_20/SUMB[25][6] ), .CO(
        \mult_20/CARRYB[26][5] ), .S(\mult_20/SUMB[26][5] ) );
  FA_X1 \mult_20/S2_26_4  ( .A(\mult_20/ab[26][4] ), .B(
        \mult_20/CARRYB[25][4] ), .CI(\mult_20/SUMB[25][5] ), .CO(
        \mult_20/CARRYB[26][4] ), .S(\mult_20/SUMB[26][4] ) );
  FA_X1 \mult_20/S2_26_3  ( .A(\mult_20/ab[26][3] ), .B(
        \mult_20/CARRYB[25][3] ), .CI(\mult_20/SUMB[25][4] ), .CO(
        \mult_20/CARRYB[26][3] ), .S(\mult_20/SUMB[26][3] ) );
  FA_X1 \mult_20/S2_26_2  ( .A(\mult_20/ab[26][2] ), .B(
        \mult_20/CARRYB[25][2] ), .CI(\mult_20/SUMB[25][3] ), .CO(
        \mult_20/CARRYB[26][2] ), .S(\mult_20/SUMB[26][2] ) );
  FA_X1 \mult_20/S2_26_1  ( .A(\mult_20/ab[26][1] ), .B(
        \mult_20/CARRYB[25][1] ), .CI(\mult_20/SUMB[25][2] ), .CO(
        \mult_20/CARRYB[26][1] ), .S(\mult_20/SUMB[26][1] ) );
  FA_X1 \mult_20/S1_26_0  ( .A(\mult_20/ab[26][0] ), .B(
        \mult_20/CARRYB[25][0] ), .CI(\mult_20/SUMB[25][1] ), .CO(
        \mult_20/CARRYB[26][0] ), .S(N90) );
  FA_X1 \mult_20/S3_27_30  ( .A(\mult_20/ab[27][30] ), .B(
        \mult_20/CARRYB[26][30] ), .CI(\mult_20/ab[26][31] ), .CO(
        \mult_20/CARRYB[27][30] ), .S(\mult_20/SUMB[27][30] ) );
  FA_X1 \mult_20/S2_27_29  ( .A(\mult_20/ab[27][29] ), .B(
        \mult_20/CARRYB[26][29] ), .CI(\mult_20/SUMB[26][30] ), .CO(
        \mult_20/CARRYB[27][29] ), .S(\mult_20/SUMB[27][29] ) );
  FA_X1 \mult_20/S2_27_28  ( .A(\mult_20/ab[27][28] ), .B(
        \mult_20/CARRYB[26][28] ), .CI(\mult_20/SUMB[26][29] ), .CO(
        \mult_20/CARRYB[27][28] ), .S(\mult_20/SUMB[27][28] ) );
  FA_X1 \mult_20/S2_27_27  ( .A(\mult_20/ab[27][27] ), .B(
        \mult_20/CARRYB[26][27] ), .CI(\mult_20/SUMB[26][28] ), .CO(
        \mult_20/CARRYB[27][27] ), .S(\mult_20/SUMB[27][27] ) );
  FA_X1 \mult_20/S2_27_26  ( .A(\mult_20/ab[27][26] ), .B(
        \mult_20/CARRYB[26][26] ), .CI(\mult_20/SUMB[26][27] ), .CO(
        \mult_20/CARRYB[27][26] ), .S(\mult_20/SUMB[27][26] ) );
  FA_X1 \mult_20/S2_27_25  ( .A(\mult_20/ab[27][25] ), .B(
        \mult_20/CARRYB[26][25] ), .CI(\mult_20/SUMB[26][26] ), .CO(
        \mult_20/CARRYB[27][25] ), .S(\mult_20/SUMB[27][25] ) );
  FA_X1 \mult_20/S2_27_24  ( .A(\mult_20/ab[27][24] ), .B(
        \mult_20/CARRYB[26][24] ), .CI(\mult_20/SUMB[26][25] ), .CO(
        \mult_20/CARRYB[27][24] ), .S(\mult_20/SUMB[27][24] ) );
  FA_X1 \mult_20/S2_27_23  ( .A(\mult_20/ab[27][23] ), .B(
        \mult_20/CARRYB[26][23] ), .CI(\mult_20/SUMB[26][24] ), .CO(
        \mult_20/CARRYB[27][23] ), .S(\mult_20/SUMB[27][23] ) );
  FA_X1 \mult_20/S2_27_22  ( .A(\mult_20/ab[27][22] ), .B(
        \mult_20/CARRYB[26][22] ), .CI(\mult_20/SUMB[26][23] ), .CO(
        \mult_20/CARRYB[27][22] ), .S(\mult_20/SUMB[27][22] ) );
  FA_X1 \mult_20/S2_27_21  ( .A(\mult_20/ab[27][21] ), .B(
        \mult_20/CARRYB[26][21] ), .CI(\mult_20/SUMB[26][22] ), .CO(
        \mult_20/CARRYB[27][21] ), .S(\mult_20/SUMB[27][21] ) );
  FA_X1 \mult_20/S2_27_20  ( .A(\mult_20/ab[27][20] ), .B(
        \mult_20/CARRYB[26][20] ), .CI(\mult_20/SUMB[26][21] ), .CO(
        \mult_20/CARRYB[27][20] ), .S(\mult_20/SUMB[27][20] ) );
  FA_X1 \mult_20/S2_27_19  ( .A(\mult_20/ab[27][19] ), .B(
        \mult_20/CARRYB[26][19] ), .CI(\mult_20/SUMB[26][20] ), .CO(
        \mult_20/CARRYB[27][19] ), .S(\mult_20/SUMB[27][19] ) );
  FA_X1 \mult_20/S2_27_18  ( .A(\mult_20/ab[27][18] ), .B(
        \mult_20/CARRYB[26][18] ), .CI(\mult_20/SUMB[26][19] ), .CO(
        \mult_20/CARRYB[27][18] ), .S(\mult_20/SUMB[27][18] ) );
  FA_X1 \mult_20/S2_27_17  ( .A(\mult_20/ab[27][17] ), .B(
        \mult_20/CARRYB[26][17] ), .CI(\mult_20/SUMB[26][18] ), .CO(
        \mult_20/CARRYB[27][17] ), .S(\mult_20/SUMB[27][17] ) );
  FA_X1 \mult_20/S2_27_16  ( .A(\mult_20/ab[27][16] ), .B(
        \mult_20/CARRYB[26][16] ), .CI(\mult_20/SUMB[26][17] ), .CO(
        \mult_20/CARRYB[27][16] ), .S(\mult_20/SUMB[27][16] ) );
  FA_X1 \mult_20/S2_27_15  ( .A(\mult_20/ab[27][15] ), .B(
        \mult_20/CARRYB[26][15] ), .CI(\mult_20/SUMB[26][16] ), .CO(
        \mult_20/CARRYB[27][15] ), .S(\mult_20/SUMB[27][15] ) );
  FA_X1 \mult_20/S2_27_14  ( .A(\mult_20/ab[27][14] ), .B(
        \mult_20/CARRYB[26][14] ), .CI(\mult_20/SUMB[26][15] ), .CO(
        \mult_20/CARRYB[27][14] ), .S(\mult_20/SUMB[27][14] ) );
  FA_X1 \mult_20/S2_27_13  ( .A(\mult_20/ab[27][13] ), .B(
        \mult_20/CARRYB[26][13] ), .CI(\mult_20/SUMB[26][14] ), .CO(
        \mult_20/CARRYB[27][13] ), .S(\mult_20/SUMB[27][13] ) );
  FA_X1 \mult_20/S2_27_12  ( .A(\mult_20/ab[27][12] ), .B(
        \mult_20/CARRYB[26][12] ), .CI(\mult_20/SUMB[26][13] ), .CO(
        \mult_20/CARRYB[27][12] ), .S(\mult_20/SUMB[27][12] ) );
  FA_X1 \mult_20/S2_27_11  ( .A(\mult_20/ab[27][11] ), .B(
        \mult_20/CARRYB[26][11] ), .CI(\mult_20/SUMB[26][12] ), .CO(
        \mult_20/CARRYB[27][11] ), .S(\mult_20/SUMB[27][11] ) );
  FA_X1 \mult_20/S2_27_10  ( .A(\mult_20/ab[27][10] ), .B(
        \mult_20/CARRYB[26][10] ), .CI(\mult_20/SUMB[26][11] ), .CO(
        \mult_20/CARRYB[27][10] ), .S(\mult_20/SUMB[27][10] ) );
  FA_X1 \mult_20/S2_27_9  ( .A(\mult_20/ab[27][9] ), .B(
        \mult_20/CARRYB[26][9] ), .CI(\mult_20/SUMB[26][10] ), .CO(
        \mult_20/CARRYB[27][9] ), .S(\mult_20/SUMB[27][9] ) );
  FA_X1 \mult_20/S2_27_8  ( .A(\mult_20/ab[27][8] ), .B(
        \mult_20/CARRYB[26][8] ), .CI(\mult_20/SUMB[26][9] ), .CO(
        \mult_20/CARRYB[27][8] ), .S(\mult_20/SUMB[27][8] ) );
  FA_X1 \mult_20/S2_27_7  ( .A(\mult_20/ab[27][7] ), .B(
        \mult_20/CARRYB[26][7] ), .CI(\mult_20/SUMB[26][8] ), .CO(
        \mult_20/CARRYB[27][7] ), .S(\mult_20/SUMB[27][7] ) );
  FA_X1 \mult_20/S2_27_6  ( .A(\mult_20/ab[27][6] ), .B(
        \mult_20/CARRYB[26][6] ), .CI(\mult_20/SUMB[26][7] ), .CO(
        \mult_20/CARRYB[27][6] ), .S(\mult_20/SUMB[27][6] ) );
  FA_X1 \mult_20/S2_27_5  ( .A(\mult_20/ab[27][5] ), .B(
        \mult_20/CARRYB[26][5] ), .CI(\mult_20/SUMB[26][6] ), .CO(
        \mult_20/CARRYB[27][5] ), .S(\mult_20/SUMB[27][5] ) );
  FA_X1 \mult_20/S2_27_4  ( .A(\mult_20/ab[27][4] ), .B(
        \mult_20/CARRYB[26][4] ), .CI(\mult_20/SUMB[26][5] ), .CO(
        \mult_20/CARRYB[27][4] ), .S(\mult_20/SUMB[27][4] ) );
  FA_X1 \mult_20/S2_27_3  ( .A(\mult_20/ab[27][3] ), .B(
        \mult_20/CARRYB[26][3] ), .CI(\mult_20/SUMB[26][4] ), .CO(
        \mult_20/CARRYB[27][3] ), .S(\mult_20/SUMB[27][3] ) );
  FA_X1 \mult_20/S2_27_2  ( .A(\mult_20/ab[27][2] ), .B(
        \mult_20/CARRYB[26][2] ), .CI(\mult_20/SUMB[26][3] ), .CO(
        \mult_20/CARRYB[27][2] ), .S(\mult_20/SUMB[27][2] ) );
  FA_X1 \mult_20/S2_27_1  ( .A(\mult_20/ab[27][1] ), .B(
        \mult_20/CARRYB[26][1] ), .CI(\mult_20/SUMB[26][2] ), .CO(
        \mult_20/CARRYB[27][1] ), .S(\mult_20/SUMB[27][1] ) );
  FA_X1 \mult_20/S1_27_0  ( .A(\mult_20/ab[27][0] ), .B(
        \mult_20/CARRYB[26][0] ), .CI(\mult_20/SUMB[26][1] ), .CO(
        \mult_20/CARRYB[27][0] ), .S(N91) );
  FA_X1 \mult_20/S3_28_30  ( .A(\mult_20/ab[28][30] ), .B(
        \mult_20/CARRYB[27][30] ), .CI(\mult_20/ab[27][31] ), .CO(
        \mult_20/CARRYB[28][30] ), .S(\mult_20/SUMB[28][30] ) );
  FA_X1 \mult_20/S2_28_29  ( .A(\mult_20/ab[28][29] ), .B(
        \mult_20/CARRYB[27][29] ), .CI(\mult_20/SUMB[27][30] ), .CO(
        \mult_20/CARRYB[28][29] ), .S(\mult_20/SUMB[28][29] ) );
  FA_X1 \mult_20/S2_28_28  ( .A(\mult_20/ab[28][28] ), .B(
        \mult_20/CARRYB[27][28] ), .CI(\mult_20/SUMB[27][29] ), .CO(
        \mult_20/CARRYB[28][28] ), .S(\mult_20/SUMB[28][28] ) );
  FA_X1 \mult_20/S2_28_27  ( .A(\mult_20/ab[28][27] ), .B(
        \mult_20/CARRYB[27][27] ), .CI(\mult_20/SUMB[27][28] ), .CO(
        \mult_20/CARRYB[28][27] ), .S(\mult_20/SUMB[28][27] ) );
  FA_X1 \mult_20/S2_28_26  ( .A(\mult_20/ab[28][26] ), .B(
        \mult_20/CARRYB[27][26] ), .CI(\mult_20/SUMB[27][27] ), .CO(
        \mult_20/CARRYB[28][26] ), .S(\mult_20/SUMB[28][26] ) );
  FA_X1 \mult_20/S2_28_25  ( .A(\mult_20/ab[28][25] ), .B(
        \mult_20/CARRYB[27][25] ), .CI(\mult_20/SUMB[27][26] ), .CO(
        \mult_20/CARRYB[28][25] ), .S(\mult_20/SUMB[28][25] ) );
  FA_X1 \mult_20/S2_28_24  ( .A(\mult_20/ab[28][24] ), .B(
        \mult_20/CARRYB[27][24] ), .CI(\mult_20/SUMB[27][25] ), .CO(
        \mult_20/CARRYB[28][24] ), .S(\mult_20/SUMB[28][24] ) );
  FA_X1 \mult_20/S2_28_23  ( .A(\mult_20/ab[28][23] ), .B(
        \mult_20/CARRYB[27][23] ), .CI(\mult_20/SUMB[27][24] ), .CO(
        \mult_20/CARRYB[28][23] ), .S(\mult_20/SUMB[28][23] ) );
  FA_X1 \mult_20/S2_28_22  ( .A(\mult_20/ab[28][22] ), .B(
        \mult_20/CARRYB[27][22] ), .CI(\mult_20/SUMB[27][23] ), .CO(
        \mult_20/CARRYB[28][22] ), .S(\mult_20/SUMB[28][22] ) );
  FA_X1 \mult_20/S2_28_21  ( .A(\mult_20/ab[28][21] ), .B(
        \mult_20/CARRYB[27][21] ), .CI(\mult_20/SUMB[27][22] ), .CO(
        \mult_20/CARRYB[28][21] ), .S(\mult_20/SUMB[28][21] ) );
  FA_X1 \mult_20/S2_28_20  ( .A(\mult_20/ab[28][20] ), .B(
        \mult_20/CARRYB[27][20] ), .CI(\mult_20/SUMB[27][21] ), .CO(
        \mult_20/CARRYB[28][20] ), .S(\mult_20/SUMB[28][20] ) );
  FA_X1 \mult_20/S2_28_19  ( .A(\mult_20/ab[28][19] ), .B(
        \mult_20/CARRYB[27][19] ), .CI(\mult_20/SUMB[27][20] ), .CO(
        \mult_20/CARRYB[28][19] ), .S(\mult_20/SUMB[28][19] ) );
  FA_X1 \mult_20/S2_28_18  ( .A(\mult_20/ab[28][18] ), .B(
        \mult_20/CARRYB[27][18] ), .CI(\mult_20/SUMB[27][19] ), .CO(
        \mult_20/CARRYB[28][18] ), .S(\mult_20/SUMB[28][18] ) );
  FA_X1 \mult_20/S2_28_17  ( .A(\mult_20/ab[28][17] ), .B(
        \mult_20/CARRYB[27][17] ), .CI(\mult_20/SUMB[27][18] ), .CO(
        \mult_20/CARRYB[28][17] ), .S(\mult_20/SUMB[28][17] ) );
  FA_X1 \mult_20/S2_28_16  ( .A(\mult_20/ab[28][16] ), .B(
        \mult_20/CARRYB[27][16] ), .CI(\mult_20/SUMB[27][17] ), .CO(
        \mult_20/CARRYB[28][16] ), .S(\mult_20/SUMB[28][16] ) );
  FA_X1 \mult_20/S2_28_15  ( .A(\mult_20/ab[28][15] ), .B(
        \mult_20/CARRYB[27][15] ), .CI(\mult_20/SUMB[27][16] ), .CO(
        \mult_20/CARRYB[28][15] ), .S(\mult_20/SUMB[28][15] ) );
  FA_X1 \mult_20/S2_28_14  ( .A(\mult_20/ab[28][14] ), .B(
        \mult_20/CARRYB[27][14] ), .CI(\mult_20/SUMB[27][15] ), .CO(
        \mult_20/CARRYB[28][14] ), .S(\mult_20/SUMB[28][14] ) );
  FA_X1 \mult_20/S2_28_13  ( .A(\mult_20/ab[28][13] ), .B(
        \mult_20/CARRYB[27][13] ), .CI(\mult_20/SUMB[27][14] ), .CO(
        \mult_20/CARRYB[28][13] ), .S(\mult_20/SUMB[28][13] ) );
  FA_X1 \mult_20/S2_28_12  ( .A(\mult_20/ab[28][12] ), .B(
        \mult_20/CARRYB[27][12] ), .CI(\mult_20/SUMB[27][13] ), .CO(
        \mult_20/CARRYB[28][12] ), .S(\mult_20/SUMB[28][12] ) );
  FA_X1 \mult_20/S2_28_11  ( .A(\mult_20/ab[28][11] ), .B(
        \mult_20/CARRYB[27][11] ), .CI(\mult_20/SUMB[27][12] ), .CO(
        \mult_20/CARRYB[28][11] ), .S(\mult_20/SUMB[28][11] ) );
  FA_X1 \mult_20/S2_28_10  ( .A(\mult_20/ab[28][10] ), .B(
        \mult_20/CARRYB[27][10] ), .CI(\mult_20/SUMB[27][11] ), .CO(
        \mult_20/CARRYB[28][10] ), .S(\mult_20/SUMB[28][10] ) );
  FA_X1 \mult_20/S2_28_9  ( .A(\mult_20/ab[28][9] ), .B(
        \mult_20/CARRYB[27][9] ), .CI(\mult_20/SUMB[27][10] ), .CO(
        \mult_20/CARRYB[28][9] ), .S(\mult_20/SUMB[28][9] ) );
  FA_X1 \mult_20/S2_28_8  ( .A(\mult_20/ab[28][8] ), .B(
        \mult_20/CARRYB[27][8] ), .CI(\mult_20/SUMB[27][9] ), .CO(
        \mult_20/CARRYB[28][8] ), .S(\mult_20/SUMB[28][8] ) );
  FA_X1 \mult_20/S2_28_7  ( .A(\mult_20/ab[28][7] ), .B(
        \mult_20/CARRYB[27][7] ), .CI(\mult_20/SUMB[27][8] ), .CO(
        \mult_20/CARRYB[28][7] ), .S(\mult_20/SUMB[28][7] ) );
  FA_X1 \mult_20/S2_28_6  ( .A(\mult_20/ab[28][6] ), .B(
        \mult_20/CARRYB[27][6] ), .CI(\mult_20/SUMB[27][7] ), .CO(
        \mult_20/CARRYB[28][6] ), .S(\mult_20/SUMB[28][6] ) );
  FA_X1 \mult_20/S2_28_5  ( .A(\mult_20/ab[28][5] ), .B(
        \mult_20/CARRYB[27][5] ), .CI(\mult_20/SUMB[27][6] ), .CO(
        \mult_20/CARRYB[28][5] ), .S(\mult_20/SUMB[28][5] ) );
  FA_X1 \mult_20/S2_28_4  ( .A(\mult_20/ab[28][4] ), .B(
        \mult_20/CARRYB[27][4] ), .CI(\mult_20/SUMB[27][5] ), .CO(
        \mult_20/CARRYB[28][4] ), .S(\mult_20/SUMB[28][4] ) );
  FA_X1 \mult_20/S2_28_3  ( .A(\mult_20/ab[28][3] ), .B(
        \mult_20/CARRYB[27][3] ), .CI(\mult_20/SUMB[27][4] ), .CO(
        \mult_20/CARRYB[28][3] ), .S(\mult_20/SUMB[28][3] ) );
  FA_X1 \mult_20/S2_28_2  ( .A(\mult_20/ab[28][2] ), .B(
        \mult_20/CARRYB[27][2] ), .CI(\mult_20/SUMB[27][3] ), .CO(
        \mult_20/CARRYB[28][2] ), .S(\mult_20/SUMB[28][2] ) );
  FA_X1 \mult_20/S2_28_1  ( .A(\mult_20/ab[28][1] ), .B(
        \mult_20/CARRYB[27][1] ), .CI(\mult_20/SUMB[27][2] ), .CO(
        \mult_20/CARRYB[28][1] ), .S(\mult_20/SUMB[28][1] ) );
  FA_X1 \mult_20/S1_28_0  ( .A(\mult_20/ab[28][0] ), .B(
        \mult_20/CARRYB[27][0] ), .CI(\mult_20/SUMB[27][1] ), .CO(
        \mult_20/CARRYB[28][0] ), .S(N92) );
  FA_X1 \mult_20/S3_29_30  ( .A(\mult_20/ab[29][30] ), .B(
        \mult_20/CARRYB[28][30] ), .CI(\mult_20/ab[28][31] ), .CO(
        \mult_20/CARRYB[29][30] ), .S(\mult_20/SUMB[29][30] ) );
  FA_X1 \mult_20/S2_29_29  ( .A(\mult_20/ab[29][29] ), .B(
        \mult_20/CARRYB[28][29] ), .CI(\mult_20/SUMB[28][30] ), .CO(
        \mult_20/CARRYB[29][29] ), .S(\mult_20/SUMB[29][29] ) );
  FA_X1 \mult_20/S2_29_28  ( .A(\mult_20/ab[29][28] ), .B(
        \mult_20/CARRYB[28][28] ), .CI(\mult_20/SUMB[28][29] ), .CO(
        \mult_20/CARRYB[29][28] ), .S(\mult_20/SUMB[29][28] ) );
  FA_X1 \mult_20/S2_29_27  ( .A(\mult_20/ab[29][27] ), .B(
        \mult_20/CARRYB[28][27] ), .CI(\mult_20/SUMB[28][28] ), .CO(
        \mult_20/CARRYB[29][27] ), .S(\mult_20/SUMB[29][27] ) );
  FA_X1 \mult_20/S2_29_26  ( .A(\mult_20/ab[29][26] ), .B(
        \mult_20/CARRYB[28][26] ), .CI(\mult_20/SUMB[28][27] ), .CO(
        \mult_20/CARRYB[29][26] ), .S(\mult_20/SUMB[29][26] ) );
  FA_X1 \mult_20/S2_29_25  ( .A(\mult_20/ab[29][25] ), .B(
        \mult_20/CARRYB[28][25] ), .CI(\mult_20/SUMB[28][26] ), .CO(
        \mult_20/CARRYB[29][25] ), .S(\mult_20/SUMB[29][25] ) );
  FA_X1 \mult_20/S2_29_24  ( .A(\mult_20/ab[29][24] ), .B(
        \mult_20/CARRYB[28][24] ), .CI(\mult_20/SUMB[28][25] ), .CO(
        \mult_20/CARRYB[29][24] ), .S(\mult_20/SUMB[29][24] ) );
  FA_X1 \mult_20/S2_29_23  ( .A(\mult_20/ab[29][23] ), .B(
        \mult_20/CARRYB[28][23] ), .CI(\mult_20/SUMB[28][24] ), .CO(
        \mult_20/CARRYB[29][23] ), .S(\mult_20/SUMB[29][23] ) );
  FA_X1 \mult_20/S2_29_22  ( .A(\mult_20/ab[29][22] ), .B(
        \mult_20/CARRYB[28][22] ), .CI(\mult_20/SUMB[28][23] ), .CO(
        \mult_20/CARRYB[29][22] ), .S(\mult_20/SUMB[29][22] ) );
  FA_X1 \mult_20/S2_29_21  ( .A(\mult_20/ab[29][21] ), .B(
        \mult_20/CARRYB[28][21] ), .CI(\mult_20/SUMB[28][22] ), .CO(
        \mult_20/CARRYB[29][21] ), .S(\mult_20/SUMB[29][21] ) );
  FA_X1 \mult_20/S2_29_20  ( .A(\mult_20/ab[29][20] ), .B(
        \mult_20/CARRYB[28][20] ), .CI(\mult_20/SUMB[28][21] ), .CO(
        \mult_20/CARRYB[29][20] ), .S(\mult_20/SUMB[29][20] ) );
  FA_X1 \mult_20/S2_29_19  ( .A(\mult_20/ab[29][19] ), .B(
        \mult_20/CARRYB[28][19] ), .CI(\mult_20/SUMB[28][20] ), .CO(
        \mult_20/CARRYB[29][19] ), .S(\mult_20/SUMB[29][19] ) );
  FA_X1 \mult_20/S2_29_18  ( .A(\mult_20/ab[29][18] ), .B(
        \mult_20/CARRYB[28][18] ), .CI(\mult_20/SUMB[28][19] ), .CO(
        \mult_20/CARRYB[29][18] ), .S(\mult_20/SUMB[29][18] ) );
  FA_X1 \mult_20/S2_29_17  ( .A(\mult_20/ab[29][17] ), .B(
        \mult_20/CARRYB[28][17] ), .CI(\mult_20/SUMB[28][18] ), .CO(
        \mult_20/CARRYB[29][17] ), .S(\mult_20/SUMB[29][17] ) );
  FA_X1 \mult_20/S2_29_16  ( .A(\mult_20/ab[29][16] ), .B(
        \mult_20/CARRYB[28][16] ), .CI(\mult_20/SUMB[28][17] ), .CO(
        \mult_20/CARRYB[29][16] ), .S(\mult_20/SUMB[29][16] ) );
  FA_X1 \mult_20/S2_29_15  ( .A(\mult_20/ab[29][15] ), .B(
        \mult_20/CARRYB[28][15] ), .CI(\mult_20/SUMB[28][16] ), .CO(
        \mult_20/CARRYB[29][15] ), .S(\mult_20/SUMB[29][15] ) );
  FA_X1 \mult_20/S2_29_14  ( .A(\mult_20/ab[29][14] ), .B(
        \mult_20/CARRYB[28][14] ), .CI(\mult_20/SUMB[28][15] ), .CO(
        \mult_20/CARRYB[29][14] ), .S(\mult_20/SUMB[29][14] ) );
  FA_X1 \mult_20/S2_29_13  ( .A(\mult_20/ab[29][13] ), .B(
        \mult_20/CARRYB[28][13] ), .CI(\mult_20/SUMB[28][14] ), .CO(
        \mult_20/CARRYB[29][13] ), .S(\mult_20/SUMB[29][13] ) );
  FA_X1 \mult_20/S2_29_12  ( .A(\mult_20/ab[29][12] ), .B(
        \mult_20/CARRYB[28][12] ), .CI(\mult_20/SUMB[28][13] ), .CO(
        \mult_20/CARRYB[29][12] ), .S(\mult_20/SUMB[29][12] ) );
  FA_X1 \mult_20/S2_29_11  ( .A(\mult_20/ab[29][11] ), .B(
        \mult_20/CARRYB[28][11] ), .CI(\mult_20/SUMB[28][12] ), .CO(
        \mult_20/CARRYB[29][11] ), .S(\mult_20/SUMB[29][11] ) );
  FA_X1 \mult_20/S2_29_10  ( .A(\mult_20/ab[29][10] ), .B(
        \mult_20/CARRYB[28][10] ), .CI(\mult_20/SUMB[28][11] ), .CO(
        \mult_20/CARRYB[29][10] ), .S(\mult_20/SUMB[29][10] ) );
  FA_X1 \mult_20/S2_29_9  ( .A(\mult_20/ab[29][9] ), .B(
        \mult_20/CARRYB[28][9] ), .CI(\mult_20/SUMB[28][10] ), .CO(
        \mult_20/CARRYB[29][9] ), .S(\mult_20/SUMB[29][9] ) );
  FA_X1 \mult_20/S2_29_8  ( .A(\mult_20/ab[29][8] ), .B(
        \mult_20/CARRYB[28][8] ), .CI(\mult_20/SUMB[28][9] ), .CO(
        \mult_20/CARRYB[29][8] ), .S(\mult_20/SUMB[29][8] ) );
  FA_X1 \mult_20/S2_29_7  ( .A(\mult_20/ab[29][7] ), .B(
        \mult_20/CARRYB[28][7] ), .CI(\mult_20/SUMB[28][8] ), .CO(
        \mult_20/CARRYB[29][7] ), .S(\mult_20/SUMB[29][7] ) );
  FA_X1 \mult_20/S2_29_6  ( .A(\mult_20/ab[29][6] ), .B(
        \mult_20/CARRYB[28][6] ), .CI(\mult_20/SUMB[28][7] ), .CO(
        \mult_20/CARRYB[29][6] ), .S(\mult_20/SUMB[29][6] ) );
  FA_X1 \mult_20/S2_29_5  ( .A(\mult_20/ab[29][5] ), .B(
        \mult_20/CARRYB[28][5] ), .CI(\mult_20/SUMB[28][6] ), .CO(
        \mult_20/CARRYB[29][5] ), .S(\mult_20/SUMB[29][5] ) );
  FA_X1 \mult_20/S2_29_4  ( .A(\mult_20/ab[29][4] ), .B(
        \mult_20/CARRYB[28][4] ), .CI(\mult_20/SUMB[28][5] ), .CO(
        \mult_20/CARRYB[29][4] ), .S(\mult_20/SUMB[29][4] ) );
  FA_X1 \mult_20/S2_29_3  ( .A(\mult_20/ab[29][3] ), .B(
        \mult_20/CARRYB[28][3] ), .CI(\mult_20/SUMB[28][4] ), .CO(
        \mult_20/CARRYB[29][3] ), .S(\mult_20/SUMB[29][3] ) );
  FA_X1 \mult_20/S2_29_2  ( .A(\mult_20/ab[29][2] ), .B(
        \mult_20/CARRYB[28][2] ), .CI(\mult_20/SUMB[28][3] ), .CO(
        \mult_20/CARRYB[29][2] ), .S(\mult_20/SUMB[29][2] ) );
  FA_X1 \mult_20/S2_29_1  ( .A(\mult_20/ab[29][1] ), .B(
        \mult_20/CARRYB[28][1] ), .CI(\mult_20/SUMB[28][2] ), .CO(
        \mult_20/CARRYB[29][1] ), .S(\mult_20/SUMB[29][1] ) );
  FA_X1 \mult_20/S1_29_0  ( .A(\mult_20/ab[29][0] ), .B(
        \mult_20/CARRYB[28][0] ), .CI(\mult_20/SUMB[28][1] ), .CO(
        \mult_20/CARRYB[29][0] ), .S(N93) );
  FA_X1 \mult_20/S3_30_30  ( .A(\mult_20/ab[30][30] ), .B(
        \mult_20/CARRYB[29][30] ), .CI(\mult_20/ab[29][31] ), .CO(
        \mult_20/CARRYB[30][30] ), .S(\mult_20/SUMB[30][30] ) );
  FA_X1 \mult_20/S2_30_29  ( .A(\mult_20/ab[30][29] ), .B(
        \mult_20/CARRYB[29][29] ), .CI(\mult_20/SUMB[29][30] ), .CO(
        \mult_20/CARRYB[30][29] ), .S(\mult_20/SUMB[30][29] ) );
  FA_X1 \mult_20/S2_30_28  ( .A(\mult_20/ab[30][28] ), .B(
        \mult_20/CARRYB[29][28] ), .CI(\mult_20/SUMB[29][29] ), .CO(
        \mult_20/CARRYB[30][28] ), .S(\mult_20/SUMB[30][28] ) );
  FA_X1 \mult_20/S2_30_27  ( .A(\mult_20/ab[30][27] ), .B(
        \mult_20/CARRYB[29][27] ), .CI(\mult_20/SUMB[29][28] ), .CO(
        \mult_20/CARRYB[30][27] ), .S(\mult_20/SUMB[30][27] ) );
  FA_X1 \mult_20/S2_30_26  ( .A(\mult_20/ab[30][26] ), .B(
        \mult_20/CARRYB[29][26] ), .CI(\mult_20/SUMB[29][27] ), .CO(
        \mult_20/CARRYB[30][26] ), .S(\mult_20/SUMB[30][26] ) );
  FA_X1 \mult_20/S2_30_25  ( .A(\mult_20/ab[30][25] ), .B(
        \mult_20/CARRYB[29][25] ), .CI(\mult_20/SUMB[29][26] ), .CO(
        \mult_20/CARRYB[30][25] ), .S(\mult_20/SUMB[30][25] ) );
  FA_X1 \mult_20/S2_30_24  ( .A(\mult_20/ab[30][24] ), .B(
        \mult_20/CARRYB[29][24] ), .CI(\mult_20/SUMB[29][25] ), .CO(
        \mult_20/CARRYB[30][24] ), .S(\mult_20/SUMB[30][24] ) );
  FA_X1 \mult_20/S2_30_23  ( .A(\mult_20/ab[30][23] ), .B(
        \mult_20/CARRYB[29][23] ), .CI(\mult_20/SUMB[29][24] ), .CO(
        \mult_20/CARRYB[30][23] ), .S(\mult_20/SUMB[30][23] ) );
  FA_X1 \mult_20/S2_30_22  ( .A(\mult_20/ab[30][22] ), .B(
        \mult_20/CARRYB[29][22] ), .CI(\mult_20/SUMB[29][23] ), .CO(
        \mult_20/CARRYB[30][22] ), .S(\mult_20/SUMB[30][22] ) );
  FA_X1 \mult_20/S2_30_21  ( .A(\mult_20/ab[30][21] ), .B(
        \mult_20/CARRYB[29][21] ), .CI(\mult_20/SUMB[29][22] ), .CO(
        \mult_20/CARRYB[30][21] ), .S(\mult_20/SUMB[30][21] ) );
  FA_X1 \mult_20/S2_30_20  ( .A(\mult_20/ab[30][20] ), .B(
        \mult_20/CARRYB[29][20] ), .CI(\mult_20/SUMB[29][21] ), .CO(
        \mult_20/CARRYB[30][20] ), .S(\mult_20/SUMB[30][20] ) );
  FA_X1 \mult_20/S2_30_19  ( .A(\mult_20/ab[30][19] ), .B(
        \mult_20/CARRYB[29][19] ), .CI(\mult_20/SUMB[29][20] ), .CO(
        \mult_20/CARRYB[30][19] ), .S(\mult_20/SUMB[30][19] ) );
  FA_X1 \mult_20/S2_30_18  ( .A(\mult_20/ab[30][18] ), .B(
        \mult_20/CARRYB[29][18] ), .CI(\mult_20/SUMB[29][19] ), .CO(
        \mult_20/CARRYB[30][18] ), .S(\mult_20/SUMB[30][18] ) );
  FA_X1 \mult_20/S2_30_17  ( .A(\mult_20/ab[30][17] ), .B(
        \mult_20/CARRYB[29][17] ), .CI(\mult_20/SUMB[29][18] ), .CO(
        \mult_20/CARRYB[30][17] ), .S(\mult_20/SUMB[30][17] ) );
  FA_X1 \mult_20/S2_30_16  ( .A(\mult_20/ab[30][16] ), .B(
        \mult_20/CARRYB[29][16] ), .CI(\mult_20/SUMB[29][17] ), .CO(
        \mult_20/CARRYB[30][16] ), .S(\mult_20/SUMB[30][16] ) );
  FA_X1 \mult_20/S2_30_15  ( .A(\mult_20/ab[30][15] ), .B(
        \mult_20/CARRYB[29][15] ), .CI(\mult_20/SUMB[29][16] ), .CO(
        \mult_20/CARRYB[30][15] ), .S(\mult_20/SUMB[30][15] ) );
  FA_X1 \mult_20/S2_30_14  ( .A(\mult_20/ab[30][14] ), .B(
        \mult_20/CARRYB[29][14] ), .CI(\mult_20/SUMB[29][15] ), .CO(
        \mult_20/CARRYB[30][14] ), .S(\mult_20/SUMB[30][14] ) );
  FA_X1 \mult_20/S2_30_13  ( .A(\mult_20/ab[30][13] ), .B(
        \mult_20/CARRYB[29][13] ), .CI(\mult_20/SUMB[29][14] ), .CO(
        \mult_20/CARRYB[30][13] ), .S(\mult_20/SUMB[30][13] ) );
  FA_X1 \mult_20/S2_30_12  ( .A(\mult_20/ab[30][12] ), .B(
        \mult_20/CARRYB[29][12] ), .CI(\mult_20/SUMB[29][13] ), .CO(
        \mult_20/CARRYB[30][12] ), .S(\mult_20/SUMB[30][12] ) );
  FA_X1 \mult_20/S2_30_11  ( .A(\mult_20/ab[30][11] ), .B(
        \mult_20/CARRYB[29][11] ), .CI(\mult_20/SUMB[29][12] ), .CO(
        \mult_20/CARRYB[30][11] ), .S(\mult_20/SUMB[30][11] ) );
  FA_X1 \mult_20/S2_30_10  ( .A(\mult_20/ab[30][10] ), .B(
        \mult_20/CARRYB[29][10] ), .CI(\mult_20/SUMB[29][11] ), .CO(
        \mult_20/CARRYB[30][10] ), .S(\mult_20/SUMB[30][10] ) );
  FA_X1 \mult_20/S2_30_9  ( .A(\mult_20/ab[30][9] ), .B(
        \mult_20/CARRYB[29][9] ), .CI(\mult_20/SUMB[29][10] ), .CO(
        \mult_20/CARRYB[30][9] ), .S(\mult_20/SUMB[30][9] ) );
  FA_X1 \mult_20/S2_30_8  ( .A(\mult_20/ab[30][8] ), .B(
        \mult_20/CARRYB[29][8] ), .CI(\mult_20/SUMB[29][9] ), .CO(
        \mult_20/CARRYB[30][8] ), .S(\mult_20/SUMB[30][8] ) );
  FA_X1 \mult_20/S2_30_7  ( .A(\mult_20/ab[30][7] ), .B(
        \mult_20/CARRYB[29][7] ), .CI(\mult_20/SUMB[29][8] ), .CO(
        \mult_20/CARRYB[30][7] ), .S(\mult_20/SUMB[30][7] ) );
  FA_X1 \mult_20/S2_30_6  ( .A(\mult_20/ab[30][6] ), .B(
        \mult_20/CARRYB[29][6] ), .CI(\mult_20/SUMB[29][7] ), .CO(
        \mult_20/CARRYB[30][6] ), .S(\mult_20/SUMB[30][6] ) );
  FA_X1 \mult_20/S2_30_5  ( .A(\mult_20/ab[30][5] ), .B(
        \mult_20/CARRYB[29][5] ), .CI(\mult_20/SUMB[29][6] ), .CO(
        \mult_20/CARRYB[30][5] ), .S(\mult_20/SUMB[30][5] ) );
  FA_X1 \mult_20/S2_30_4  ( .A(\mult_20/ab[30][4] ), .B(
        \mult_20/CARRYB[29][4] ), .CI(\mult_20/SUMB[29][5] ), .CO(
        \mult_20/CARRYB[30][4] ), .S(\mult_20/SUMB[30][4] ) );
  FA_X1 \mult_20/S2_30_3  ( .A(\mult_20/ab[30][3] ), .B(
        \mult_20/CARRYB[29][3] ), .CI(\mult_20/SUMB[29][4] ), .CO(
        \mult_20/CARRYB[30][3] ), .S(\mult_20/SUMB[30][3] ) );
  FA_X1 \mult_20/S2_30_2  ( .A(\mult_20/ab[30][2] ), .B(
        \mult_20/CARRYB[29][2] ), .CI(\mult_20/SUMB[29][3] ), .CO(
        \mult_20/CARRYB[30][2] ), .S(\mult_20/SUMB[30][2] ) );
  FA_X1 \mult_20/S2_30_1  ( .A(\mult_20/ab[30][1] ), .B(
        \mult_20/CARRYB[29][1] ), .CI(\mult_20/SUMB[29][2] ), .CO(
        \mult_20/CARRYB[30][1] ), .S(\mult_20/SUMB[30][1] ) );
  FA_X1 \mult_20/S1_30_0  ( .A(\mult_20/ab[30][0] ), .B(
        \mult_20/CARRYB[29][0] ), .CI(\mult_20/SUMB[29][1] ), .CO(
        \mult_20/CARRYB[30][0] ), .S(N94) );
  FA_X1 \mult_20/S5_30  ( .A(\mult_20/ab[31][30] ), .B(
        \mult_20/CARRYB[30][30] ), .CI(\mult_20/ab[30][31] ), .CO(
        \mult_20/CARRYB[31][30] ), .S(\mult_20/SUMB[31][30] ) );
  FA_X1 \mult_20/S4_29  ( .A(\mult_20/ab[31][29] ), .B(
        \mult_20/CARRYB[30][29] ), .CI(\mult_20/SUMB[30][30] ), .CO(
        \mult_20/CARRYB[31][29] ), .S(\mult_20/SUMB[31][29] ) );
  FA_X1 \mult_20/S4_28  ( .A(\mult_20/ab[31][28] ), .B(
        \mult_20/CARRYB[30][28] ), .CI(\mult_20/SUMB[30][29] ), .CO(
        \mult_20/CARRYB[31][28] ), .S(\mult_20/SUMB[31][28] ) );
  FA_X1 \mult_20/S4_27  ( .A(\mult_20/ab[31][27] ), .B(
        \mult_20/CARRYB[30][27] ), .CI(\mult_20/SUMB[30][28] ), .CO(
        \mult_20/CARRYB[31][27] ), .S(\mult_20/SUMB[31][27] ) );
  FA_X1 \mult_20/S4_26  ( .A(\mult_20/ab[31][26] ), .B(
        \mult_20/CARRYB[30][26] ), .CI(\mult_20/SUMB[30][27] ), .CO(
        \mult_20/CARRYB[31][26] ), .S(\mult_20/SUMB[31][26] ) );
  FA_X1 \mult_20/S4_25  ( .A(\mult_20/ab[31][25] ), .B(
        \mult_20/CARRYB[30][25] ), .CI(\mult_20/SUMB[30][26] ), .CO(
        \mult_20/CARRYB[31][25] ), .S(\mult_20/SUMB[31][25] ) );
  FA_X1 \mult_20/S4_24  ( .A(\mult_20/ab[31][24] ), .B(
        \mult_20/CARRYB[30][24] ), .CI(\mult_20/SUMB[30][25] ), .CO(
        \mult_20/CARRYB[31][24] ), .S(\mult_20/SUMB[31][24] ) );
  FA_X1 \mult_20/S4_23  ( .A(\mult_20/ab[31][23] ), .B(
        \mult_20/CARRYB[30][23] ), .CI(\mult_20/SUMB[30][24] ), .CO(
        \mult_20/CARRYB[31][23] ), .S(\mult_20/SUMB[31][23] ) );
  FA_X1 \mult_20/S4_22  ( .A(\mult_20/ab[31][22] ), .B(
        \mult_20/CARRYB[30][22] ), .CI(\mult_20/SUMB[30][23] ), .CO(
        \mult_20/CARRYB[31][22] ), .S(\mult_20/SUMB[31][22] ) );
  FA_X1 \mult_20/S4_21  ( .A(\mult_20/ab[31][21] ), .B(
        \mult_20/CARRYB[30][21] ), .CI(\mult_20/SUMB[30][22] ), .CO(
        \mult_20/CARRYB[31][21] ), .S(\mult_20/SUMB[31][21] ) );
  FA_X1 \mult_20/S4_20  ( .A(\mult_20/ab[31][20] ), .B(
        \mult_20/CARRYB[30][20] ), .CI(\mult_20/SUMB[30][21] ), .CO(
        \mult_20/CARRYB[31][20] ), .S(\mult_20/SUMB[31][20] ) );
  FA_X1 \mult_20/S4_19  ( .A(\mult_20/ab[31][19] ), .B(
        \mult_20/CARRYB[30][19] ), .CI(\mult_20/SUMB[30][20] ), .CO(
        \mult_20/CARRYB[31][19] ), .S(\mult_20/SUMB[31][19] ) );
  FA_X1 \mult_20/S4_18  ( .A(\mult_20/ab[31][18] ), .B(
        \mult_20/CARRYB[30][18] ), .CI(\mult_20/SUMB[30][19] ), .CO(
        \mult_20/CARRYB[31][18] ), .S(\mult_20/SUMB[31][18] ) );
  FA_X1 \mult_20/S4_17  ( .A(\mult_20/ab[31][17] ), .B(
        \mult_20/CARRYB[30][17] ), .CI(\mult_20/SUMB[30][18] ), .CO(
        \mult_20/CARRYB[31][17] ), .S(\mult_20/SUMB[31][17] ) );
  FA_X1 \mult_20/S4_16  ( .A(\mult_20/ab[31][16] ), .B(
        \mult_20/CARRYB[30][16] ), .CI(\mult_20/SUMB[30][17] ), .CO(
        \mult_20/CARRYB[31][16] ), .S(\mult_20/SUMB[31][16] ) );
  FA_X1 \mult_20/S4_15  ( .A(\mult_20/ab[31][15] ), .B(
        \mult_20/CARRYB[30][15] ), .CI(\mult_20/SUMB[30][16] ), .CO(
        \mult_20/CARRYB[31][15] ), .S(\mult_20/SUMB[31][15] ) );
  FA_X1 \mult_20/S4_14  ( .A(\mult_20/ab[31][14] ), .B(
        \mult_20/CARRYB[30][14] ), .CI(\mult_20/SUMB[30][15] ), .CO(
        \mult_20/CARRYB[31][14] ), .S(\mult_20/SUMB[31][14] ) );
  FA_X1 \mult_20/S4_13  ( .A(\mult_20/ab[31][13] ), .B(
        \mult_20/CARRYB[30][13] ), .CI(\mult_20/SUMB[30][14] ), .CO(
        \mult_20/CARRYB[31][13] ), .S(\mult_20/SUMB[31][13] ) );
  FA_X1 \mult_20/S4_12  ( .A(\mult_20/ab[31][12] ), .B(
        \mult_20/CARRYB[30][12] ), .CI(\mult_20/SUMB[30][13] ), .CO(
        \mult_20/CARRYB[31][12] ), .S(\mult_20/SUMB[31][12] ) );
  FA_X1 \mult_20/S4_11  ( .A(\mult_20/ab[31][11] ), .B(
        \mult_20/CARRYB[30][11] ), .CI(\mult_20/SUMB[30][12] ), .CO(
        \mult_20/CARRYB[31][11] ), .S(\mult_20/SUMB[31][11] ) );
  FA_X1 \mult_20/S4_10  ( .A(\mult_20/ab[31][10] ), .B(
        \mult_20/CARRYB[30][10] ), .CI(\mult_20/SUMB[30][11] ), .CO(
        \mult_20/CARRYB[31][10] ), .S(\mult_20/SUMB[31][10] ) );
  FA_X1 \mult_20/S4_9  ( .A(\mult_20/ab[31][9] ), .B(\mult_20/CARRYB[30][9] ), 
        .CI(\mult_20/SUMB[30][10] ), .CO(\mult_20/CARRYB[31][9] ), .S(
        \mult_20/SUMB[31][9] ) );
  FA_X1 \mult_20/S4_8  ( .A(\mult_20/ab[31][8] ), .B(\mult_20/CARRYB[30][8] ), 
        .CI(\mult_20/SUMB[30][9] ), .CO(\mult_20/CARRYB[31][8] ), .S(
        \mult_20/SUMB[31][8] ) );
  FA_X1 \mult_20/S4_7  ( .A(\mult_20/ab[31][7] ), .B(\mult_20/CARRYB[30][7] ), 
        .CI(\mult_20/SUMB[30][8] ), .CO(\mult_20/CARRYB[31][7] ), .S(
        \mult_20/SUMB[31][7] ) );
  FA_X1 \mult_20/S4_6  ( .A(\mult_20/ab[31][6] ), .B(\mult_20/CARRYB[30][6] ), 
        .CI(\mult_20/SUMB[30][7] ), .CO(\mult_20/CARRYB[31][6] ), .S(
        \mult_20/SUMB[31][6] ) );
  FA_X1 \mult_20/S4_5  ( .A(\mult_20/ab[31][5] ), .B(\mult_20/CARRYB[30][5] ), 
        .CI(\mult_20/SUMB[30][6] ), .CO(\mult_20/CARRYB[31][5] ), .S(
        \mult_20/SUMB[31][5] ) );
  FA_X1 \mult_20/S4_4  ( .A(\mult_20/ab[31][4] ), .B(\mult_20/CARRYB[30][4] ), 
        .CI(\mult_20/SUMB[30][5] ), .CO(\mult_20/CARRYB[31][4] ), .S(
        \mult_20/SUMB[31][4] ) );
  FA_X1 \mult_20/S4_3  ( .A(\mult_20/ab[31][3] ), .B(\mult_20/CARRYB[30][3] ), 
        .CI(\mult_20/SUMB[30][4] ), .CO(\mult_20/CARRYB[31][3] ), .S(
        \mult_20/SUMB[31][3] ) );
  FA_X1 \mult_20/S4_2  ( .A(\mult_20/ab[31][2] ), .B(\mult_20/CARRYB[30][2] ), 
        .CI(\mult_20/SUMB[30][3] ), .CO(\mult_20/CARRYB[31][2] ), .S(
        \mult_20/SUMB[31][2] ) );
  FA_X1 \mult_20/S4_1  ( .A(\mult_20/ab[31][1] ), .B(\mult_20/CARRYB[30][1] ), 
        .CI(\mult_20/SUMB[30][2] ), .CO(\mult_20/CARRYB[31][1] ), .S(
        \mult_20/SUMB[31][1] ) );
  FA_X1 \mult_20/S4_0  ( .A(\mult_20/ab[31][0] ), .B(\mult_20/CARRYB[30][0] ), 
        .CI(\mult_20/SUMB[30][1] ), .CO(\mult_20/CARRYB[31][0] ), .S(N95) );
  FA_X1 \mult_19/S3_2_30  ( .A(\mult_19/ab[2][30] ), .B(\mult_19/n33 ), .CI(
        \mult_19/ab[1][31] ), .CO(\mult_19/CARRYB[2][30] ), .S(
        \mult_19/SUMB[2][30] ) );
  FA_X1 \mult_19/S2_2_29  ( .A(\mult_19/ab[2][29] ), .B(\mult_19/n3 ), .CI(
        \mult_19/n34 ), .CO(\mult_19/CARRYB[2][29] ), .S(\mult_19/SUMB[2][29] ) );
  FA_X1 \mult_19/S2_2_28  ( .A(\mult_19/ab[2][28] ), .B(\mult_19/n4 ), .CI(
        \mult_19/n35 ), .CO(\mult_19/CARRYB[2][28] ), .S(\mult_19/SUMB[2][28] ) );
  FA_X1 \mult_19/S2_2_27  ( .A(\mult_19/ab[2][27] ), .B(\mult_19/n5 ), .CI(
        \mult_19/n36 ), .CO(\mult_19/CARRYB[2][27] ), .S(\mult_19/SUMB[2][27] ) );
  FA_X1 \mult_19/S2_2_26  ( .A(\mult_19/ab[2][26] ), .B(\mult_19/n6 ), .CI(
        \mult_19/n37 ), .CO(\mult_19/CARRYB[2][26] ), .S(\mult_19/SUMB[2][26] ) );
  FA_X1 \mult_19/S2_2_25  ( .A(\mult_19/ab[2][25] ), .B(\mult_19/n7 ), .CI(
        \mult_19/n38 ), .CO(\mult_19/CARRYB[2][25] ), .S(\mult_19/SUMB[2][25] ) );
  FA_X1 \mult_19/S2_2_24  ( .A(\mult_19/ab[2][24] ), .B(\mult_19/n8 ), .CI(
        \mult_19/n39 ), .CO(\mult_19/CARRYB[2][24] ), .S(\mult_19/SUMB[2][24] ) );
  FA_X1 \mult_19/S2_2_23  ( .A(\mult_19/ab[2][23] ), .B(\mult_19/n9 ), .CI(
        \mult_19/n40 ), .CO(\mult_19/CARRYB[2][23] ), .S(\mult_19/SUMB[2][23] ) );
  FA_X1 \mult_19/S2_2_22  ( .A(\mult_19/ab[2][22] ), .B(\mult_19/n10 ), .CI(
        \mult_19/n41 ), .CO(\mult_19/CARRYB[2][22] ), .S(\mult_19/SUMB[2][22] ) );
  FA_X1 \mult_19/S2_2_21  ( .A(\mult_19/ab[2][21] ), .B(\mult_19/n11 ), .CI(
        \mult_19/n42 ), .CO(\mult_19/CARRYB[2][21] ), .S(\mult_19/SUMB[2][21] ) );
  FA_X1 \mult_19/S2_2_20  ( .A(\mult_19/ab[2][20] ), .B(\mult_19/n12 ), .CI(
        \mult_19/n43 ), .CO(\mult_19/CARRYB[2][20] ), .S(\mult_19/SUMB[2][20] ) );
  FA_X1 \mult_19/S2_2_19  ( .A(\mult_19/ab[2][19] ), .B(\mult_19/n13 ), .CI(
        \mult_19/n44 ), .CO(\mult_19/CARRYB[2][19] ), .S(\mult_19/SUMB[2][19] ) );
  FA_X1 \mult_19/S2_2_18  ( .A(\mult_19/ab[2][18] ), .B(\mult_19/n14 ), .CI(
        \mult_19/n45 ), .CO(\mult_19/CARRYB[2][18] ), .S(\mult_19/SUMB[2][18] ) );
  FA_X1 \mult_19/S2_2_17  ( .A(\mult_19/ab[2][17] ), .B(\mult_19/n15 ), .CI(
        \mult_19/n46 ), .CO(\mult_19/CARRYB[2][17] ), .S(\mult_19/SUMB[2][17] ) );
  FA_X1 \mult_19/S2_2_16  ( .A(\mult_19/ab[2][16] ), .B(\mult_19/n16 ), .CI(
        \mult_19/n47 ), .CO(\mult_19/CARRYB[2][16] ), .S(\mult_19/SUMB[2][16] ) );
  FA_X1 \mult_19/S2_2_15  ( .A(\mult_19/ab[2][15] ), .B(\mult_19/n17 ), .CI(
        \mult_19/n48 ), .CO(\mult_19/CARRYB[2][15] ), .S(\mult_19/SUMB[2][15] ) );
  FA_X1 \mult_19/S2_2_14  ( .A(\mult_19/ab[2][14] ), .B(\mult_19/n18 ), .CI(
        \mult_19/n49 ), .CO(\mult_19/CARRYB[2][14] ), .S(\mult_19/SUMB[2][14] ) );
  FA_X1 \mult_19/S2_2_13  ( .A(\mult_19/ab[2][13] ), .B(\mult_19/n19 ), .CI(
        \mult_19/n50 ), .CO(\mult_19/CARRYB[2][13] ), .S(\mult_19/SUMB[2][13] ) );
  FA_X1 \mult_19/S2_2_12  ( .A(\mult_19/ab[2][12] ), .B(\mult_19/n20 ), .CI(
        \mult_19/n51 ), .CO(\mult_19/CARRYB[2][12] ), .S(\mult_19/SUMB[2][12] ) );
  FA_X1 \mult_19/S2_2_11  ( .A(\mult_19/ab[2][11] ), .B(\mult_19/n21 ), .CI(
        \mult_19/n52 ), .CO(\mult_19/CARRYB[2][11] ), .S(\mult_19/SUMB[2][11] ) );
  FA_X1 \mult_19/S2_2_10  ( .A(\mult_19/ab[2][10] ), .B(\mult_19/n22 ), .CI(
        \mult_19/n53 ), .CO(\mult_19/CARRYB[2][10] ), .S(\mult_19/SUMB[2][10] ) );
  FA_X1 \mult_19/S2_2_9  ( .A(\mult_19/ab[2][9] ), .B(\mult_19/n23 ), .CI(
        \mult_19/n54 ), .CO(\mult_19/CARRYB[2][9] ), .S(\mult_19/SUMB[2][9] )
         );
  FA_X1 \mult_19/S2_2_8  ( .A(\mult_19/ab[2][8] ), .B(\mult_19/n24 ), .CI(
        \mult_19/n55 ), .CO(\mult_19/CARRYB[2][8] ), .S(\mult_19/SUMB[2][8] )
         );
  FA_X1 \mult_19/S2_2_7  ( .A(\mult_19/ab[2][7] ), .B(\mult_19/n25 ), .CI(
        \mult_19/n56 ), .CO(\mult_19/CARRYB[2][7] ), .S(\mult_19/SUMB[2][7] )
         );
  FA_X1 \mult_19/S2_2_6  ( .A(\mult_19/ab[2][6] ), .B(\mult_19/n26 ), .CI(
        \mult_19/n57 ), .CO(\mult_19/CARRYB[2][6] ), .S(\mult_19/SUMB[2][6] )
         );
  FA_X1 \mult_19/S2_2_5  ( .A(\mult_19/ab[2][5] ), .B(\mult_19/n27 ), .CI(
        \mult_19/n58 ), .CO(\mult_19/CARRYB[2][5] ), .S(\mult_19/SUMB[2][5] )
         );
  FA_X1 \mult_19/S2_2_4  ( .A(\mult_19/ab[2][4] ), .B(\mult_19/n28 ), .CI(
        \mult_19/n59 ), .CO(\mult_19/CARRYB[2][4] ), .S(\mult_19/SUMB[2][4] )
         );
  FA_X1 \mult_19/S2_2_3  ( .A(\mult_19/ab[2][3] ), .B(\mult_19/n29 ), .CI(
        \mult_19/n60 ), .CO(\mult_19/CARRYB[2][3] ), .S(\mult_19/SUMB[2][3] )
         );
  FA_X1 \mult_19/S2_2_2  ( .A(\mult_19/ab[2][2] ), .B(\mult_19/n30 ), .CI(
        \mult_19/n61 ), .CO(\mult_19/CARRYB[2][2] ), .S(\mult_19/SUMB[2][2] )
         );
  FA_X1 \mult_19/S2_2_1  ( .A(\mult_19/ab[2][1] ), .B(\mult_19/n31 ), .CI(
        \mult_19/n62 ), .CO(\mult_19/CARRYB[2][1] ), .S(\mult_19/SUMB[2][1] )
         );
  FA_X1 \mult_19/S1_2_0  ( .A(\mult_19/ab[2][0] ), .B(\mult_19/n32 ), .CI(
        \mult_19/n63 ), .CO(\mult_19/CARRYB[2][0] ), .S(N2) );
  FA_X1 \mult_19/S3_3_30  ( .A(\mult_19/ab[3][30] ), .B(
        \mult_19/CARRYB[2][30] ), .CI(\mult_19/ab[2][31] ), .CO(
        \mult_19/CARRYB[3][30] ), .S(\mult_19/SUMB[3][30] ) );
  FA_X1 \mult_19/S2_3_29  ( .A(\mult_19/ab[3][29] ), .B(
        \mult_19/CARRYB[2][29] ), .CI(\mult_19/SUMB[2][30] ), .CO(
        \mult_19/CARRYB[3][29] ), .S(\mult_19/SUMB[3][29] ) );
  FA_X1 \mult_19/S2_3_28  ( .A(\mult_19/ab[3][28] ), .B(
        \mult_19/CARRYB[2][28] ), .CI(\mult_19/SUMB[2][29] ), .CO(
        \mult_19/CARRYB[3][28] ), .S(\mult_19/SUMB[3][28] ) );
  FA_X1 \mult_19/S2_3_27  ( .A(\mult_19/ab[3][27] ), .B(
        \mult_19/CARRYB[2][27] ), .CI(\mult_19/SUMB[2][28] ), .CO(
        \mult_19/CARRYB[3][27] ), .S(\mult_19/SUMB[3][27] ) );
  FA_X1 \mult_19/S2_3_26  ( .A(\mult_19/ab[3][26] ), .B(
        \mult_19/CARRYB[2][26] ), .CI(\mult_19/SUMB[2][27] ), .CO(
        \mult_19/CARRYB[3][26] ), .S(\mult_19/SUMB[3][26] ) );
  FA_X1 \mult_19/S2_3_25  ( .A(\mult_19/ab[3][25] ), .B(
        \mult_19/CARRYB[2][25] ), .CI(\mult_19/SUMB[2][26] ), .CO(
        \mult_19/CARRYB[3][25] ), .S(\mult_19/SUMB[3][25] ) );
  FA_X1 \mult_19/S2_3_24  ( .A(\mult_19/ab[3][24] ), .B(
        \mult_19/CARRYB[2][24] ), .CI(\mult_19/SUMB[2][25] ), .CO(
        \mult_19/CARRYB[3][24] ), .S(\mult_19/SUMB[3][24] ) );
  FA_X1 \mult_19/S2_3_23  ( .A(\mult_19/ab[3][23] ), .B(
        \mult_19/CARRYB[2][23] ), .CI(\mult_19/SUMB[2][24] ), .CO(
        \mult_19/CARRYB[3][23] ), .S(\mult_19/SUMB[3][23] ) );
  FA_X1 \mult_19/S2_3_22  ( .A(\mult_19/ab[3][22] ), .B(
        \mult_19/CARRYB[2][22] ), .CI(\mult_19/SUMB[2][23] ), .CO(
        \mult_19/CARRYB[3][22] ), .S(\mult_19/SUMB[3][22] ) );
  FA_X1 \mult_19/S2_3_21  ( .A(\mult_19/ab[3][21] ), .B(
        \mult_19/CARRYB[2][21] ), .CI(\mult_19/SUMB[2][22] ), .CO(
        \mult_19/CARRYB[3][21] ), .S(\mult_19/SUMB[3][21] ) );
  FA_X1 \mult_19/S2_3_20  ( .A(\mult_19/ab[3][20] ), .B(
        \mult_19/CARRYB[2][20] ), .CI(\mult_19/SUMB[2][21] ), .CO(
        \mult_19/CARRYB[3][20] ), .S(\mult_19/SUMB[3][20] ) );
  FA_X1 \mult_19/S2_3_19  ( .A(\mult_19/ab[3][19] ), .B(
        \mult_19/CARRYB[2][19] ), .CI(\mult_19/SUMB[2][20] ), .CO(
        \mult_19/CARRYB[3][19] ), .S(\mult_19/SUMB[3][19] ) );
  FA_X1 \mult_19/S2_3_18  ( .A(\mult_19/ab[3][18] ), .B(
        \mult_19/CARRYB[2][18] ), .CI(\mult_19/SUMB[2][19] ), .CO(
        \mult_19/CARRYB[3][18] ), .S(\mult_19/SUMB[3][18] ) );
  FA_X1 \mult_19/S2_3_17  ( .A(\mult_19/ab[3][17] ), .B(
        \mult_19/CARRYB[2][17] ), .CI(\mult_19/SUMB[2][18] ), .CO(
        \mult_19/CARRYB[3][17] ), .S(\mult_19/SUMB[3][17] ) );
  FA_X1 \mult_19/S2_3_16  ( .A(\mult_19/ab[3][16] ), .B(
        \mult_19/CARRYB[2][16] ), .CI(\mult_19/SUMB[2][17] ), .CO(
        \mult_19/CARRYB[3][16] ), .S(\mult_19/SUMB[3][16] ) );
  FA_X1 \mult_19/S2_3_15  ( .A(\mult_19/ab[3][15] ), .B(
        \mult_19/CARRYB[2][15] ), .CI(\mult_19/SUMB[2][16] ), .CO(
        \mult_19/CARRYB[3][15] ), .S(\mult_19/SUMB[3][15] ) );
  FA_X1 \mult_19/S2_3_14  ( .A(\mult_19/ab[3][14] ), .B(
        \mult_19/CARRYB[2][14] ), .CI(\mult_19/SUMB[2][15] ), .CO(
        \mult_19/CARRYB[3][14] ), .S(\mult_19/SUMB[3][14] ) );
  FA_X1 \mult_19/S2_3_13  ( .A(\mult_19/ab[3][13] ), .B(
        \mult_19/CARRYB[2][13] ), .CI(\mult_19/SUMB[2][14] ), .CO(
        \mult_19/CARRYB[3][13] ), .S(\mult_19/SUMB[3][13] ) );
  FA_X1 \mult_19/S2_3_12  ( .A(\mult_19/ab[3][12] ), .B(
        \mult_19/CARRYB[2][12] ), .CI(\mult_19/SUMB[2][13] ), .CO(
        \mult_19/CARRYB[3][12] ), .S(\mult_19/SUMB[3][12] ) );
  FA_X1 \mult_19/S2_3_11  ( .A(\mult_19/ab[3][11] ), .B(
        \mult_19/CARRYB[2][11] ), .CI(\mult_19/SUMB[2][12] ), .CO(
        \mult_19/CARRYB[3][11] ), .S(\mult_19/SUMB[3][11] ) );
  FA_X1 \mult_19/S2_3_10  ( .A(\mult_19/ab[3][10] ), .B(
        \mult_19/CARRYB[2][10] ), .CI(\mult_19/SUMB[2][11] ), .CO(
        \mult_19/CARRYB[3][10] ), .S(\mult_19/SUMB[3][10] ) );
  FA_X1 \mult_19/S2_3_9  ( .A(\mult_19/ab[3][9] ), .B(\mult_19/CARRYB[2][9] ), 
        .CI(\mult_19/SUMB[2][10] ), .CO(\mult_19/CARRYB[3][9] ), .S(
        \mult_19/SUMB[3][9] ) );
  FA_X1 \mult_19/S2_3_8  ( .A(\mult_19/ab[3][8] ), .B(\mult_19/CARRYB[2][8] ), 
        .CI(\mult_19/SUMB[2][9] ), .CO(\mult_19/CARRYB[3][8] ), .S(
        \mult_19/SUMB[3][8] ) );
  FA_X1 \mult_19/S2_3_7  ( .A(\mult_19/ab[3][7] ), .B(\mult_19/CARRYB[2][7] ), 
        .CI(\mult_19/SUMB[2][8] ), .CO(\mult_19/CARRYB[3][7] ), .S(
        \mult_19/SUMB[3][7] ) );
  FA_X1 \mult_19/S2_3_6  ( .A(\mult_19/ab[3][6] ), .B(\mult_19/CARRYB[2][6] ), 
        .CI(\mult_19/SUMB[2][7] ), .CO(\mult_19/CARRYB[3][6] ), .S(
        \mult_19/SUMB[3][6] ) );
  FA_X1 \mult_19/S2_3_5  ( .A(\mult_19/ab[3][5] ), .B(\mult_19/CARRYB[2][5] ), 
        .CI(\mult_19/SUMB[2][6] ), .CO(\mult_19/CARRYB[3][5] ), .S(
        \mult_19/SUMB[3][5] ) );
  FA_X1 \mult_19/S2_3_4  ( .A(\mult_19/ab[3][4] ), .B(\mult_19/CARRYB[2][4] ), 
        .CI(\mult_19/SUMB[2][5] ), .CO(\mult_19/CARRYB[3][4] ), .S(
        \mult_19/SUMB[3][4] ) );
  FA_X1 \mult_19/S2_3_3  ( .A(\mult_19/ab[3][3] ), .B(\mult_19/CARRYB[2][3] ), 
        .CI(\mult_19/SUMB[2][4] ), .CO(\mult_19/CARRYB[3][3] ), .S(
        \mult_19/SUMB[3][3] ) );
  FA_X1 \mult_19/S2_3_2  ( .A(\mult_19/ab[3][2] ), .B(\mult_19/CARRYB[2][2] ), 
        .CI(\mult_19/SUMB[2][3] ), .CO(\mult_19/CARRYB[3][2] ), .S(
        \mult_19/SUMB[3][2] ) );
  FA_X1 \mult_19/S2_3_1  ( .A(\mult_19/ab[3][1] ), .B(\mult_19/CARRYB[2][1] ), 
        .CI(\mult_19/SUMB[2][2] ), .CO(\mult_19/CARRYB[3][1] ), .S(
        \mult_19/SUMB[3][1] ) );
  FA_X1 \mult_19/S1_3_0  ( .A(\mult_19/ab[3][0] ), .B(\mult_19/CARRYB[2][0] ), 
        .CI(\mult_19/SUMB[2][1] ), .CO(\mult_19/CARRYB[3][0] ), .S(N3) );
  FA_X1 \mult_19/S3_4_30  ( .A(\mult_19/ab[4][30] ), .B(
        \mult_19/CARRYB[3][30] ), .CI(\mult_19/ab[3][31] ), .CO(
        \mult_19/CARRYB[4][30] ), .S(\mult_19/SUMB[4][30] ) );
  FA_X1 \mult_19/S2_4_29  ( .A(\mult_19/ab[4][29] ), .B(
        \mult_19/CARRYB[3][29] ), .CI(\mult_19/SUMB[3][30] ), .CO(
        \mult_19/CARRYB[4][29] ), .S(\mult_19/SUMB[4][29] ) );
  FA_X1 \mult_19/S2_4_28  ( .A(\mult_19/ab[4][28] ), .B(
        \mult_19/CARRYB[3][28] ), .CI(\mult_19/SUMB[3][29] ), .CO(
        \mult_19/CARRYB[4][28] ), .S(\mult_19/SUMB[4][28] ) );
  FA_X1 \mult_19/S2_4_27  ( .A(\mult_19/ab[4][27] ), .B(
        \mult_19/CARRYB[3][27] ), .CI(\mult_19/SUMB[3][28] ), .CO(
        \mult_19/CARRYB[4][27] ), .S(\mult_19/SUMB[4][27] ) );
  FA_X1 \mult_19/S2_4_26  ( .A(\mult_19/ab[4][26] ), .B(
        \mult_19/CARRYB[3][26] ), .CI(\mult_19/SUMB[3][27] ), .CO(
        \mult_19/CARRYB[4][26] ), .S(\mult_19/SUMB[4][26] ) );
  FA_X1 \mult_19/S2_4_25  ( .A(\mult_19/ab[4][25] ), .B(
        \mult_19/CARRYB[3][25] ), .CI(\mult_19/SUMB[3][26] ), .CO(
        \mult_19/CARRYB[4][25] ), .S(\mult_19/SUMB[4][25] ) );
  FA_X1 \mult_19/S2_4_24  ( .A(\mult_19/ab[4][24] ), .B(
        \mult_19/CARRYB[3][24] ), .CI(\mult_19/SUMB[3][25] ), .CO(
        \mult_19/CARRYB[4][24] ), .S(\mult_19/SUMB[4][24] ) );
  FA_X1 \mult_19/S2_4_23  ( .A(\mult_19/ab[4][23] ), .B(
        \mult_19/CARRYB[3][23] ), .CI(\mult_19/SUMB[3][24] ), .CO(
        \mult_19/CARRYB[4][23] ), .S(\mult_19/SUMB[4][23] ) );
  FA_X1 \mult_19/S2_4_22  ( .A(\mult_19/ab[4][22] ), .B(
        \mult_19/CARRYB[3][22] ), .CI(\mult_19/SUMB[3][23] ), .CO(
        \mult_19/CARRYB[4][22] ), .S(\mult_19/SUMB[4][22] ) );
  FA_X1 \mult_19/S2_4_21  ( .A(\mult_19/ab[4][21] ), .B(
        \mult_19/CARRYB[3][21] ), .CI(\mult_19/SUMB[3][22] ), .CO(
        \mult_19/CARRYB[4][21] ), .S(\mult_19/SUMB[4][21] ) );
  FA_X1 \mult_19/S2_4_20  ( .A(\mult_19/ab[4][20] ), .B(
        \mult_19/CARRYB[3][20] ), .CI(\mult_19/SUMB[3][21] ), .CO(
        \mult_19/CARRYB[4][20] ), .S(\mult_19/SUMB[4][20] ) );
  FA_X1 \mult_19/S2_4_19  ( .A(\mult_19/ab[4][19] ), .B(
        \mult_19/CARRYB[3][19] ), .CI(\mult_19/SUMB[3][20] ), .CO(
        \mult_19/CARRYB[4][19] ), .S(\mult_19/SUMB[4][19] ) );
  FA_X1 \mult_19/S2_4_18  ( .A(\mult_19/ab[4][18] ), .B(
        \mult_19/CARRYB[3][18] ), .CI(\mult_19/SUMB[3][19] ), .CO(
        \mult_19/CARRYB[4][18] ), .S(\mult_19/SUMB[4][18] ) );
  FA_X1 \mult_19/S2_4_17  ( .A(\mult_19/ab[4][17] ), .B(
        \mult_19/CARRYB[3][17] ), .CI(\mult_19/SUMB[3][18] ), .CO(
        \mult_19/CARRYB[4][17] ), .S(\mult_19/SUMB[4][17] ) );
  FA_X1 \mult_19/S2_4_16  ( .A(\mult_19/ab[4][16] ), .B(
        \mult_19/CARRYB[3][16] ), .CI(\mult_19/SUMB[3][17] ), .CO(
        \mult_19/CARRYB[4][16] ), .S(\mult_19/SUMB[4][16] ) );
  FA_X1 \mult_19/S2_4_15  ( .A(\mult_19/ab[4][15] ), .B(
        \mult_19/CARRYB[3][15] ), .CI(\mult_19/SUMB[3][16] ), .CO(
        \mult_19/CARRYB[4][15] ), .S(\mult_19/SUMB[4][15] ) );
  FA_X1 \mult_19/S2_4_14  ( .A(\mult_19/ab[4][14] ), .B(
        \mult_19/CARRYB[3][14] ), .CI(\mult_19/SUMB[3][15] ), .CO(
        \mult_19/CARRYB[4][14] ), .S(\mult_19/SUMB[4][14] ) );
  FA_X1 \mult_19/S2_4_13  ( .A(\mult_19/ab[4][13] ), .B(
        \mult_19/CARRYB[3][13] ), .CI(\mult_19/SUMB[3][14] ), .CO(
        \mult_19/CARRYB[4][13] ), .S(\mult_19/SUMB[4][13] ) );
  FA_X1 \mult_19/S2_4_12  ( .A(\mult_19/ab[4][12] ), .B(
        \mult_19/CARRYB[3][12] ), .CI(\mult_19/SUMB[3][13] ), .CO(
        \mult_19/CARRYB[4][12] ), .S(\mult_19/SUMB[4][12] ) );
  FA_X1 \mult_19/S2_4_11  ( .A(\mult_19/ab[4][11] ), .B(
        \mult_19/CARRYB[3][11] ), .CI(\mult_19/SUMB[3][12] ), .CO(
        \mult_19/CARRYB[4][11] ), .S(\mult_19/SUMB[4][11] ) );
  FA_X1 \mult_19/S2_4_10  ( .A(\mult_19/ab[4][10] ), .B(
        \mult_19/CARRYB[3][10] ), .CI(\mult_19/SUMB[3][11] ), .CO(
        \mult_19/CARRYB[4][10] ), .S(\mult_19/SUMB[4][10] ) );
  FA_X1 \mult_19/S2_4_9  ( .A(\mult_19/ab[4][9] ), .B(\mult_19/CARRYB[3][9] ), 
        .CI(\mult_19/SUMB[3][10] ), .CO(\mult_19/CARRYB[4][9] ), .S(
        \mult_19/SUMB[4][9] ) );
  FA_X1 \mult_19/S2_4_8  ( .A(\mult_19/ab[4][8] ), .B(\mult_19/CARRYB[3][8] ), 
        .CI(\mult_19/SUMB[3][9] ), .CO(\mult_19/CARRYB[4][8] ), .S(
        \mult_19/SUMB[4][8] ) );
  FA_X1 \mult_19/S2_4_7  ( .A(\mult_19/ab[4][7] ), .B(\mult_19/CARRYB[3][7] ), 
        .CI(\mult_19/SUMB[3][8] ), .CO(\mult_19/CARRYB[4][7] ), .S(
        \mult_19/SUMB[4][7] ) );
  FA_X1 \mult_19/S2_4_6  ( .A(\mult_19/ab[4][6] ), .B(\mult_19/CARRYB[3][6] ), 
        .CI(\mult_19/SUMB[3][7] ), .CO(\mult_19/CARRYB[4][6] ), .S(
        \mult_19/SUMB[4][6] ) );
  FA_X1 \mult_19/S2_4_5  ( .A(\mult_19/ab[4][5] ), .B(\mult_19/CARRYB[3][5] ), 
        .CI(\mult_19/SUMB[3][6] ), .CO(\mult_19/CARRYB[4][5] ), .S(
        \mult_19/SUMB[4][5] ) );
  FA_X1 \mult_19/S2_4_4  ( .A(\mult_19/ab[4][4] ), .B(\mult_19/CARRYB[3][4] ), 
        .CI(\mult_19/SUMB[3][5] ), .CO(\mult_19/CARRYB[4][4] ), .S(
        \mult_19/SUMB[4][4] ) );
  FA_X1 \mult_19/S2_4_3  ( .A(\mult_19/ab[4][3] ), .B(\mult_19/CARRYB[3][3] ), 
        .CI(\mult_19/SUMB[3][4] ), .CO(\mult_19/CARRYB[4][3] ), .S(
        \mult_19/SUMB[4][3] ) );
  FA_X1 \mult_19/S2_4_2  ( .A(\mult_19/ab[4][2] ), .B(\mult_19/CARRYB[3][2] ), 
        .CI(\mult_19/SUMB[3][3] ), .CO(\mult_19/CARRYB[4][2] ), .S(
        \mult_19/SUMB[4][2] ) );
  FA_X1 \mult_19/S2_4_1  ( .A(\mult_19/ab[4][1] ), .B(\mult_19/CARRYB[3][1] ), 
        .CI(\mult_19/SUMB[3][2] ), .CO(\mult_19/CARRYB[4][1] ), .S(
        \mult_19/SUMB[4][1] ) );
  FA_X1 \mult_19/S1_4_0  ( .A(\mult_19/ab[4][0] ), .B(\mult_19/CARRYB[3][0] ), 
        .CI(\mult_19/SUMB[3][1] ), .CO(\mult_19/CARRYB[4][0] ), .S(N4) );
  FA_X1 \mult_19/S3_5_30  ( .A(\mult_19/ab[5][30] ), .B(
        \mult_19/CARRYB[4][30] ), .CI(\mult_19/ab[4][31] ), .CO(
        \mult_19/CARRYB[5][30] ), .S(\mult_19/SUMB[5][30] ) );
  FA_X1 \mult_19/S2_5_29  ( .A(\mult_19/ab[5][29] ), .B(
        \mult_19/CARRYB[4][29] ), .CI(\mult_19/SUMB[4][30] ), .CO(
        \mult_19/CARRYB[5][29] ), .S(\mult_19/SUMB[5][29] ) );
  FA_X1 \mult_19/S2_5_28  ( .A(\mult_19/ab[5][28] ), .B(
        \mult_19/CARRYB[4][28] ), .CI(\mult_19/SUMB[4][29] ), .CO(
        \mult_19/CARRYB[5][28] ), .S(\mult_19/SUMB[5][28] ) );
  FA_X1 \mult_19/S2_5_27  ( .A(\mult_19/ab[5][27] ), .B(
        \mult_19/CARRYB[4][27] ), .CI(\mult_19/SUMB[4][28] ), .CO(
        \mult_19/CARRYB[5][27] ), .S(\mult_19/SUMB[5][27] ) );
  FA_X1 \mult_19/S2_5_26  ( .A(\mult_19/ab[5][26] ), .B(
        \mult_19/CARRYB[4][26] ), .CI(\mult_19/SUMB[4][27] ), .CO(
        \mult_19/CARRYB[5][26] ), .S(\mult_19/SUMB[5][26] ) );
  FA_X1 \mult_19/S2_5_25  ( .A(\mult_19/ab[5][25] ), .B(
        \mult_19/CARRYB[4][25] ), .CI(\mult_19/SUMB[4][26] ), .CO(
        \mult_19/CARRYB[5][25] ), .S(\mult_19/SUMB[5][25] ) );
  FA_X1 \mult_19/S2_5_24  ( .A(\mult_19/ab[5][24] ), .B(
        \mult_19/CARRYB[4][24] ), .CI(\mult_19/SUMB[4][25] ), .CO(
        \mult_19/CARRYB[5][24] ), .S(\mult_19/SUMB[5][24] ) );
  FA_X1 \mult_19/S2_5_23  ( .A(\mult_19/ab[5][23] ), .B(
        \mult_19/CARRYB[4][23] ), .CI(\mult_19/SUMB[4][24] ), .CO(
        \mult_19/CARRYB[5][23] ), .S(\mult_19/SUMB[5][23] ) );
  FA_X1 \mult_19/S2_5_22  ( .A(\mult_19/ab[5][22] ), .B(
        \mult_19/CARRYB[4][22] ), .CI(\mult_19/SUMB[4][23] ), .CO(
        \mult_19/CARRYB[5][22] ), .S(\mult_19/SUMB[5][22] ) );
  FA_X1 \mult_19/S2_5_21  ( .A(\mult_19/ab[5][21] ), .B(
        \mult_19/CARRYB[4][21] ), .CI(\mult_19/SUMB[4][22] ), .CO(
        \mult_19/CARRYB[5][21] ), .S(\mult_19/SUMB[5][21] ) );
  FA_X1 \mult_19/S2_5_20  ( .A(\mult_19/ab[5][20] ), .B(
        \mult_19/CARRYB[4][20] ), .CI(\mult_19/SUMB[4][21] ), .CO(
        \mult_19/CARRYB[5][20] ), .S(\mult_19/SUMB[5][20] ) );
  FA_X1 \mult_19/S2_5_19  ( .A(\mult_19/ab[5][19] ), .B(
        \mult_19/CARRYB[4][19] ), .CI(\mult_19/SUMB[4][20] ), .CO(
        \mult_19/CARRYB[5][19] ), .S(\mult_19/SUMB[5][19] ) );
  FA_X1 \mult_19/S2_5_18  ( .A(\mult_19/ab[5][18] ), .B(
        \mult_19/CARRYB[4][18] ), .CI(\mult_19/SUMB[4][19] ), .CO(
        \mult_19/CARRYB[5][18] ), .S(\mult_19/SUMB[5][18] ) );
  FA_X1 \mult_19/S2_5_17  ( .A(\mult_19/ab[5][17] ), .B(
        \mult_19/CARRYB[4][17] ), .CI(\mult_19/SUMB[4][18] ), .CO(
        \mult_19/CARRYB[5][17] ), .S(\mult_19/SUMB[5][17] ) );
  FA_X1 \mult_19/S2_5_16  ( .A(\mult_19/ab[5][16] ), .B(
        \mult_19/CARRYB[4][16] ), .CI(\mult_19/SUMB[4][17] ), .CO(
        \mult_19/CARRYB[5][16] ), .S(\mult_19/SUMB[5][16] ) );
  FA_X1 \mult_19/S2_5_15  ( .A(\mult_19/ab[5][15] ), .B(
        \mult_19/CARRYB[4][15] ), .CI(\mult_19/SUMB[4][16] ), .CO(
        \mult_19/CARRYB[5][15] ), .S(\mult_19/SUMB[5][15] ) );
  FA_X1 \mult_19/S2_5_14  ( .A(\mult_19/ab[5][14] ), .B(
        \mult_19/CARRYB[4][14] ), .CI(\mult_19/SUMB[4][15] ), .CO(
        \mult_19/CARRYB[5][14] ), .S(\mult_19/SUMB[5][14] ) );
  FA_X1 \mult_19/S2_5_13  ( .A(\mult_19/ab[5][13] ), .B(
        \mult_19/CARRYB[4][13] ), .CI(\mult_19/SUMB[4][14] ), .CO(
        \mult_19/CARRYB[5][13] ), .S(\mult_19/SUMB[5][13] ) );
  FA_X1 \mult_19/S2_5_12  ( .A(\mult_19/ab[5][12] ), .B(
        \mult_19/CARRYB[4][12] ), .CI(\mult_19/SUMB[4][13] ), .CO(
        \mult_19/CARRYB[5][12] ), .S(\mult_19/SUMB[5][12] ) );
  FA_X1 \mult_19/S2_5_11  ( .A(\mult_19/ab[5][11] ), .B(
        \mult_19/CARRYB[4][11] ), .CI(\mult_19/SUMB[4][12] ), .CO(
        \mult_19/CARRYB[5][11] ), .S(\mult_19/SUMB[5][11] ) );
  FA_X1 \mult_19/S2_5_10  ( .A(\mult_19/ab[5][10] ), .B(
        \mult_19/CARRYB[4][10] ), .CI(\mult_19/SUMB[4][11] ), .CO(
        \mult_19/CARRYB[5][10] ), .S(\mult_19/SUMB[5][10] ) );
  FA_X1 \mult_19/S2_5_9  ( .A(\mult_19/ab[5][9] ), .B(\mult_19/CARRYB[4][9] ), 
        .CI(\mult_19/SUMB[4][10] ), .CO(\mult_19/CARRYB[5][9] ), .S(
        \mult_19/SUMB[5][9] ) );
  FA_X1 \mult_19/S2_5_8  ( .A(\mult_19/ab[5][8] ), .B(\mult_19/CARRYB[4][8] ), 
        .CI(\mult_19/SUMB[4][9] ), .CO(\mult_19/CARRYB[5][8] ), .S(
        \mult_19/SUMB[5][8] ) );
  FA_X1 \mult_19/S2_5_7  ( .A(\mult_19/ab[5][7] ), .B(\mult_19/CARRYB[4][7] ), 
        .CI(\mult_19/SUMB[4][8] ), .CO(\mult_19/CARRYB[5][7] ), .S(
        \mult_19/SUMB[5][7] ) );
  FA_X1 \mult_19/S2_5_6  ( .A(\mult_19/ab[5][6] ), .B(\mult_19/CARRYB[4][6] ), 
        .CI(\mult_19/SUMB[4][7] ), .CO(\mult_19/CARRYB[5][6] ), .S(
        \mult_19/SUMB[5][6] ) );
  FA_X1 \mult_19/S2_5_5  ( .A(\mult_19/ab[5][5] ), .B(\mult_19/CARRYB[4][5] ), 
        .CI(\mult_19/SUMB[4][6] ), .CO(\mult_19/CARRYB[5][5] ), .S(
        \mult_19/SUMB[5][5] ) );
  FA_X1 \mult_19/S2_5_4  ( .A(\mult_19/ab[5][4] ), .B(\mult_19/CARRYB[4][4] ), 
        .CI(\mult_19/SUMB[4][5] ), .CO(\mult_19/CARRYB[5][4] ), .S(
        \mult_19/SUMB[5][4] ) );
  FA_X1 \mult_19/S2_5_3  ( .A(\mult_19/ab[5][3] ), .B(\mult_19/CARRYB[4][3] ), 
        .CI(\mult_19/SUMB[4][4] ), .CO(\mult_19/CARRYB[5][3] ), .S(
        \mult_19/SUMB[5][3] ) );
  FA_X1 \mult_19/S2_5_2  ( .A(\mult_19/ab[5][2] ), .B(\mult_19/CARRYB[4][2] ), 
        .CI(\mult_19/SUMB[4][3] ), .CO(\mult_19/CARRYB[5][2] ), .S(
        \mult_19/SUMB[5][2] ) );
  FA_X1 \mult_19/S2_5_1  ( .A(\mult_19/ab[5][1] ), .B(\mult_19/CARRYB[4][1] ), 
        .CI(\mult_19/SUMB[4][2] ), .CO(\mult_19/CARRYB[5][1] ), .S(
        \mult_19/SUMB[5][1] ) );
  FA_X1 \mult_19/S1_5_0  ( .A(\mult_19/ab[5][0] ), .B(\mult_19/CARRYB[4][0] ), 
        .CI(\mult_19/SUMB[4][1] ), .CO(\mult_19/CARRYB[5][0] ), .S(N5) );
  FA_X1 \mult_19/S3_6_30  ( .A(\mult_19/ab[6][30] ), .B(
        \mult_19/CARRYB[5][30] ), .CI(\mult_19/ab[5][31] ), .CO(
        \mult_19/CARRYB[6][30] ), .S(\mult_19/SUMB[6][30] ) );
  FA_X1 \mult_19/S2_6_29  ( .A(\mult_19/ab[6][29] ), .B(
        \mult_19/CARRYB[5][29] ), .CI(\mult_19/SUMB[5][30] ), .CO(
        \mult_19/CARRYB[6][29] ), .S(\mult_19/SUMB[6][29] ) );
  FA_X1 \mult_19/S2_6_28  ( .A(\mult_19/ab[6][28] ), .B(
        \mult_19/CARRYB[5][28] ), .CI(\mult_19/SUMB[5][29] ), .CO(
        \mult_19/CARRYB[6][28] ), .S(\mult_19/SUMB[6][28] ) );
  FA_X1 \mult_19/S2_6_27  ( .A(\mult_19/ab[6][27] ), .B(
        \mult_19/CARRYB[5][27] ), .CI(\mult_19/SUMB[5][28] ), .CO(
        \mult_19/CARRYB[6][27] ), .S(\mult_19/SUMB[6][27] ) );
  FA_X1 \mult_19/S2_6_26  ( .A(\mult_19/ab[6][26] ), .B(
        \mult_19/CARRYB[5][26] ), .CI(\mult_19/SUMB[5][27] ), .CO(
        \mult_19/CARRYB[6][26] ), .S(\mult_19/SUMB[6][26] ) );
  FA_X1 \mult_19/S2_6_25  ( .A(\mult_19/ab[6][25] ), .B(
        \mult_19/CARRYB[5][25] ), .CI(\mult_19/SUMB[5][26] ), .CO(
        \mult_19/CARRYB[6][25] ), .S(\mult_19/SUMB[6][25] ) );
  FA_X1 \mult_19/S2_6_24  ( .A(\mult_19/ab[6][24] ), .B(
        \mult_19/CARRYB[5][24] ), .CI(\mult_19/SUMB[5][25] ), .CO(
        \mult_19/CARRYB[6][24] ), .S(\mult_19/SUMB[6][24] ) );
  FA_X1 \mult_19/S2_6_23  ( .A(\mult_19/ab[6][23] ), .B(
        \mult_19/CARRYB[5][23] ), .CI(\mult_19/SUMB[5][24] ), .CO(
        \mult_19/CARRYB[6][23] ), .S(\mult_19/SUMB[6][23] ) );
  FA_X1 \mult_19/S2_6_22  ( .A(\mult_19/ab[6][22] ), .B(
        \mult_19/CARRYB[5][22] ), .CI(\mult_19/SUMB[5][23] ), .CO(
        \mult_19/CARRYB[6][22] ), .S(\mult_19/SUMB[6][22] ) );
  FA_X1 \mult_19/S2_6_21  ( .A(\mult_19/ab[6][21] ), .B(
        \mult_19/CARRYB[5][21] ), .CI(\mult_19/SUMB[5][22] ), .CO(
        \mult_19/CARRYB[6][21] ), .S(\mult_19/SUMB[6][21] ) );
  FA_X1 \mult_19/S2_6_20  ( .A(\mult_19/ab[6][20] ), .B(
        \mult_19/CARRYB[5][20] ), .CI(\mult_19/SUMB[5][21] ), .CO(
        \mult_19/CARRYB[6][20] ), .S(\mult_19/SUMB[6][20] ) );
  FA_X1 \mult_19/S2_6_19  ( .A(\mult_19/ab[6][19] ), .B(
        \mult_19/CARRYB[5][19] ), .CI(\mult_19/SUMB[5][20] ), .CO(
        \mult_19/CARRYB[6][19] ), .S(\mult_19/SUMB[6][19] ) );
  FA_X1 \mult_19/S2_6_18  ( .A(\mult_19/ab[6][18] ), .B(
        \mult_19/CARRYB[5][18] ), .CI(\mult_19/SUMB[5][19] ), .CO(
        \mult_19/CARRYB[6][18] ), .S(\mult_19/SUMB[6][18] ) );
  FA_X1 \mult_19/S2_6_17  ( .A(\mult_19/ab[6][17] ), .B(
        \mult_19/CARRYB[5][17] ), .CI(\mult_19/SUMB[5][18] ), .CO(
        \mult_19/CARRYB[6][17] ), .S(\mult_19/SUMB[6][17] ) );
  FA_X1 \mult_19/S2_6_16  ( .A(\mult_19/ab[6][16] ), .B(
        \mult_19/CARRYB[5][16] ), .CI(\mult_19/SUMB[5][17] ), .CO(
        \mult_19/CARRYB[6][16] ), .S(\mult_19/SUMB[6][16] ) );
  FA_X1 \mult_19/S2_6_15  ( .A(\mult_19/ab[6][15] ), .B(
        \mult_19/CARRYB[5][15] ), .CI(\mult_19/SUMB[5][16] ), .CO(
        \mult_19/CARRYB[6][15] ), .S(\mult_19/SUMB[6][15] ) );
  FA_X1 \mult_19/S2_6_14  ( .A(\mult_19/ab[6][14] ), .B(
        \mult_19/CARRYB[5][14] ), .CI(\mult_19/SUMB[5][15] ), .CO(
        \mult_19/CARRYB[6][14] ), .S(\mult_19/SUMB[6][14] ) );
  FA_X1 \mult_19/S2_6_13  ( .A(\mult_19/ab[6][13] ), .B(
        \mult_19/CARRYB[5][13] ), .CI(\mult_19/SUMB[5][14] ), .CO(
        \mult_19/CARRYB[6][13] ), .S(\mult_19/SUMB[6][13] ) );
  FA_X1 \mult_19/S2_6_12  ( .A(\mult_19/ab[6][12] ), .B(
        \mult_19/CARRYB[5][12] ), .CI(\mult_19/SUMB[5][13] ), .CO(
        \mult_19/CARRYB[6][12] ), .S(\mult_19/SUMB[6][12] ) );
  FA_X1 \mult_19/S2_6_11  ( .A(\mult_19/ab[6][11] ), .B(
        \mult_19/CARRYB[5][11] ), .CI(\mult_19/SUMB[5][12] ), .CO(
        \mult_19/CARRYB[6][11] ), .S(\mult_19/SUMB[6][11] ) );
  FA_X1 \mult_19/S2_6_10  ( .A(\mult_19/ab[6][10] ), .B(
        \mult_19/CARRYB[5][10] ), .CI(\mult_19/SUMB[5][11] ), .CO(
        \mult_19/CARRYB[6][10] ), .S(\mult_19/SUMB[6][10] ) );
  FA_X1 \mult_19/S2_6_9  ( .A(\mult_19/ab[6][9] ), .B(\mult_19/CARRYB[5][9] ), 
        .CI(\mult_19/SUMB[5][10] ), .CO(\mult_19/CARRYB[6][9] ), .S(
        \mult_19/SUMB[6][9] ) );
  FA_X1 \mult_19/S2_6_8  ( .A(\mult_19/ab[6][8] ), .B(\mult_19/CARRYB[5][8] ), 
        .CI(\mult_19/SUMB[5][9] ), .CO(\mult_19/CARRYB[6][8] ), .S(
        \mult_19/SUMB[6][8] ) );
  FA_X1 \mult_19/S2_6_7  ( .A(\mult_19/ab[6][7] ), .B(\mult_19/CARRYB[5][7] ), 
        .CI(\mult_19/SUMB[5][8] ), .CO(\mult_19/CARRYB[6][7] ), .S(
        \mult_19/SUMB[6][7] ) );
  FA_X1 \mult_19/S2_6_6  ( .A(\mult_19/ab[6][6] ), .B(\mult_19/CARRYB[5][6] ), 
        .CI(\mult_19/SUMB[5][7] ), .CO(\mult_19/CARRYB[6][6] ), .S(
        \mult_19/SUMB[6][6] ) );
  FA_X1 \mult_19/S2_6_5  ( .A(\mult_19/ab[6][5] ), .B(\mult_19/CARRYB[5][5] ), 
        .CI(\mult_19/SUMB[5][6] ), .CO(\mult_19/CARRYB[6][5] ), .S(
        \mult_19/SUMB[6][5] ) );
  FA_X1 \mult_19/S2_6_4  ( .A(\mult_19/ab[6][4] ), .B(\mult_19/CARRYB[5][4] ), 
        .CI(\mult_19/SUMB[5][5] ), .CO(\mult_19/CARRYB[6][4] ), .S(
        \mult_19/SUMB[6][4] ) );
  FA_X1 \mult_19/S2_6_3  ( .A(\mult_19/ab[6][3] ), .B(\mult_19/CARRYB[5][3] ), 
        .CI(\mult_19/SUMB[5][4] ), .CO(\mult_19/CARRYB[6][3] ), .S(
        \mult_19/SUMB[6][3] ) );
  FA_X1 \mult_19/S2_6_2  ( .A(\mult_19/ab[6][2] ), .B(\mult_19/CARRYB[5][2] ), 
        .CI(\mult_19/SUMB[5][3] ), .CO(\mult_19/CARRYB[6][2] ), .S(
        \mult_19/SUMB[6][2] ) );
  FA_X1 \mult_19/S2_6_1  ( .A(\mult_19/ab[6][1] ), .B(\mult_19/CARRYB[5][1] ), 
        .CI(\mult_19/SUMB[5][2] ), .CO(\mult_19/CARRYB[6][1] ), .S(
        \mult_19/SUMB[6][1] ) );
  FA_X1 \mult_19/S1_6_0  ( .A(\mult_19/ab[6][0] ), .B(\mult_19/CARRYB[5][0] ), 
        .CI(\mult_19/SUMB[5][1] ), .CO(\mult_19/CARRYB[6][0] ), .S(N6) );
  FA_X1 \mult_19/S3_7_30  ( .A(\mult_19/ab[7][30] ), .B(
        \mult_19/CARRYB[6][30] ), .CI(\mult_19/ab[6][31] ), .CO(
        \mult_19/CARRYB[7][30] ), .S(\mult_19/SUMB[7][30] ) );
  FA_X1 \mult_19/S2_7_29  ( .A(\mult_19/ab[7][29] ), .B(
        \mult_19/CARRYB[6][29] ), .CI(\mult_19/SUMB[6][30] ), .CO(
        \mult_19/CARRYB[7][29] ), .S(\mult_19/SUMB[7][29] ) );
  FA_X1 \mult_19/S2_7_28  ( .A(\mult_19/ab[7][28] ), .B(
        \mult_19/CARRYB[6][28] ), .CI(\mult_19/SUMB[6][29] ), .CO(
        \mult_19/CARRYB[7][28] ), .S(\mult_19/SUMB[7][28] ) );
  FA_X1 \mult_19/S2_7_27  ( .A(\mult_19/ab[7][27] ), .B(
        \mult_19/CARRYB[6][27] ), .CI(\mult_19/SUMB[6][28] ), .CO(
        \mult_19/CARRYB[7][27] ), .S(\mult_19/SUMB[7][27] ) );
  FA_X1 \mult_19/S2_7_26  ( .A(\mult_19/ab[7][26] ), .B(
        \mult_19/CARRYB[6][26] ), .CI(\mult_19/SUMB[6][27] ), .CO(
        \mult_19/CARRYB[7][26] ), .S(\mult_19/SUMB[7][26] ) );
  FA_X1 \mult_19/S2_7_25  ( .A(\mult_19/ab[7][25] ), .B(
        \mult_19/CARRYB[6][25] ), .CI(\mult_19/SUMB[6][26] ), .CO(
        \mult_19/CARRYB[7][25] ), .S(\mult_19/SUMB[7][25] ) );
  FA_X1 \mult_19/S2_7_24  ( .A(\mult_19/ab[7][24] ), .B(
        \mult_19/CARRYB[6][24] ), .CI(\mult_19/SUMB[6][25] ), .CO(
        \mult_19/CARRYB[7][24] ), .S(\mult_19/SUMB[7][24] ) );
  FA_X1 \mult_19/S2_7_23  ( .A(\mult_19/ab[7][23] ), .B(
        \mult_19/CARRYB[6][23] ), .CI(\mult_19/SUMB[6][24] ), .CO(
        \mult_19/CARRYB[7][23] ), .S(\mult_19/SUMB[7][23] ) );
  FA_X1 \mult_19/S2_7_22  ( .A(\mult_19/ab[7][22] ), .B(
        \mult_19/CARRYB[6][22] ), .CI(\mult_19/SUMB[6][23] ), .CO(
        \mult_19/CARRYB[7][22] ), .S(\mult_19/SUMB[7][22] ) );
  FA_X1 \mult_19/S2_7_21  ( .A(\mult_19/ab[7][21] ), .B(
        \mult_19/CARRYB[6][21] ), .CI(\mult_19/SUMB[6][22] ), .CO(
        \mult_19/CARRYB[7][21] ), .S(\mult_19/SUMB[7][21] ) );
  FA_X1 \mult_19/S2_7_20  ( .A(\mult_19/ab[7][20] ), .B(
        \mult_19/CARRYB[6][20] ), .CI(\mult_19/SUMB[6][21] ), .CO(
        \mult_19/CARRYB[7][20] ), .S(\mult_19/SUMB[7][20] ) );
  FA_X1 \mult_19/S2_7_19  ( .A(\mult_19/ab[7][19] ), .B(
        \mult_19/CARRYB[6][19] ), .CI(\mult_19/SUMB[6][20] ), .CO(
        \mult_19/CARRYB[7][19] ), .S(\mult_19/SUMB[7][19] ) );
  FA_X1 \mult_19/S2_7_18  ( .A(\mult_19/ab[7][18] ), .B(
        \mult_19/CARRYB[6][18] ), .CI(\mult_19/SUMB[6][19] ), .CO(
        \mult_19/CARRYB[7][18] ), .S(\mult_19/SUMB[7][18] ) );
  FA_X1 \mult_19/S2_7_17  ( .A(\mult_19/ab[7][17] ), .B(
        \mult_19/CARRYB[6][17] ), .CI(\mult_19/SUMB[6][18] ), .CO(
        \mult_19/CARRYB[7][17] ), .S(\mult_19/SUMB[7][17] ) );
  FA_X1 \mult_19/S2_7_16  ( .A(\mult_19/ab[7][16] ), .B(
        \mult_19/CARRYB[6][16] ), .CI(\mult_19/SUMB[6][17] ), .CO(
        \mult_19/CARRYB[7][16] ), .S(\mult_19/SUMB[7][16] ) );
  FA_X1 \mult_19/S2_7_15  ( .A(\mult_19/ab[7][15] ), .B(
        \mult_19/CARRYB[6][15] ), .CI(\mult_19/SUMB[6][16] ), .CO(
        \mult_19/CARRYB[7][15] ), .S(\mult_19/SUMB[7][15] ) );
  FA_X1 \mult_19/S2_7_14  ( .A(\mult_19/ab[7][14] ), .B(
        \mult_19/CARRYB[6][14] ), .CI(\mult_19/SUMB[6][15] ), .CO(
        \mult_19/CARRYB[7][14] ), .S(\mult_19/SUMB[7][14] ) );
  FA_X1 \mult_19/S2_7_13  ( .A(\mult_19/ab[7][13] ), .B(
        \mult_19/CARRYB[6][13] ), .CI(\mult_19/SUMB[6][14] ), .CO(
        \mult_19/CARRYB[7][13] ), .S(\mult_19/SUMB[7][13] ) );
  FA_X1 \mult_19/S2_7_12  ( .A(\mult_19/ab[7][12] ), .B(
        \mult_19/CARRYB[6][12] ), .CI(\mult_19/SUMB[6][13] ), .CO(
        \mult_19/CARRYB[7][12] ), .S(\mult_19/SUMB[7][12] ) );
  FA_X1 \mult_19/S2_7_11  ( .A(\mult_19/ab[7][11] ), .B(
        \mult_19/CARRYB[6][11] ), .CI(\mult_19/SUMB[6][12] ), .CO(
        \mult_19/CARRYB[7][11] ), .S(\mult_19/SUMB[7][11] ) );
  FA_X1 \mult_19/S2_7_10  ( .A(\mult_19/ab[7][10] ), .B(
        \mult_19/CARRYB[6][10] ), .CI(\mult_19/SUMB[6][11] ), .CO(
        \mult_19/CARRYB[7][10] ), .S(\mult_19/SUMB[7][10] ) );
  FA_X1 \mult_19/S2_7_9  ( .A(\mult_19/ab[7][9] ), .B(\mult_19/CARRYB[6][9] ), 
        .CI(\mult_19/SUMB[6][10] ), .CO(\mult_19/CARRYB[7][9] ), .S(
        \mult_19/SUMB[7][9] ) );
  FA_X1 \mult_19/S2_7_8  ( .A(\mult_19/ab[7][8] ), .B(\mult_19/CARRYB[6][8] ), 
        .CI(\mult_19/SUMB[6][9] ), .CO(\mult_19/CARRYB[7][8] ), .S(
        \mult_19/SUMB[7][8] ) );
  FA_X1 \mult_19/S2_7_7  ( .A(\mult_19/ab[7][7] ), .B(\mult_19/CARRYB[6][7] ), 
        .CI(\mult_19/SUMB[6][8] ), .CO(\mult_19/CARRYB[7][7] ), .S(
        \mult_19/SUMB[7][7] ) );
  FA_X1 \mult_19/S2_7_6  ( .A(\mult_19/ab[7][6] ), .B(\mult_19/CARRYB[6][6] ), 
        .CI(\mult_19/SUMB[6][7] ), .CO(\mult_19/CARRYB[7][6] ), .S(
        \mult_19/SUMB[7][6] ) );
  FA_X1 \mult_19/S2_7_5  ( .A(\mult_19/ab[7][5] ), .B(\mult_19/CARRYB[6][5] ), 
        .CI(\mult_19/SUMB[6][6] ), .CO(\mult_19/CARRYB[7][5] ), .S(
        \mult_19/SUMB[7][5] ) );
  FA_X1 \mult_19/S2_7_4  ( .A(\mult_19/ab[7][4] ), .B(\mult_19/CARRYB[6][4] ), 
        .CI(\mult_19/SUMB[6][5] ), .CO(\mult_19/CARRYB[7][4] ), .S(
        \mult_19/SUMB[7][4] ) );
  FA_X1 \mult_19/S2_7_3  ( .A(\mult_19/ab[7][3] ), .B(\mult_19/CARRYB[6][3] ), 
        .CI(\mult_19/SUMB[6][4] ), .CO(\mult_19/CARRYB[7][3] ), .S(
        \mult_19/SUMB[7][3] ) );
  FA_X1 \mult_19/S2_7_2  ( .A(\mult_19/ab[7][2] ), .B(\mult_19/CARRYB[6][2] ), 
        .CI(\mult_19/SUMB[6][3] ), .CO(\mult_19/CARRYB[7][2] ), .S(
        \mult_19/SUMB[7][2] ) );
  FA_X1 \mult_19/S2_7_1  ( .A(\mult_19/ab[7][1] ), .B(\mult_19/CARRYB[6][1] ), 
        .CI(\mult_19/SUMB[6][2] ), .CO(\mult_19/CARRYB[7][1] ), .S(
        \mult_19/SUMB[7][1] ) );
  FA_X1 \mult_19/S1_7_0  ( .A(\mult_19/ab[7][0] ), .B(\mult_19/CARRYB[6][0] ), 
        .CI(\mult_19/SUMB[6][1] ), .CO(\mult_19/CARRYB[7][0] ), .S(N7) );
  FA_X1 \mult_19/S3_8_30  ( .A(\mult_19/ab[8][30] ), .B(
        \mult_19/CARRYB[7][30] ), .CI(\mult_19/ab[7][31] ), .CO(
        \mult_19/CARRYB[8][30] ), .S(\mult_19/SUMB[8][30] ) );
  FA_X1 \mult_19/S2_8_29  ( .A(\mult_19/ab[8][29] ), .B(
        \mult_19/CARRYB[7][29] ), .CI(\mult_19/SUMB[7][30] ), .CO(
        \mult_19/CARRYB[8][29] ), .S(\mult_19/SUMB[8][29] ) );
  FA_X1 \mult_19/S2_8_28  ( .A(\mult_19/ab[8][28] ), .B(
        \mult_19/CARRYB[7][28] ), .CI(\mult_19/SUMB[7][29] ), .CO(
        \mult_19/CARRYB[8][28] ), .S(\mult_19/SUMB[8][28] ) );
  FA_X1 \mult_19/S2_8_27  ( .A(\mult_19/ab[8][27] ), .B(
        \mult_19/CARRYB[7][27] ), .CI(\mult_19/SUMB[7][28] ), .CO(
        \mult_19/CARRYB[8][27] ), .S(\mult_19/SUMB[8][27] ) );
  FA_X1 \mult_19/S2_8_26  ( .A(\mult_19/ab[8][26] ), .B(
        \mult_19/CARRYB[7][26] ), .CI(\mult_19/SUMB[7][27] ), .CO(
        \mult_19/CARRYB[8][26] ), .S(\mult_19/SUMB[8][26] ) );
  FA_X1 \mult_19/S2_8_25  ( .A(\mult_19/ab[8][25] ), .B(
        \mult_19/CARRYB[7][25] ), .CI(\mult_19/SUMB[7][26] ), .CO(
        \mult_19/CARRYB[8][25] ), .S(\mult_19/SUMB[8][25] ) );
  FA_X1 \mult_19/S2_8_24  ( .A(\mult_19/ab[8][24] ), .B(
        \mult_19/CARRYB[7][24] ), .CI(\mult_19/SUMB[7][25] ), .CO(
        \mult_19/CARRYB[8][24] ), .S(\mult_19/SUMB[8][24] ) );
  FA_X1 \mult_19/S2_8_23  ( .A(\mult_19/ab[8][23] ), .B(
        \mult_19/CARRYB[7][23] ), .CI(\mult_19/SUMB[7][24] ), .CO(
        \mult_19/CARRYB[8][23] ), .S(\mult_19/SUMB[8][23] ) );
  FA_X1 \mult_19/S2_8_22  ( .A(\mult_19/ab[8][22] ), .B(
        \mult_19/CARRYB[7][22] ), .CI(\mult_19/SUMB[7][23] ), .CO(
        \mult_19/CARRYB[8][22] ), .S(\mult_19/SUMB[8][22] ) );
  FA_X1 \mult_19/S2_8_21  ( .A(\mult_19/ab[8][21] ), .B(
        \mult_19/CARRYB[7][21] ), .CI(\mult_19/SUMB[7][22] ), .CO(
        \mult_19/CARRYB[8][21] ), .S(\mult_19/SUMB[8][21] ) );
  FA_X1 \mult_19/S2_8_20  ( .A(\mult_19/ab[8][20] ), .B(
        \mult_19/CARRYB[7][20] ), .CI(\mult_19/SUMB[7][21] ), .CO(
        \mult_19/CARRYB[8][20] ), .S(\mult_19/SUMB[8][20] ) );
  FA_X1 \mult_19/S2_8_19  ( .A(\mult_19/ab[8][19] ), .B(
        \mult_19/CARRYB[7][19] ), .CI(\mult_19/SUMB[7][20] ), .CO(
        \mult_19/CARRYB[8][19] ), .S(\mult_19/SUMB[8][19] ) );
  FA_X1 \mult_19/S2_8_18  ( .A(\mult_19/ab[8][18] ), .B(
        \mult_19/CARRYB[7][18] ), .CI(\mult_19/SUMB[7][19] ), .CO(
        \mult_19/CARRYB[8][18] ), .S(\mult_19/SUMB[8][18] ) );
  FA_X1 \mult_19/S2_8_17  ( .A(\mult_19/ab[8][17] ), .B(
        \mult_19/CARRYB[7][17] ), .CI(\mult_19/SUMB[7][18] ), .CO(
        \mult_19/CARRYB[8][17] ), .S(\mult_19/SUMB[8][17] ) );
  FA_X1 \mult_19/S2_8_16  ( .A(\mult_19/ab[8][16] ), .B(
        \mult_19/CARRYB[7][16] ), .CI(\mult_19/SUMB[7][17] ), .CO(
        \mult_19/CARRYB[8][16] ), .S(\mult_19/SUMB[8][16] ) );
  FA_X1 \mult_19/S2_8_15  ( .A(\mult_19/ab[8][15] ), .B(
        \mult_19/CARRYB[7][15] ), .CI(\mult_19/SUMB[7][16] ), .CO(
        \mult_19/CARRYB[8][15] ), .S(\mult_19/SUMB[8][15] ) );
  FA_X1 \mult_19/S2_8_14  ( .A(\mult_19/ab[8][14] ), .B(
        \mult_19/CARRYB[7][14] ), .CI(\mult_19/SUMB[7][15] ), .CO(
        \mult_19/CARRYB[8][14] ), .S(\mult_19/SUMB[8][14] ) );
  FA_X1 \mult_19/S2_8_13  ( .A(\mult_19/ab[8][13] ), .B(
        \mult_19/CARRYB[7][13] ), .CI(\mult_19/SUMB[7][14] ), .CO(
        \mult_19/CARRYB[8][13] ), .S(\mult_19/SUMB[8][13] ) );
  FA_X1 \mult_19/S2_8_12  ( .A(\mult_19/ab[8][12] ), .B(
        \mult_19/CARRYB[7][12] ), .CI(\mult_19/SUMB[7][13] ), .CO(
        \mult_19/CARRYB[8][12] ), .S(\mult_19/SUMB[8][12] ) );
  FA_X1 \mult_19/S2_8_11  ( .A(\mult_19/ab[8][11] ), .B(
        \mult_19/CARRYB[7][11] ), .CI(\mult_19/SUMB[7][12] ), .CO(
        \mult_19/CARRYB[8][11] ), .S(\mult_19/SUMB[8][11] ) );
  FA_X1 \mult_19/S2_8_10  ( .A(\mult_19/ab[8][10] ), .B(
        \mult_19/CARRYB[7][10] ), .CI(\mult_19/SUMB[7][11] ), .CO(
        \mult_19/CARRYB[8][10] ), .S(\mult_19/SUMB[8][10] ) );
  FA_X1 \mult_19/S2_8_9  ( .A(\mult_19/ab[8][9] ), .B(\mult_19/CARRYB[7][9] ), 
        .CI(\mult_19/SUMB[7][10] ), .CO(\mult_19/CARRYB[8][9] ), .S(
        \mult_19/SUMB[8][9] ) );
  FA_X1 \mult_19/S2_8_8  ( .A(\mult_19/ab[8][8] ), .B(\mult_19/CARRYB[7][8] ), 
        .CI(\mult_19/SUMB[7][9] ), .CO(\mult_19/CARRYB[8][8] ), .S(
        \mult_19/SUMB[8][8] ) );
  FA_X1 \mult_19/S2_8_7  ( .A(\mult_19/ab[8][7] ), .B(\mult_19/CARRYB[7][7] ), 
        .CI(\mult_19/SUMB[7][8] ), .CO(\mult_19/CARRYB[8][7] ), .S(
        \mult_19/SUMB[8][7] ) );
  FA_X1 \mult_19/S2_8_6  ( .A(\mult_19/ab[8][6] ), .B(\mult_19/CARRYB[7][6] ), 
        .CI(\mult_19/SUMB[7][7] ), .CO(\mult_19/CARRYB[8][6] ), .S(
        \mult_19/SUMB[8][6] ) );
  FA_X1 \mult_19/S2_8_5  ( .A(\mult_19/ab[8][5] ), .B(\mult_19/CARRYB[7][5] ), 
        .CI(\mult_19/SUMB[7][6] ), .CO(\mult_19/CARRYB[8][5] ), .S(
        \mult_19/SUMB[8][5] ) );
  FA_X1 \mult_19/S2_8_4  ( .A(\mult_19/ab[8][4] ), .B(\mult_19/CARRYB[7][4] ), 
        .CI(\mult_19/SUMB[7][5] ), .CO(\mult_19/CARRYB[8][4] ), .S(
        \mult_19/SUMB[8][4] ) );
  FA_X1 \mult_19/S2_8_3  ( .A(\mult_19/ab[8][3] ), .B(\mult_19/CARRYB[7][3] ), 
        .CI(\mult_19/SUMB[7][4] ), .CO(\mult_19/CARRYB[8][3] ), .S(
        \mult_19/SUMB[8][3] ) );
  FA_X1 \mult_19/S2_8_2  ( .A(\mult_19/ab[8][2] ), .B(\mult_19/CARRYB[7][2] ), 
        .CI(\mult_19/SUMB[7][3] ), .CO(\mult_19/CARRYB[8][2] ), .S(
        \mult_19/SUMB[8][2] ) );
  FA_X1 \mult_19/S2_8_1  ( .A(\mult_19/ab[8][1] ), .B(\mult_19/CARRYB[7][1] ), 
        .CI(\mult_19/SUMB[7][2] ), .CO(\mult_19/CARRYB[8][1] ), .S(
        \mult_19/SUMB[8][1] ) );
  FA_X1 \mult_19/S1_8_0  ( .A(\mult_19/ab[8][0] ), .B(\mult_19/CARRYB[7][0] ), 
        .CI(\mult_19/SUMB[7][1] ), .CO(\mult_19/CARRYB[8][0] ), .S(N8) );
  FA_X1 \mult_19/S3_9_30  ( .A(\mult_19/ab[9][30] ), .B(
        \mult_19/CARRYB[8][30] ), .CI(\mult_19/ab[8][31] ), .CO(
        \mult_19/CARRYB[9][30] ), .S(\mult_19/SUMB[9][30] ) );
  FA_X1 \mult_19/S2_9_29  ( .A(\mult_19/ab[9][29] ), .B(
        \mult_19/CARRYB[8][29] ), .CI(\mult_19/SUMB[8][30] ), .CO(
        \mult_19/CARRYB[9][29] ), .S(\mult_19/SUMB[9][29] ) );
  FA_X1 \mult_19/S2_9_28  ( .A(\mult_19/ab[9][28] ), .B(
        \mult_19/CARRYB[8][28] ), .CI(\mult_19/SUMB[8][29] ), .CO(
        \mult_19/CARRYB[9][28] ), .S(\mult_19/SUMB[9][28] ) );
  FA_X1 \mult_19/S2_9_27  ( .A(\mult_19/ab[9][27] ), .B(
        \mult_19/CARRYB[8][27] ), .CI(\mult_19/SUMB[8][28] ), .CO(
        \mult_19/CARRYB[9][27] ), .S(\mult_19/SUMB[9][27] ) );
  FA_X1 \mult_19/S2_9_26  ( .A(\mult_19/ab[9][26] ), .B(
        \mult_19/CARRYB[8][26] ), .CI(\mult_19/SUMB[8][27] ), .CO(
        \mult_19/CARRYB[9][26] ), .S(\mult_19/SUMB[9][26] ) );
  FA_X1 \mult_19/S2_9_25  ( .A(\mult_19/ab[9][25] ), .B(
        \mult_19/CARRYB[8][25] ), .CI(\mult_19/SUMB[8][26] ), .CO(
        \mult_19/CARRYB[9][25] ), .S(\mult_19/SUMB[9][25] ) );
  FA_X1 \mult_19/S2_9_24  ( .A(\mult_19/ab[9][24] ), .B(
        \mult_19/CARRYB[8][24] ), .CI(\mult_19/SUMB[8][25] ), .CO(
        \mult_19/CARRYB[9][24] ), .S(\mult_19/SUMB[9][24] ) );
  FA_X1 \mult_19/S2_9_23  ( .A(\mult_19/ab[9][23] ), .B(
        \mult_19/CARRYB[8][23] ), .CI(\mult_19/SUMB[8][24] ), .CO(
        \mult_19/CARRYB[9][23] ), .S(\mult_19/SUMB[9][23] ) );
  FA_X1 \mult_19/S2_9_22  ( .A(\mult_19/ab[9][22] ), .B(
        \mult_19/CARRYB[8][22] ), .CI(\mult_19/SUMB[8][23] ), .CO(
        \mult_19/CARRYB[9][22] ), .S(\mult_19/SUMB[9][22] ) );
  FA_X1 \mult_19/S2_9_21  ( .A(\mult_19/ab[9][21] ), .B(
        \mult_19/CARRYB[8][21] ), .CI(\mult_19/SUMB[8][22] ), .CO(
        \mult_19/CARRYB[9][21] ), .S(\mult_19/SUMB[9][21] ) );
  FA_X1 \mult_19/S2_9_20  ( .A(\mult_19/ab[9][20] ), .B(
        \mult_19/CARRYB[8][20] ), .CI(\mult_19/SUMB[8][21] ), .CO(
        \mult_19/CARRYB[9][20] ), .S(\mult_19/SUMB[9][20] ) );
  FA_X1 \mult_19/S2_9_19  ( .A(\mult_19/ab[9][19] ), .B(
        \mult_19/CARRYB[8][19] ), .CI(\mult_19/SUMB[8][20] ), .CO(
        \mult_19/CARRYB[9][19] ), .S(\mult_19/SUMB[9][19] ) );
  FA_X1 \mult_19/S2_9_18  ( .A(\mult_19/ab[9][18] ), .B(
        \mult_19/CARRYB[8][18] ), .CI(\mult_19/SUMB[8][19] ), .CO(
        \mult_19/CARRYB[9][18] ), .S(\mult_19/SUMB[9][18] ) );
  FA_X1 \mult_19/S2_9_17  ( .A(\mult_19/ab[9][17] ), .B(
        \mult_19/CARRYB[8][17] ), .CI(\mult_19/SUMB[8][18] ), .CO(
        \mult_19/CARRYB[9][17] ), .S(\mult_19/SUMB[9][17] ) );
  FA_X1 \mult_19/S2_9_16  ( .A(\mult_19/ab[9][16] ), .B(
        \mult_19/CARRYB[8][16] ), .CI(\mult_19/SUMB[8][17] ), .CO(
        \mult_19/CARRYB[9][16] ), .S(\mult_19/SUMB[9][16] ) );
  FA_X1 \mult_19/S2_9_15  ( .A(\mult_19/ab[9][15] ), .B(
        \mult_19/CARRYB[8][15] ), .CI(\mult_19/SUMB[8][16] ), .CO(
        \mult_19/CARRYB[9][15] ), .S(\mult_19/SUMB[9][15] ) );
  FA_X1 \mult_19/S2_9_14  ( .A(\mult_19/ab[9][14] ), .B(
        \mult_19/CARRYB[8][14] ), .CI(\mult_19/SUMB[8][15] ), .CO(
        \mult_19/CARRYB[9][14] ), .S(\mult_19/SUMB[9][14] ) );
  FA_X1 \mult_19/S2_9_13  ( .A(\mult_19/ab[9][13] ), .B(
        \mult_19/CARRYB[8][13] ), .CI(\mult_19/SUMB[8][14] ), .CO(
        \mult_19/CARRYB[9][13] ), .S(\mult_19/SUMB[9][13] ) );
  FA_X1 \mult_19/S2_9_12  ( .A(\mult_19/ab[9][12] ), .B(
        \mult_19/CARRYB[8][12] ), .CI(\mult_19/SUMB[8][13] ), .CO(
        \mult_19/CARRYB[9][12] ), .S(\mult_19/SUMB[9][12] ) );
  FA_X1 \mult_19/S2_9_11  ( .A(\mult_19/ab[9][11] ), .B(
        \mult_19/CARRYB[8][11] ), .CI(\mult_19/SUMB[8][12] ), .CO(
        \mult_19/CARRYB[9][11] ), .S(\mult_19/SUMB[9][11] ) );
  FA_X1 \mult_19/S2_9_10  ( .A(\mult_19/ab[9][10] ), .B(
        \mult_19/CARRYB[8][10] ), .CI(\mult_19/SUMB[8][11] ), .CO(
        \mult_19/CARRYB[9][10] ), .S(\mult_19/SUMB[9][10] ) );
  FA_X1 \mult_19/S2_9_9  ( .A(\mult_19/ab[9][9] ), .B(\mult_19/CARRYB[8][9] ), 
        .CI(\mult_19/SUMB[8][10] ), .CO(\mult_19/CARRYB[9][9] ), .S(
        \mult_19/SUMB[9][9] ) );
  FA_X1 \mult_19/S2_9_8  ( .A(\mult_19/ab[9][8] ), .B(\mult_19/CARRYB[8][8] ), 
        .CI(\mult_19/SUMB[8][9] ), .CO(\mult_19/CARRYB[9][8] ), .S(
        \mult_19/SUMB[9][8] ) );
  FA_X1 \mult_19/S2_9_7  ( .A(\mult_19/ab[9][7] ), .B(\mult_19/CARRYB[8][7] ), 
        .CI(\mult_19/SUMB[8][8] ), .CO(\mult_19/CARRYB[9][7] ), .S(
        \mult_19/SUMB[9][7] ) );
  FA_X1 \mult_19/S2_9_6  ( .A(\mult_19/ab[9][6] ), .B(\mult_19/CARRYB[8][6] ), 
        .CI(\mult_19/SUMB[8][7] ), .CO(\mult_19/CARRYB[9][6] ), .S(
        \mult_19/SUMB[9][6] ) );
  FA_X1 \mult_19/S2_9_5  ( .A(\mult_19/ab[9][5] ), .B(\mult_19/CARRYB[8][5] ), 
        .CI(\mult_19/SUMB[8][6] ), .CO(\mult_19/CARRYB[9][5] ), .S(
        \mult_19/SUMB[9][5] ) );
  FA_X1 \mult_19/S2_9_4  ( .A(\mult_19/ab[9][4] ), .B(\mult_19/CARRYB[8][4] ), 
        .CI(\mult_19/SUMB[8][5] ), .CO(\mult_19/CARRYB[9][4] ), .S(
        \mult_19/SUMB[9][4] ) );
  FA_X1 \mult_19/S2_9_3  ( .A(\mult_19/ab[9][3] ), .B(\mult_19/CARRYB[8][3] ), 
        .CI(\mult_19/SUMB[8][4] ), .CO(\mult_19/CARRYB[9][3] ), .S(
        \mult_19/SUMB[9][3] ) );
  FA_X1 \mult_19/S2_9_2  ( .A(\mult_19/ab[9][2] ), .B(\mult_19/CARRYB[8][2] ), 
        .CI(\mult_19/SUMB[8][3] ), .CO(\mult_19/CARRYB[9][2] ), .S(
        \mult_19/SUMB[9][2] ) );
  FA_X1 \mult_19/S2_9_1  ( .A(\mult_19/ab[9][1] ), .B(\mult_19/CARRYB[8][1] ), 
        .CI(\mult_19/SUMB[8][2] ), .CO(\mult_19/CARRYB[9][1] ), .S(
        \mult_19/SUMB[9][1] ) );
  FA_X1 \mult_19/S1_9_0  ( .A(\mult_19/ab[9][0] ), .B(\mult_19/CARRYB[8][0] ), 
        .CI(\mult_19/SUMB[8][1] ), .CO(\mult_19/CARRYB[9][0] ), .S(N9) );
  FA_X1 \mult_19/S3_10_30  ( .A(\mult_19/ab[10][30] ), .B(
        \mult_19/CARRYB[9][30] ), .CI(\mult_19/ab[9][31] ), .CO(
        \mult_19/CARRYB[10][30] ), .S(\mult_19/SUMB[10][30] ) );
  FA_X1 \mult_19/S2_10_29  ( .A(\mult_19/ab[10][29] ), .B(
        \mult_19/CARRYB[9][29] ), .CI(\mult_19/SUMB[9][30] ), .CO(
        \mult_19/CARRYB[10][29] ), .S(\mult_19/SUMB[10][29] ) );
  FA_X1 \mult_19/S2_10_28  ( .A(\mult_19/ab[10][28] ), .B(
        \mult_19/CARRYB[9][28] ), .CI(\mult_19/SUMB[9][29] ), .CO(
        \mult_19/CARRYB[10][28] ), .S(\mult_19/SUMB[10][28] ) );
  FA_X1 \mult_19/S2_10_27  ( .A(\mult_19/ab[10][27] ), .B(
        \mult_19/CARRYB[9][27] ), .CI(\mult_19/SUMB[9][28] ), .CO(
        \mult_19/CARRYB[10][27] ), .S(\mult_19/SUMB[10][27] ) );
  FA_X1 \mult_19/S2_10_26  ( .A(\mult_19/ab[10][26] ), .B(
        \mult_19/CARRYB[9][26] ), .CI(\mult_19/SUMB[9][27] ), .CO(
        \mult_19/CARRYB[10][26] ), .S(\mult_19/SUMB[10][26] ) );
  FA_X1 \mult_19/S2_10_25  ( .A(\mult_19/ab[10][25] ), .B(
        \mult_19/CARRYB[9][25] ), .CI(\mult_19/SUMB[9][26] ), .CO(
        \mult_19/CARRYB[10][25] ), .S(\mult_19/SUMB[10][25] ) );
  FA_X1 \mult_19/S2_10_24  ( .A(\mult_19/ab[10][24] ), .B(
        \mult_19/CARRYB[9][24] ), .CI(\mult_19/SUMB[9][25] ), .CO(
        \mult_19/CARRYB[10][24] ), .S(\mult_19/SUMB[10][24] ) );
  FA_X1 \mult_19/S2_10_23  ( .A(\mult_19/ab[10][23] ), .B(
        \mult_19/CARRYB[9][23] ), .CI(\mult_19/SUMB[9][24] ), .CO(
        \mult_19/CARRYB[10][23] ), .S(\mult_19/SUMB[10][23] ) );
  FA_X1 \mult_19/S2_10_22  ( .A(\mult_19/ab[10][22] ), .B(
        \mult_19/CARRYB[9][22] ), .CI(\mult_19/SUMB[9][23] ), .CO(
        \mult_19/CARRYB[10][22] ), .S(\mult_19/SUMB[10][22] ) );
  FA_X1 \mult_19/S2_10_21  ( .A(\mult_19/ab[10][21] ), .B(
        \mult_19/CARRYB[9][21] ), .CI(\mult_19/SUMB[9][22] ), .CO(
        \mult_19/CARRYB[10][21] ), .S(\mult_19/SUMB[10][21] ) );
  FA_X1 \mult_19/S2_10_20  ( .A(\mult_19/ab[10][20] ), .B(
        \mult_19/CARRYB[9][20] ), .CI(\mult_19/SUMB[9][21] ), .CO(
        \mult_19/CARRYB[10][20] ), .S(\mult_19/SUMB[10][20] ) );
  FA_X1 \mult_19/S2_10_19  ( .A(\mult_19/ab[10][19] ), .B(
        \mult_19/CARRYB[9][19] ), .CI(\mult_19/SUMB[9][20] ), .CO(
        \mult_19/CARRYB[10][19] ), .S(\mult_19/SUMB[10][19] ) );
  FA_X1 \mult_19/S2_10_18  ( .A(\mult_19/ab[10][18] ), .B(
        \mult_19/CARRYB[9][18] ), .CI(\mult_19/SUMB[9][19] ), .CO(
        \mult_19/CARRYB[10][18] ), .S(\mult_19/SUMB[10][18] ) );
  FA_X1 \mult_19/S2_10_17  ( .A(\mult_19/ab[10][17] ), .B(
        \mult_19/CARRYB[9][17] ), .CI(\mult_19/SUMB[9][18] ), .CO(
        \mult_19/CARRYB[10][17] ), .S(\mult_19/SUMB[10][17] ) );
  FA_X1 \mult_19/S2_10_16  ( .A(\mult_19/ab[10][16] ), .B(
        \mult_19/CARRYB[9][16] ), .CI(\mult_19/SUMB[9][17] ), .CO(
        \mult_19/CARRYB[10][16] ), .S(\mult_19/SUMB[10][16] ) );
  FA_X1 \mult_19/S2_10_15  ( .A(\mult_19/ab[10][15] ), .B(
        \mult_19/CARRYB[9][15] ), .CI(\mult_19/SUMB[9][16] ), .CO(
        \mult_19/CARRYB[10][15] ), .S(\mult_19/SUMB[10][15] ) );
  FA_X1 \mult_19/S2_10_14  ( .A(\mult_19/ab[10][14] ), .B(
        \mult_19/CARRYB[9][14] ), .CI(\mult_19/SUMB[9][15] ), .CO(
        \mult_19/CARRYB[10][14] ), .S(\mult_19/SUMB[10][14] ) );
  FA_X1 \mult_19/S2_10_13  ( .A(\mult_19/ab[10][13] ), .B(
        \mult_19/CARRYB[9][13] ), .CI(\mult_19/SUMB[9][14] ), .CO(
        \mult_19/CARRYB[10][13] ), .S(\mult_19/SUMB[10][13] ) );
  FA_X1 \mult_19/S2_10_12  ( .A(\mult_19/ab[10][12] ), .B(
        \mult_19/CARRYB[9][12] ), .CI(\mult_19/SUMB[9][13] ), .CO(
        \mult_19/CARRYB[10][12] ), .S(\mult_19/SUMB[10][12] ) );
  FA_X1 \mult_19/S2_10_11  ( .A(\mult_19/ab[10][11] ), .B(
        \mult_19/CARRYB[9][11] ), .CI(\mult_19/SUMB[9][12] ), .CO(
        \mult_19/CARRYB[10][11] ), .S(\mult_19/SUMB[10][11] ) );
  FA_X1 \mult_19/S2_10_10  ( .A(\mult_19/ab[10][10] ), .B(
        \mult_19/CARRYB[9][10] ), .CI(\mult_19/SUMB[9][11] ), .CO(
        \mult_19/CARRYB[10][10] ), .S(\mult_19/SUMB[10][10] ) );
  FA_X1 \mult_19/S2_10_9  ( .A(\mult_19/ab[10][9] ), .B(\mult_19/CARRYB[9][9] ), .CI(\mult_19/SUMB[9][10] ), .CO(\mult_19/CARRYB[10][9] ), .S(
        \mult_19/SUMB[10][9] ) );
  FA_X1 \mult_19/S2_10_8  ( .A(\mult_19/ab[10][8] ), .B(\mult_19/CARRYB[9][8] ), .CI(\mult_19/SUMB[9][9] ), .CO(\mult_19/CARRYB[10][8] ), .S(
        \mult_19/SUMB[10][8] ) );
  FA_X1 \mult_19/S2_10_7  ( .A(\mult_19/ab[10][7] ), .B(\mult_19/CARRYB[9][7] ), .CI(\mult_19/SUMB[9][8] ), .CO(\mult_19/CARRYB[10][7] ), .S(
        \mult_19/SUMB[10][7] ) );
  FA_X1 \mult_19/S2_10_6  ( .A(\mult_19/ab[10][6] ), .B(\mult_19/CARRYB[9][6] ), .CI(\mult_19/SUMB[9][7] ), .CO(\mult_19/CARRYB[10][6] ), .S(
        \mult_19/SUMB[10][6] ) );
  FA_X1 \mult_19/S2_10_5  ( .A(\mult_19/ab[10][5] ), .B(\mult_19/CARRYB[9][5] ), .CI(\mult_19/SUMB[9][6] ), .CO(\mult_19/CARRYB[10][5] ), .S(
        \mult_19/SUMB[10][5] ) );
  FA_X1 \mult_19/S2_10_4  ( .A(\mult_19/ab[10][4] ), .B(\mult_19/CARRYB[9][4] ), .CI(\mult_19/SUMB[9][5] ), .CO(\mult_19/CARRYB[10][4] ), .S(
        \mult_19/SUMB[10][4] ) );
  FA_X1 \mult_19/S2_10_3  ( .A(\mult_19/ab[10][3] ), .B(\mult_19/CARRYB[9][3] ), .CI(\mult_19/SUMB[9][4] ), .CO(\mult_19/CARRYB[10][3] ), .S(
        \mult_19/SUMB[10][3] ) );
  FA_X1 \mult_19/S2_10_2  ( .A(\mult_19/ab[10][2] ), .B(\mult_19/CARRYB[9][2] ), .CI(\mult_19/SUMB[9][3] ), .CO(\mult_19/CARRYB[10][2] ), .S(
        \mult_19/SUMB[10][2] ) );
  FA_X1 \mult_19/S2_10_1  ( .A(\mult_19/ab[10][1] ), .B(\mult_19/CARRYB[9][1] ), .CI(\mult_19/SUMB[9][2] ), .CO(\mult_19/CARRYB[10][1] ), .S(
        \mult_19/SUMB[10][1] ) );
  FA_X1 \mult_19/S1_10_0  ( .A(\mult_19/ab[10][0] ), .B(\mult_19/CARRYB[9][0] ), .CI(\mult_19/SUMB[9][1] ), .CO(\mult_19/CARRYB[10][0] ), .S(N10) );
  FA_X1 \mult_19/S3_11_30  ( .A(\mult_19/ab[11][30] ), .B(
        \mult_19/CARRYB[10][30] ), .CI(\mult_19/ab[10][31] ), .CO(
        \mult_19/CARRYB[11][30] ), .S(\mult_19/SUMB[11][30] ) );
  FA_X1 \mult_19/S2_11_29  ( .A(\mult_19/ab[11][29] ), .B(
        \mult_19/CARRYB[10][29] ), .CI(\mult_19/SUMB[10][30] ), .CO(
        \mult_19/CARRYB[11][29] ), .S(\mult_19/SUMB[11][29] ) );
  FA_X1 \mult_19/S2_11_28  ( .A(\mult_19/ab[11][28] ), .B(
        \mult_19/CARRYB[10][28] ), .CI(\mult_19/SUMB[10][29] ), .CO(
        \mult_19/CARRYB[11][28] ), .S(\mult_19/SUMB[11][28] ) );
  FA_X1 \mult_19/S2_11_27  ( .A(\mult_19/ab[11][27] ), .B(
        \mult_19/CARRYB[10][27] ), .CI(\mult_19/SUMB[10][28] ), .CO(
        \mult_19/CARRYB[11][27] ), .S(\mult_19/SUMB[11][27] ) );
  FA_X1 \mult_19/S2_11_26  ( .A(\mult_19/ab[11][26] ), .B(
        \mult_19/CARRYB[10][26] ), .CI(\mult_19/SUMB[10][27] ), .CO(
        \mult_19/CARRYB[11][26] ), .S(\mult_19/SUMB[11][26] ) );
  FA_X1 \mult_19/S2_11_25  ( .A(\mult_19/ab[11][25] ), .B(
        \mult_19/CARRYB[10][25] ), .CI(\mult_19/SUMB[10][26] ), .CO(
        \mult_19/CARRYB[11][25] ), .S(\mult_19/SUMB[11][25] ) );
  FA_X1 \mult_19/S2_11_24  ( .A(\mult_19/ab[11][24] ), .B(
        \mult_19/CARRYB[10][24] ), .CI(\mult_19/SUMB[10][25] ), .CO(
        \mult_19/CARRYB[11][24] ), .S(\mult_19/SUMB[11][24] ) );
  FA_X1 \mult_19/S2_11_23  ( .A(\mult_19/ab[11][23] ), .B(
        \mult_19/CARRYB[10][23] ), .CI(\mult_19/SUMB[10][24] ), .CO(
        \mult_19/CARRYB[11][23] ), .S(\mult_19/SUMB[11][23] ) );
  FA_X1 \mult_19/S2_11_22  ( .A(\mult_19/ab[11][22] ), .B(
        \mult_19/CARRYB[10][22] ), .CI(\mult_19/SUMB[10][23] ), .CO(
        \mult_19/CARRYB[11][22] ), .S(\mult_19/SUMB[11][22] ) );
  FA_X1 \mult_19/S2_11_21  ( .A(\mult_19/ab[11][21] ), .B(
        \mult_19/CARRYB[10][21] ), .CI(\mult_19/SUMB[10][22] ), .CO(
        \mult_19/CARRYB[11][21] ), .S(\mult_19/SUMB[11][21] ) );
  FA_X1 \mult_19/S2_11_20  ( .A(\mult_19/ab[11][20] ), .B(
        \mult_19/CARRYB[10][20] ), .CI(\mult_19/SUMB[10][21] ), .CO(
        \mult_19/CARRYB[11][20] ), .S(\mult_19/SUMB[11][20] ) );
  FA_X1 \mult_19/S2_11_19  ( .A(\mult_19/ab[11][19] ), .B(
        \mult_19/CARRYB[10][19] ), .CI(\mult_19/SUMB[10][20] ), .CO(
        \mult_19/CARRYB[11][19] ), .S(\mult_19/SUMB[11][19] ) );
  FA_X1 \mult_19/S2_11_18  ( .A(\mult_19/ab[11][18] ), .B(
        \mult_19/CARRYB[10][18] ), .CI(\mult_19/SUMB[10][19] ), .CO(
        \mult_19/CARRYB[11][18] ), .S(\mult_19/SUMB[11][18] ) );
  FA_X1 \mult_19/S2_11_17  ( .A(\mult_19/ab[11][17] ), .B(
        \mult_19/CARRYB[10][17] ), .CI(\mult_19/SUMB[10][18] ), .CO(
        \mult_19/CARRYB[11][17] ), .S(\mult_19/SUMB[11][17] ) );
  FA_X1 \mult_19/S2_11_16  ( .A(\mult_19/ab[11][16] ), .B(
        \mult_19/CARRYB[10][16] ), .CI(\mult_19/SUMB[10][17] ), .CO(
        \mult_19/CARRYB[11][16] ), .S(\mult_19/SUMB[11][16] ) );
  FA_X1 \mult_19/S2_11_15  ( .A(\mult_19/ab[11][15] ), .B(
        \mult_19/CARRYB[10][15] ), .CI(\mult_19/SUMB[10][16] ), .CO(
        \mult_19/CARRYB[11][15] ), .S(\mult_19/SUMB[11][15] ) );
  FA_X1 \mult_19/S2_11_14  ( .A(\mult_19/ab[11][14] ), .B(
        \mult_19/CARRYB[10][14] ), .CI(\mult_19/SUMB[10][15] ), .CO(
        \mult_19/CARRYB[11][14] ), .S(\mult_19/SUMB[11][14] ) );
  FA_X1 \mult_19/S2_11_13  ( .A(\mult_19/ab[11][13] ), .B(
        \mult_19/CARRYB[10][13] ), .CI(\mult_19/SUMB[10][14] ), .CO(
        \mult_19/CARRYB[11][13] ), .S(\mult_19/SUMB[11][13] ) );
  FA_X1 \mult_19/S2_11_12  ( .A(\mult_19/ab[11][12] ), .B(
        \mult_19/CARRYB[10][12] ), .CI(\mult_19/SUMB[10][13] ), .CO(
        \mult_19/CARRYB[11][12] ), .S(\mult_19/SUMB[11][12] ) );
  FA_X1 \mult_19/S2_11_11  ( .A(\mult_19/ab[11][11] ), .B(
        \mult_19/CARRYB[10][11] ), .CI(\mult_19/SUMB[10][12] ), .CO(
        \mult_19/CARRYB[11][11] ), .S(\mult_19/SUMB[11][11] ) );
  FA_X1 \mult_19/S2_11_10  ( .A(\mult_19/ab[11][10] ), .B(
        \mult_19/CARRYB[10][10] ), .CI(\mult_19/SUMB[10][11] ), .CO(
        \mult_19/CARRYB[11][10] ), .S(\mult_19/SUMB[11][10] ) );
  FA_X1 \mult_19/S2_11_9  ( .A(\mult_19/ab[11][9] ), .B(
        \mult_19/CARRYB[10][9] ), .CI(\mult_19/SUMB[10][10] ), .CO(
        \mult_19/CARRYB[11][9] ), .S(\mult_19/SUMB[11][9] ) );
  FA_X1 \mult_19/S2_11_8  ( .A(\mult_19/ab[11][8] ), .B(
        \mult_19/CARRYB[10][8] ), .CI(\mult_19/SUMB[10][9] ), .CO(
        \mult_19/CARRYB[11][8] ), .S(\mult_19/SUMB[11][8] ) );
  FA_X1 \mult_19/S2_11_7  ( .A(\mult_19/ab[11][7] ), .B(
        \mult_19/CARRYB[10][7] ), .CI(\mult_19/SUMB[10][8] ), .CO(
        \mult_19/CARRYB[11][7] ), .S(\mult_19/SUMB[11][7] ) );
  FA_X1 \mult_19/S2_11_6  ( .A(\mult_19/ab[11][6] ), .B(
        \mult_19/CARRYB[10][6] ), .CI(\mult_19/SUMB[10][7] ), .CO(
        \mult_19/CARRYB[11][6] ), .S(\mult_19/SUMB[11][6] ) );
  FA_X1 \mult_19/S2_11_5  ( .A(\mult_19/ab[11][5] ), .B(
        \mult_19/CARRYB[10][5] ), .CI(\mult_19/SUMB[10][6] ), .CO(
        \mult_19/CARRYB[11][5] ), .S(\mult_19/SUMB[11][5] ) );
  FA_X1 \mult_19/S2_11_4  ( .A(\mult_19/ab[11][4] ), .B(
        \mult_19/CARRYB[10][4] ), .CI(\mult_19/SUMB[10][5] ), .CO(
        \mult_19/CARRYB[11][4] ), .S(\mult_19/SUMB[11][4] ) );
  FA_X1 \mult_19/S2_11_3  ( .A(\mult_19/ab[11][3] ), .B(
        \mult_19/CARRYB[10][3] ), .CI(\mult_19/SUMB[10][4] ), .CO(
        \mult_19/CARRYB[11][3] ), .S(\mult_19/SUMB[11][3] ) );
  FA_X1 \mult_19/S2_11_2  ( .A(\mult_19/ab[11][2] ), .B(
        \mult_19/CARRYB[10][2] ), .CI(\mult_19/SUMB[10][3] ), .CO(
        \mult_19/CARRYB[11][2] ), .S(\mult_19/SUMB[11][2] ) );
  FA_X1 \mult_19/S2_11_1  ( .A(\mult_19/ab[11][1] ), .B(
        \mult_19/CARRYB[10][1] ), .CI(\mult_19/SUMB[10][2] ), .CO(
        \mult_19/CARRYB[11][1] ), .S(\mult_19/SUMB[11][1] ) );
  FA_X1 \mult_19/S1_11_0  ( .A(\mult_19/ab[11][0] ), .B(
        \mult_19/CARRYB[10][0] ), .CI(\mult_19/SUMB[10][1] ), .CO(
        \mult_19/CARRYB[11][0] ), .S(N11) );
  FA_X1 \mult_19/S3_12_30  ( .A(\mult_19/ab[12][30] ), .B(
        \mult_19/CARRYB[11][30] ), .CI(\mult_19/ab[11][31] ), .CO(
        \mult_19/CARRYB[12][30] ), .S(\mult_19/SUMB[12][30] ) );
  FA_X1 \mult_19/S2_12_29  ( .A(\mult_19/ab[12][29] ), .B(
        \mult_19/CARRYB[11][29] ), .CI(\mult_19/SUMB[11][30] ), .CO(
        \mult_19/CARRYB[12][29] ), .S(\mult_19/SUMB[12][29] ) );
  FA_X1 \mult_19/S2_12_28  ( .A(\mult_19/ab[12][28] ), .B(
        \mult_19/CARRYB[11][28] ), .CI(\mult_19/SUMB[11][29] ), .CO(
        \mult_19/CARRYB[12][28] ), .S(\mult_19/SUMB[12][28] ) );
  FA_X1 \mult_19/S2_12_27  ( .A(\mult_19/ab[12][27] ), .B(
        \mult_19/CARRYB[11][27] ), .CI(\mult_19/SUMB[11][28] ), .CO(
        \mult_19/CARRYB[12][27] ), .S(\mult_19/SUMB[12][27] ) );
  FA_X1 \mult_19/S2_12_26  ( .A(\mult_19/ab[12][26] ), .B(
        \mult_19/CARRYB[11][26] ), .CI(\mult_19/SUMB[11][27] ), .CO(
        \mult_19/CARRYB[12][26] ), .S(\mult_19/SUMB[12][26] ) );
  FA_X1 \mult_19/S2_12_25  ( .A(\mult_19/ab[12][25] ), .B(
        \mult_19/CARRYB[11][25] ), .CI(\mult_19/SUMB[11][26] ), .CO(
        \mult_19/CARRYB[12][25] ), .S(\mult_19/SUMB[12][25] ) );
  FA_X1 \mult_19/S2_12_24  ( .A(\mult_19/ab[12][24] ), .B(
        \mult_19/CARRYB[11][24] ), .CI(\mult_19/SUMB[11][25] ), .CO(
        \mult_19/CARRYB[12][24] ), .S(\mult_19/SUMB[12][24] ) );
  FA_X1 \mult_19/S2_12_23  ( .A(\mult_19/ab[12][23] ), .B(
        \mult_19/CARRYB[11][23] ), .CI(\mult_19/SUMB[11][24] ), .CO(
        \mult_19/CARRYB[12][23] ), .S(\mult_19/SUMB[12][23] ) );
  FA_X1 \mult_19/S2_12_22  ( .A(\mult_19/ab[12][22] ), .B(
        \mult_19/CARRYB[11][22] ), .CI(\mult_19/SUMB[11][23] ), .CO(
        \mult_19/CARRYB[12][22] ), .S(\mult_19/SUMB[12][22] ) );
  FA_X1 \mult_19/S2_12_21  ( .A(\mult_19/ab[12][21] ), .B(
        \mult_19/CARRYB[11][21] ), .CI(\mult_19/SUMB[11][22] ), .CO(
        \mult_19/CARRYB[12][21] ), .S(\mult_19/SUMB[12][21] ) );
  FA_X1 \mult_19/S2_12_20  ( .A(\mult_19/ab[12][20] ), .B(
        \mult_19/CARRYB[11][20] ), .CI(\mult_19/SUMB[11][21] ), .CO(
        \mult_19/CARRYB[12][20] ), .S(\mult_19/SUMB[12][20] ) );
  FA_X1 \mult_19/S2_12_19  ( .A(\mult_19/ab[12][19] ), .B(
        \mult_19/CARRYB[11][19] ), .CI(\mult_19/SUMB[11][20] ), .CO(
        \mult_19/CARRYB[12][19] ), .S(\mult_19/SUMB[12][19] ) );
  FA_X1 \mult_19/S2_12_18  ( .A(\mult_19/ab[12][18] ), .B(
        \mult_19/CARRYB[11][18] ), .CI(\mult_19/SUMB[11][19] ), .CO(
        \mult_19/CARRYB[12][18] ), .S(\mult_19/SUMB[12][18] ) );
  FA_X1 \mult_19/S2_12_17  ( .A(\mult_19/ab[12][17] ), .B(
        \mult_19/CARRYB[11][17] ), .CI(\mult_19/SUMB[11][18] ), .CO(
        \mult_19/CARRYB[12][17] ), .S(\mult_19/SUMB[12][17] ) );
  FA_X1 \mult_19/S2_12_16  ( .A(\mult_19/ab[12][16] ), .B(
        \mult_19/CARRYB[11][16] ), .CI(\mult_19/SUMB[11][17] ), .CO(
        \mult_19/CARRYB[12][16] ), .S(\mult_19/SUMB[12][16] ) );
  FA_X1 \mult_19/S2_12_15  ( .A(\mult_19/ab[12][15] ), .B(
        \mult_19/CARRYB[11][15] ), .CI(\mult_19/SUMB[11][16] ), .CO(
        \mult_19/CARRYB[12][15] ), .S(\mult_19/SUMB[12][15] ) );
  FA_X1 \mult_19/S2_12_14  ( .A(\mult_19/ab[12][14] ), .B(
        \mult_19/CARRYB[11][14] ), .CI(\mult_19/SUMB[11][15] ), .CO(
        \mult_19/CARRYB[12][14] ), .S(\mult_19/SUMB[12][14] ) );
  FA_X1 \mult_19/S2_12_13  ( .A(\mult_19/ab[12][13] ), .B(
        \mult_19/CARRYB[11][13] ), .CI(\mult_19/SUMB[11][14] ), .CO(
        \mult_19/CARRYB[12][13] ), .S(\mult_19/SUMB[12][13] ) );
  FA_X1 \mult_19/S2_12_12  ( .A(\mult_19/ab[12][12] ), .B(
        \mult_19/CARRYB[11][12] ), .CI(\mult_19/SUMB[11][13] ), .CO(
        \mult_19/CARRYB[12][12] ), .S(\mult_19/SUMB[12][12] ) );
  FA_X1 \mult_19/S2_12_11  ( .A(\mult_19/ab[12][11] ), .B(
        \mult_19/CARRYB[11][11] ), .CI(\mult_19/SUMB[11][12] ), .CO(
        \mult_19/CARRYB[12][11] ), .S(\mult_19/SUMB[12][11] ) );
  FA_X1 \mult_19/S2_12_10  ( .A(\mult_19/ab[12][10] ), .B(
        \mult_19/CARRYB[11][10] ), .CI(\mult_19/SUMB[11][11] ), .CO(
        \mult_19/CARRYB[12][10] ), .S(\mult_19/SUMB[12][10] ) );
  FA_X1 \mult_19/S2_12_9  ( .A(\mult_19/ab[12][9] ), .B(
        \mult_19/CARRYB[11][9] ), .CI(\mult_19/SUMB[11][10] ), .CO(
        \mult_19/CARRYB[12][9] ), .S(\mult_19/SUMB[12][9] ) );
  FA_X1 \mult_19/S2_12_8  ( .A(\mult_19/ab[12][8] ), .B(
        \mult_19/CARRYB[11][8] ), .CI(\mult_19/SUMB[11][9] ), .CO(
        \mult_19/CARRYB[12][8] ), .S(\mult_19/SUMB[12][8] ) );
  FA_X1 \mult_19/S2_12_7  ( .A(\mult_19/ab[12][7] ), .B(
        \mult_19/CARRYB[11][7] ), .CI(\mult_19/SUMB[11][8] ), .CO(
        \mult_19/CARRYB[12][7] ), .S(\mult_19/SUMB[12][7] ) );
  FA_X1 \mult_19/S2_12_6  ( .A(\mult_19/ab[12][6] ), .B(
        \mult_19/CARRYB[11][6] ), .CI(\mult_19/SUMB[11][7] ), .CO(
        \mult_19/CARRYB[12][6] ), .S(\mult_19/SUMB[12][6] ) );
  FA_X1 \mult_19/S2_12_5  ( .A(\mult_19/ab[12][5] ), .B(
        \mult_19/CARRYB[11][5] ), .CI(\mult_19/SUMB[11][6] ), .CO(
        \mult_19/CARRYB[12][5] ), .S(\mult_19/SUMB[12][5] ) );
  FA_X1 \mult_19/S2_12_4  ( .A(\mult_19/ab[12][4] ), .B(
        \mult_19/CARRYB[11][4] ), .CI(\mult_19/SUMB[11][5] ), .CO(
        \mult_19/CARRYB[12][4] ), .S(\mult_19/SUMB[12][4] ) );
  FA_X1 \mult_19/S2_12_3  ( .A(\mult_19/ab[12][3] ), .B(
        \mult_19/CARRYB[11][3] ), .CI(\mult_19/SUMB[11][4] ), .CO(
        \mult_19/CARRYB[12][3] ), .S(\mult_19/SUMB[12][3] ) );
  FA_X1 \mult_19/S2_12_2  ( .A(\mult_19/ab[12][2] ), .B(
        \mult_19/CARRYB[11][2] ), .CI(\mult_19/SUMB[11][3] ), .CO(
        \mult_19/CARRYB[12][2] ), .S(\mult_19/SUMB[12][2] ) );
  FA_X1 \mult_19/S2_12_1  ( .A(\mult_19/ab[12][1] ), .B(
        \mult_19/CARRYB[11][1] ), .CI(\mult_19/SUMB[11][2] ), .CO(
        \mult_19/CARRYB[12][1] ), .S(\mult_19/SUMB[12][1] ) );
  FA_X1 \mult_19/S1_12_0  ( .A(\mult_19/ab[12][0] ), .B(
        \mult_19/CARRYB[11][0] ), .CI(\mult_19/SUMB[11][1] ), .CO(
        \mult_19/CARRYB[12][0] ), .S(N12) );
  FA_X1 \mult_19/S3_13_30  ( .A(\mult_19/ab[13][30] ), .B(
        \mult_19/CARRYB[12][30] ), .CI(\mult_19/ab[12][31] ), .CO(
        \mult_19/CARRYB[13][30] ), .S(\mult_19/SUMB[13][30] ) );
  FA_X1 \mult_19/S2_13_29  ( .A(\mult_19/ab[13][29] ), .B(
        \mult_19/CARRYB[12][29] ), .CI(\mult_19/SUMB[12][30] ), .CO(
        \mult_19/CARRYB[13][29] ), .S(\mult_19/SUMB[13][29] ) );
  FA_X1 \mult_19/S2_13_28  ( .A(\mult_19/ab[13][28] ), .B(
        \mult_19/CARRYB[12][28] ), .CI(\mult_19/SUMB[12][29] ), .CO(
        \mult_19/CARRYB[13][28] ), .S(\mult_19/SUMB[13][28] ) );
  FA_X1 \mult_19/S2_13_27  ( .A(\mult_19/ab[13][27] ), .B(
        \mult_19/CARRYB[12][27] ), .CI(\mult_19/SUMB[12][28] ), .CO(
        \mult_19/CARRYB[13][27] ), .S(\mult_19/SUMB[13][27] ) );
  FA_X1 \mult_19/S2_13_26  ( .A(\mult_19/ab[13][26] ), .B(
        \mult_19/CARRYB[12][26] ), .CI(\mult_19/SUMB[12][27] ), .CO(
        \mult_19/CARRYB[13][26] ), .S(\mult_19/SUMB[13][26] ) );
  FA_X1 \mult_19/S2_13_25  ( .A(\mult_19/ab[13][25] ), .B(
        \mult_19/CARRYB[12][25] ), .CI(\mult_19/SUMB[12][26] ), .CO(
        \mult_19/CARRYB[13][25] ), .S(\mult_19/SUMB[13][25] ) );
  FA_X1 \mult_19/S2_13_24  ( .A(\mult_19/ab[13][24] ), .B(
        \mult_19/CARRYB[12][24] ), .CI(\mult_19/SUMB[12][25] ), .CO(
        \mult_19/CARRYB[13][24] ), .S(\mult_19/SUMB[13][24] ) );
  FA_X1 \mult_19/S2_13_23  ( .A(\mult_19/ab[13][23] ), .B(
        \mult_19/CARRYB[12][23] ), .CI(\mult_19/SUMB[12][24] ), .CO(
        \mult_19/CARRYB[13][23] ), .S(\mult_19/SUMB[13][23] ) );
  FA_X1 \mult_19/S2_13_22  ( .A(\mult_19/ab[13][22] ), .B(
        \mult_19/CARRYB[12][22] ), .CI(\mult_19/SUMB[12][23] ), .CO(
        \mult_19/CARRYB[13][22] ), .S(\mult_19/SUMB[13][22] ) );
  FA_X1 \mult_19/S2_13_21  ( .A(\mult_19/ab[13][21] ), .B(
        \mult_19/CARRYB[12][21] ), .CI(\mult_19/SUMB[12][22] ), .CO(
        \mult_19/CARRYB[13][21] ), .S(\mult_19/SUMB[13][21] ) );
  FA_X1 \mult_19/S2_13_20  ( .A(\mult_19/ab[13][20] ), .B(
        \mult_19/CARRYB[12][20] ), .CI(\mult_19/SUMB[12][21] ), .CO(
        \mult_19/CARRYB[13][20] ), .S(\mult_19/SUMB[13][20] ) );
  FA_X1 \mult_19/S2_13_19  ( .A(\mult_19/ab[13][19] ), .B(
        \mult_19/CARRYB[12][19] ), .CI(\mult_19/SUMB[12][20] ), .CO(
        \mult_19/CARRYB[13][19] ), .S(\mult_19/SUMB[13][19] ) );
  FA_X1 \mult_19/S2_13_18  ( .A(\mult_19/ab[13][18] ), .B(
        \mult_19/CARRYB[12][18] ), .CI(\mult_19/SUMB[12][19] ), .CO(
        \mult_19/CARRYB[13][18] ), .S(\mult_19/SUMB[13][18] ) );
  FA_X1 \mult_19/S2_13_17  ( .A(\mult_19/ab[13][17] ), .B(
        \mult_19/CARRYB[12][17] ), .CI(\mult_19/SUMB[12][18] ), .CO(
        \mult_19/CARRYB[13][17] ), .S(\mult_19/SUMB[13][17] ) );
  FA_X1 \mult_19/S2_13_16  ( .A(\mult_19/ab[13][16] ), .B(
        \mult_19/CARRYB[12][16] ), .CI(\mult_19/SUMB[12][17] ), .CO(
        \mult_19/CARRYB[13][16] ), .S(\mult_19/SUMB[13][16] ) );
  FA_X1 \mult_19/S2_13_15  ( .A(\mult_19/ab[13][15] ), .B(
        \mult_19/CARRYB[12][15] ), .CI(\mult_19/SUMB[12][16] ), .CO(
        \mult_19/CARRYB[13][15] ), .S(\mult_19/SUMB[13][15] ) );
  FA_X1 \mult_19/S2_13_14  ( .A(\mult_19/ab[13][14] ), .B(
        \mult_19/CARRYB[12][14] ), .CI(\mult_19/SUMB[12][15] ), .CO(
        \mult_19/CARRYB[13][14] ), .S(\mult_19/SUMB[13][14] ) );
  FA_X1 \mult_19/S2_13_13  ( .A(\mult_19/ab[13][13] ), .B(
        \mult_19/CARRYB[12][13] ), .CI(\mult_19/SUMB[12][14] ), .CO(
        \mult_19/CARRYB[13][13] ), .S(\mult_19/SUMB[13][13] ) );
  FA_X1 \mult_19/S2_13_12  ( .A(\mult_19/ab[13][12] ), .B(
        \mult_19/CARRYB[12][12] ), .CI(\mult_19/SUMB[12][13] ), .CO(
        \mult_19/CARRYB[13][12] ), .S(\mult_19/SUMB[13][12] ) );
  FA_X1 \mult_19/S2_13_11  ( .A(\mult_19/ab[13][11] ), .B(
        \mult_19/CARRYB[12][11] ), .CI(\mult_19/SUMB[12][12] ), .CO(
        \mult_19/CARRYB[13][11] ), .S(\mult_19/SUMB[13][11] ) );
  FA_X1 \mult_19/S2_13_10  ( .A(\mult_19/ab[13][10] ), .B(
        \mult_19/CARRYB[12][10] ), .CI(\mult_19/SUMB[12][11] ), .CO(
        \mult_19/CARRYB[13][10] ), .S(\mult_19/SUMB[13][10] ) );
  FA_X1 \mult_19/S2_13_9  ( .A(\mult_19/ab[13][9] ), .B(
        \mult_19/CARRYB[12][9] ), .CI(\mult_19/SUMB[12][10] ), .CO(
        \mult_19/CARRYB[13][9] ), .S(\mult_19/SUMB[13][9] ) );
  FA_X1 \mult_19/S2_13_8  ( .A(\mult_19/ab[13][8] ), .B(
        \mult_19/CARRYB[12][8] ), .CI(\mult_19/SUMB[12][9] ), .CO(
        \mult_19/CARRYB[13][8] ), .S(\mult_19/SUMB[13][8] ) );
  FA_X1 \mult_19/S2_13_7  ( .A(\mult_19/ab[13][7] ), .B(
        \mult_19/CARRYB[12][7] ), .CI(\mult_19/SUMB[12][8] ), .CO(
        \mult_19/CARRYB[13][7] ), .S(\mult_19/SUMB[13][7] ) );
  FA_X1 \mult_19/S2_13_6  ( .A(\mult_19/ab[13][6] ), .B(
        \mult_19/CARRYB[12][6] ), .CI(\mult_19/SUMB[12][7] ), .CO(
        \mult_19/CARRYB[13][6] ), .S(\mult_19/SUMB[13][6] ) );
  FA_X1 \mult_19/S2_13_5  ( .A(\mult_19/ab[13][5] ), .B(
        \mult_19/CARRYB[12][5] ), .CI(\mult_19/SUMB[12][6] ), .CO(
        \mult_19/CARRYB[13][5] ), .S(\mult_19/SUMB[13][5] ) );
  FA_X1 \mult_19/S2_13_4  ( .A(\mult_19/ab[13][4] ), .B(
        \mult_19/CARRYB[12][4] ), .CI(\mult_19/SUMB[12][5] ), .CO(
        \mult_19/CARRYB[13][4] ), .S(\mult_19/SUMB[13][4] ) );
  FA_X1 \mult_19/S2_13_3  ( .A(\mult_19/ab[13][3] ), .B(
        \mult_19/CARRYB[12][3] ), .CI(\mult_19/SUMB[12][4] ), .CO(
        \mult_19/CARRYB[13][3] ), .S(\mult_19/SUMB[13][3] ) );
  FA_X1 \mult_19/S2_13_2  ( .A(\mult_19/ab[13][2] ), .B(
        \mult_19/CARRYB[12][2] ), .CI(\mult_19/SUMB[12][3] ), .CO(
        \mult_19/CARRYB[13][2] ), .S(\mult_19/SUMB[13][2] ) );
  FA_X1 \mult_19/S2_13_1  ( .A(\mult_19/ab[13][1] ), .B(
        \mult_19/CARRYB[12][1] ), .CI(\mult_19/SUMB[12][2] ), .CO(
        \mult_19/CARRYB[13][1] ), .S(\mult_19/SUMB[13][1] ) );
  FA_X1 \mult_19/S1_13_0  ( .A(\mult_19/ab[13][0] ), .B(
        \mult_19/CARRYB[12][0] ), .CI(\mult_19/SUMB[12][1] ), .CO(
        \mult_19/CARRYB[13][0] ), .S(N13) );
  FA_X1 \mult_19/S3_14_30  ( .A(\mult_19/ab[14][30] ), .B(
        \mult_19/CARRYB[13][30] ), .CI(\mult_19/ab[13][31] ), .CO(
        \mult_19/CARRYB[14][30] ), .S(\mult_19/SUMB[14][30] ) );
  FA_X1 \mult_19/S2_14_29  ( .A(\mult_19/ab[14][29] ), .B(
        \mult_19/CARRYB[13][29] ), .CI(\mult_19/SUMB[13][30] ), .CO(
        \mult_19/CARRYB[14][29] ), .S(\mult_19/SUMB[14][29] ) );
  FA_X1 \mult_19/S2_14_28  ( .A(\mult_19/ab[14][28] ), .B(
        \mult_19/CARRYB[13][28] ), .CI(\mult_19/SUMB[13][29] ), .CO(
        \mult_19/CARRYB[14][28] ), .S(\mult_19/SUMB[14][28] ) );
  FA_X1 \mult_19/S2_14_27  ( .A(\mult_19/ab[14][27] ), .B(
        \mult_19/CARRYB[13][27] ), .CI(\mult_19/SUMB[13][28] ), .CO(
        \mult_19/CARRYB[14][27] ), .S(\mult_19/SUMB[14][27] ) );
  FA_X1 \mult_19/S2_14_26  ( .A(\mult_19/ab[14][26] ), .B(
        \mult_19/CARRYB[13][26] ), .CI(\mult_19/SUMB[13][27] ), .CO(
        \mult_19/CARRYB[14][26] ), .S(\mult_19/SUMB[14][26] ) );
  FA_X1 \mult_19/S2_14_25  ( .A(\mult_19/ab[14][25] ), .B(
        \mult_19/CARRYB[13][25] ), .CI(\mult_19/SUMB[13][26] ), .CO(
        \mult_19/CARRYB[14][25] ), .S(\mult_19/SUMB[14][25] ) );
  FA_X1 \mult_19/S2_14_24  ( .A(\mult_19/ab[14][24] ), .B(
        \mult_19/CARRYB[13][24] ), .CI(\mult_19/SUMB[13][25] ), .CO(
        \mult_19/CARRYB[14][24] ), .S(\mult_19/SUMB[14][24] ) );
  FA_X1 \mult_19/S2_14_23  ( .A(\mult_19/ab[14][23] ), .B(
        \mult_19/CARRYB[13][23] ), .CI(\mult_19/SUMB[13][24] ), .CO(
        \mult_19/CARRYB[14][23] ), .S(\mult_19/SUMB[14][23] ) );
  FA_X1 \mult_19/S2_14_22  ( .A(\mult_19/ab[14][22] ), .B(
        \mult_19/CARRYB[13][22] ), .CI(\mult_19/SUMB[13][23] ), .CO(
        \mult_19/CARRYB[14][22] ), .S(\mult_19/SUMB[14][22] ) );
  FA_X1 \mult_19/S2_14_21  ( .A(\mult_19/ab[14][21] ), .B(
        \mult_19/CARRYB[13][21] ), .CI(\mult_19/SUMB[13][22] ), .CO(
        \mult_19/CARRYB[14][21] ), .S(\mult_19/SUMB[14][21] ) );
  FA_X1 \mult_19/S2_14_20  ( .A(\mult_19/ab[14][20] ), .B(
        \mult_19/CARRYB[13][20] ), .CI(\mult_19/SUMB[13][21] ), .CO(
        \mult_19/CARRYB[14][20] ), .S(\mult_19/SUMB[14][20] ) );
  FA_X1 \mult_19/S2_14_19  ( .A(\mult_19/ab[14][19] ), .B(
        \mult_19/CARRYB[13][19] ), .CI(\mult_19/SUMB[13][20] ), .CO(
        \mult_19/CARRYB[14][19] ), .S(\mult_19/SUMB[14][19] ) );
  FA_X1 \mult_19/S2_14_18  ( .A(\mult_19/ab[14][18] ), .B(
        \mult_19/CARRYB[13][18] ), .CI(\mult_19/SUMB[13][19] ), .CO(
        \mult_19/CARRYB[14][18] ), .S(\mult_19/SUMB[14][18] ) );
  FA_X1 \mult_19/S2_14_17  ( .A(\mult_19/ab[14][17] ), .B(
        \mult_19/CARRYB[13][17] ), .CI(\mult_19/SUMB[13][18] ), .CO(
        \mult_19/CARRYB[14][17] ), .S(\mult_19/SUMB[14][17] ) );
  FA_X1 \mult_19/S2_14_16  ( .A(\mult_19/ab[14][16] ), .B(
        \mult_19/CARRYB[13][16] ), .CI(\mult_19/SUMB[13][17] ), .CO(
        \mult_19/CARRYB[14][16] ), .S(\mult_19/SUMB[14][16] ) );
  FA_X1 \mult_19/S2_14_15  ( .A(\mult_19/ab[14][15] ), .B(
        \mult_19/CARRYB[13][15] ), .CI(\mult_19/SUMB[13][16] ), .CO(
        \mult_19/CARRYB[14][15] ), .S(\mult_19/SUMB[14][15] ) );
  FA_X1 \mult_19/S2_14_14  ( .A(\mult_19/ab[14][14] ), .B(
        \mult_19/CARRYB[13][14] ), .CI(\mult_19/SUMB[13][15] ), .CO(
        \mult_19/CARRYB[14][14] ), .S(\mult_19/SUMB[14][14] ) );
  FA_X1 \mult_19/S2_14_13  ( .A(\mult_19/ab[14][13] ), .B(
        \mult_19/CARRYB[13][13] ), .CI(\mult_19/SUMB[13][14] ), .CO(
        \mult_19/CARRYB[14][13] ), .S(\mult_19/SUMB[14][13] ) );
  FA_X1 \mult_19/S2_14_12  ( .A(\mult_19/ab[14][12] ), .B(
        \mult_19/CARRYB[13][12] ), .CI(\mult_19/SUMB[13][13] ), .CO(
        \mult_19/CARRYB[14][12] ), .S(\mult_19/SUMB[14][12] ) );
  FA_X1 \mult_19/S2_14_11  ( .A(\mult_19/ab[14][11] ), .B(
        \mult_19/CARRYB[13][11] ), .CI(\mult_19/SUMB[13][12] ), .CO(
        \mult_19/CARRYB[14][11] ), .S(\mult_19/SUMB[14][11] ) );
  FA_X1 \mult_19/S2_14_10  ( .A(\mult_19/ab[14][10] ), .B(
        \mult_19/CARRYB[13][10] ), .CI(\mult_19/SUMB[13][11] ), .CO(
        \mult_19/CARRYB[14][10] ), .S(\mult_19/SUMB[14][10] ) );
  FA_X1 \mult_19/S2_14_9  ( .A(\mult_19/ab[14][9] ), .B(
        \mult_19/CARRYB[13][9] ), .CI(\mult_19/SUMB[13][10] ), .CO(
        \mult_19/CARRYB[14][9] ), .S(\mult_19/SUMB[14][9] ) );
  FA_X1 \mult_19/S2_14_8  ( .A(\mult_19/ab[14][8] ), .B(
        \mult_19/CARRYB[13][8] ), .CI(\mult_19/SUMB[13][9] ), .CO(
        \mult_19/CARRYB[14][8] ), .S(\mult_19/SUMB[14][8] ) );
  FA_X1 \mult_19/S2_14_7  ( .A(\mult_19/ab[14][7] ), .B(
        \mult_19/CARRYB[13][7] ), .CI(\mult_19/SUMB[13][8] ), .CO(
        \mult_19/CARRYB[14][7] ), .S(\mult_19/SUMB[14][7] ) );
  FA_X1 \mult_19/S2_14_6  ( .A(\mult_19/ab[14][6] ), .B(
        \mult_19/CARRYB[13][6] ), .CI(\mult_19/SUMB[13][7] ), .CO(
        \mult_19/CARRYB[14][6] ), .S(\mult_19/SUMB[14][6] ) );
  FA_X1 \mult_19/S2_14_5  ( .A(\mult_19/ab[14][5] ), .B(
        \mult_19/CARRYB[13][5] ), .CI(\mult_19/SUMB[13][6] ), .CO(
        \mult_19/CARRYB[14][5] ), .S(\mult_19/SUMB[14][5] ) );
  FA_X1 \mult_19/S2_14_4  ( .A(\mult_19/ab[14][4] ), .B(
        \mult_19/CARRYB[13][4] ), .CI(\mult_19/SUMB[13][5] ), .CO(
        \mult_19/CARRYB[14][4] ), .S(\mult_19/SUMB[14][4] ) );
  FA_X1 \mult_19/S2_14_3  ( .A(\mult_19/ab[14][3] ), .B(
        \mult_19/CARRYB[13][3] ), .CI(\mult_19/SUMB[13][4] ), .CO(
        \mult_19/CARRYB[14][3] ), .S(\mult_19/SUMB[14][3] ) );
  FA_X1 \mult_19/S2_14_2  ( .A(\mult_19/ab[14][2] ), .B(
        \mult_19/CARRYB[13][2] ), .CI(\mult_19/SUMB[13][3] ), .CO(
        \mult_19/CARRYB[14][2] ), .S(\mult_19/SUMB[14][2] ) );
  FA_X1 \mult_19/S2_14_1  ( .A(\mult_19/ab[14][1] ), .B(
        \mult_19/CARRYB[13][1] ), .CI(\mult_19/SUMB[13][2] ), .CO(
        \mult_19/CARRYB[14][1] ), .S(\mult_19/SUMB[14][1] ) );
  FA_X1 \mult_19/S1_14_0  ( .A(\mult_19/ab[14][0] ), .B(
        \mult_19/CARRYB[13][0] ), .CI(\mult_19/SUMB[13][1] ), .CO(
        \mult_19/CARRYB[14][0] ), .S(N14) );
  FA_X1 \mult_19/S3_15_30  ( .A(\mult_19/ab[15][30] ), .B(
        \mult_19/CARRYB[14][30] ), .CI(\mult_19/ab[14][31] ), .CO(
        \mult_19/CARRYB[15][30] ), .S(\mult_19/SUMB[15][30] ) );
  FA_X1 \mult_19/S2_15_29  ( .A(\mult_19/ab[15][29] ), .B(
        \mult_19/CARRYB[14][29] ), .CI(\mult_19/SUMB[14][30] ), .CO(
        \mult_19/CARRYB[15][29] ), .S(\mult_19/SUMB[15][29] ) );
  FA_X1 \mult_19/S2_15_28  ( .A(\mult_19/ab[15][28] ), .B(
        \mult_19/CARRYB[14][28] ), .CI(\mult_19/SUMB[14][29] ), .CO(
        \mult_19/CARRYB[15][28] ), .S(\mult_19/SUMB[15][28] ) );
  FA_X1 \mult_19/S2_15_27  ( .A(\mult_19/ab[15][27] ), .B(
        \mult_19/CARRYB[14][27] ), .CI(\mult_19/SUMB[14][28] ), .CO(
        \mult_19/CARRYB[15][27] ), .S(\mult_19/SUMB[15][27] ) );
  FA_X1 \mult_19/S2_15_26  ( .A(\mult_19/ab[15][26] ), .B(
        \mult_19/CARRYB[14][26] ), .CI(\mult_19/SUMB[14][27] ), .CO(
        \mult_19/CARRYB[15][26] ), .S(\mult_19/SUMB[15][26] ) );
  FA_X1 \mult_19/S2_15_25  ( .A(\mult_19/ab[15][25] ), .B(
        \mult_19/CARRYB[14][25] ), .CI(\mult_19/SUMB[14][26] ), .CO(
        \mult_19/CARRYB[15][25] ), .S(\mult_19/SUMB[15][25] ) );
  FA_X1 \mult_19/S2_15_24  ( .A(\mult_19/ab[15][24] ), .B(
        \mult_19/CARRYB[14][24] ), .CI(\mult_19/SUMB[14][25] ), .CO(
        \mult_19/CARRYB[15][24] ), .S(\mult_19/SUMB[15][24] ) );
  FA_X1 \mult_19/S2_15_23  ( .A(\mult_19/ab[15][23] ), .B(
        \mult_19/CARRYB[14][23] ), .CI(\mult_19/SUMB[14][24] ), .CO(
        \mult_19/CARRYB[15][23] ), .S(\mult_19/SUMB[15][23] ) );
  FA_X1 \mult_19/S2_15_22  ( .A(\mult_19/ab[15][22] ), .B(
        \mult_19/CARRYB[14][22] ), .CI(\mult_19/SUMB[14][23] ), .CO(
        \mult_19/CARRYB[15][22] ), .S(\mult_19/SUMB[15][22] ) );
  FA_X1 \mult_19/S2_15_21  ( .A(\mult_19/ab[15][21] ), .B(
        \mult_19/CARRYB[14][21] ), .CI(\mult_19/SUMB[14][22] ), .CO(
        \mult_19/CARRYB[15][21] ), .S(\mult_19/SUMB[15][21] ) );
  FA_X1 \mult_19/S2_15_20  ( .A(\mult_19/ab[15][20] ), .B(
        \mult_19/CARRYB[14][20] ), .CI(\mult_19/SUMB[14][21] ), .CO(
        \mult_19/CARRYB[15][20] ), .S(\mult_19/SUMB[15][20] ) );
  FA_X1 \mult_19/S2_15_19  ( .A(\mult_19/ab[15][19] ), .B(
        \mult_19/CARRYB[14][19] ), .CI(\mult_19/SUMB[14][20] ), .CO(
        \mult_19/CARRYB[15][19] ), .S(\mult_19/SUMB[15][19] ) );
  FA_X1 \mult_19/S2_15_18  ( .A(\mult_19/ab[15][18] ), .B(
        \mult_19/CARRYB[14][18] ), .CI(\mult_19/SUMB[14][19] ), .CO(
        \mult_19/CARRYB[15][18] ), .S(\mult_19/SUMB[15][18] ) );
  FA_X1 \mult_19/S2_15_17  ( .A(\mult_19/ab[15][17] ), .B(
        \mult_19/CARRYB[14][17] ), .CI(\mult_19/SUMB[14][18] ), .CO(
        \mult_19/CARRYB[15][17] ), .S(\mult_19/SUMB[15][17] ) );
  FA_X1 \mult_19/S2_15_16  ( .A(\mult_19/ab[15][16] ), .B(
        \mult_19/CARRYB[14][16] ), .CI(\mult_19/SUMB[14][17] ), .CO(
        \mult_19/CARRYB[15][16] ), .S(\mult_19/SUMB[15][16] ) );
  FA_X1 \mult_19/S2_15_15  ( .A(\mult_19/ab[15][15] ), .B(
        \mult_19/CARRYB[14][15] ), .CI(\mult_19/SUMB[14][16] ), .CO(
        \mult_19/CARRYB[15][15] ), .S(\mult_19/SUMB[15][15] ) );
  FA_X1 \mult_19/S2_15_14  ( .A(\mult_19/ab[15][14] ), .B(
        \mult_19/CARRYB[14][14] ), .CI(\mult_19/SUMB[14][15] ), .CO(
        \mult_19/CARRYB[15][14] ), .S(\mult_19/SUMB[15][14] ) );
  FA_X1 \mult_19/S2_15_13  ( .A(\mult_19/ab[15][13] ), .B(
        \mult_19/CARRYB[14][13] ), .CI(\mult_19/SUMB[14][14] ), .CO(
        \mult_19/CARRYB[15][13] ), .S(\mult_19/SUMB[15][13] ) );
  FA_X1 \mult_19/S2_15_12  ( .A(\mult_19/ab[15][12] ), .B(
        \mult_19/CARRYB[14][12] ), .CI(\mult_19/SUMB[14][13] ), .CO(
        \mult_19/CARRYB[15][12] ), .S(\mult_19/SUMB[15][12] ) );
  FA_X1 \mult_19/S2_15_11  ( .A(\mult_19/ab[15][11] ), .B(
        \mult_19/CARRYB[14][11] ), .CI(\mult_19/SUMB[14][12] ), .CO(
        \mult_19/CARRYB[15][11] ), .S(\mult_19/SUMB[15][11] ) );
  FA_X1 \mult_19/S2_15_10  ( .A(\mult_19/ab[15][10] ), .B(
        \mult_19/CARRYB[14][10] ), .CI(\mult_19/SUMB[14][11] ), .CO(
        \mult_19/CARRYB[15][10] ), .S(\mult_19/SUMB[15][10] ) );
  FA_X1 \mult_19/S2_15_9  ( .A(\mult_19/ab[15][9] ), .B(
        \mult_19/CARRYB[14][9] ), .CI(\mult_19/SUMB[14][10] ), .CO(
        \mult_19/CARRYB[15][9] ), .S(\mult_19/SUMB[15][9] ) );
  FA_X1 \mult_19/S2_15_8  ( .A(\mult_19/ab[15][8] ), .B(
        \mult_19/CARRYB[14][8] ), .CI(\mult_19/SUMB[14][9] ), .CO(
        \mult_19/CARRYB[15][8] ), .S(\mult_19/SUMB[15][8] ) );
  FA_X1 \mult_19/S2_15_7  ( .A(\mult_19/ab[15][7] ), .B(
        \mult_19/CARRYB[14][7] ), .CI(\mult_19/SUMB[14][8] ), .CO(
        \mult_19/CARRYB[15][7] ), .S(\mult_19/SUMB[15][7] ) );
  FA_X1 \mult_19/S2_15_6  ( .A(\mult_19/ab[15][6] ), .B(
        \mult_19/CARRYB[14][6] ), .CI(\mult_19/SUMB[14][7] ), .CO(
        \mult_19/CARRYB[15][6] ), .S(\mult_19/SUMB[15][6] ) );
  FA_X1 \mult_19/S2_15_5  ( .A(\mult_19/ab[15][5] ), .B(
        \mult_19/CARRYB[14][5] ), .CI(\mult_19/SUMB[14][6] ), .CO(
        \mult_19/CARRYB[15][5] ), .S(\mult_19/SUMB[15][5] ) );
  FA_X1 \mult_19/S2_15_4  ( .A(\mult_19/ab[15][4] ), .B(
        \mult_19/CARRYB[14][4] ), .CI(\mult_19/SUMB[14][5] ), .CO(
        \mult_19/CARRYB[15][4] ), .S(\mult_19/SUMB[15][4] ) );
  FA_X1 \mult_19/S2_15_3  ( .A(\mult_19/ab[15][3] ), .B(
        \mult_19/CARRYB[14][3] ), .CI(\mult_19/SUMB[14][4] ), .CO(
        \mult_19/CARRYB[15][3] ), .S(\mult_19/SUMB[15][3] ) );
  FA_X1 \mult_19/S2_15_2  ( .A(\mult_19/ab[15][2] ), .B(
        \mult_19/CARRYB[14][2] ), .CI(\mult_19/SUMB[14][3] ), .CO(
        \mult_19/CARRYB[15][2] ), .S(\mult_19/SUMB[15][2] ) );
  FA_X1 \mult_19/S2_15_1  ( .A(\mult_19/ab[15][1] ), .B(
        \mult_19/CARRYB[14][1] ), .CI(\mult_19/SUMB[14][2] ), .CO(
        \mult_19/CARRYB[15][1] ), .S(\mult_19/SUMB[15][1] ) );
  FA_X1 \mult_19/S1_15_0  ( .A(\mult_19/ab[15][0] ), .B(
        \mult_19/CARRYB[14][0] ), .CI(\mult_19/SUMB[14][1] ), .CO(
        \mult_19/CARRYB[15][0] ), .S(N15) );
  FA_X1 \mult_19/S3_16_30  ( .A(\mult_19/ab[16][30] ), .B(
        \mult_19/CARRYB[15][30] ), .CI(\mult_19/ab[15][31] ), .CO(
        \mult_19/CARRYB[16][30] ), .S(\mult_19/SUMB[16][30] ) );
  FA_X1 \mult_19/S2_16_29  ( .A(\mult_19/ab[16][29] ), .B(
        \mult_19/CARRYB[15][29] ), .CI(\mult_19/SUMB[15][30] ), .CO(
        \mult_19/CARRYB[16][29] ), .S(\mult_19/SUMB[16][29] ) );
  FA_X1 \mult_19/S2_16_28  ( .A(\mult_19/ab[16][28] ), .B(
        \mult_19/CARRYB[15][28] ), .CI(\mult_19/SUMB[15][29] ), .CO(
        \mult_19/CARRYB[16][28] ), .S(\mult_19/SUMB[16][28] ) );
  FA_X1 \mult_19/S2_16_27  ( .A(\mult_19/ab[16][27] ), .B(
        \mult_19/CARRYB[15][27] ), .CI(\mult_19/SUMB[15][28] ), .CO(
        \mult_19/CARRYB[16][27] ), .S(\mult_19/SUMB[16][27] ) );
  FA_X1 \mult_19/S2_16_26  ( .A(\mult_19/ab[16][26] ), .B(
        \mult_19/CARRYB[15][26] ), .CI(\mult_19/SUMB[15][27] ), .CO(
        \mult_19/CARRYB[16][26] ), .S(\mult_19/SUMB[16][26] ) );
  FA_X1 \mult_19/S2_16_25  ( .A(\mult_19/ab[16][25] ), .B(
        \mult_19/CARRYB[15][25] ), .CI(\mult_19/SUMB[15][26] ), .CO(
        \mult_19/CARRYB[16][25] ), .S(\mult_19/SUMB[16][25] ) );
  FA_X1 \mult_19/S2_16_24  ( .A(\mult_19/ab[16][24] ), .B(
        \mult_19/CARRYB[15][24] ), .CI(\mult_19/SUMB[15][25] ), .CO(
        \mult_19/CARRYB[16][24] ), .S(\mult_19/SUMB[16][24] ) );
  FA_X1 \mult_19/S2_16_23  ( .A(\mult_19/ab[16][23] ), .B(
        \mult_19/CARRYB[15][23] ), .CI(\mult_19/SUMB[15][24] ), .CO(
        \mult_19/CARRYB[16][23] ), .S(\mult_19/SUMB[16][23] ) );
  FA_X1 \mult_19/S2_16_22  ( .A(\mult_19/ab[16][22] ), .B(
        \mult_19/CARRYB[15][22] ), .CI(\mult_19/SUMB[15][23] ), .CO(
        \mult_19/CARRYB[16][22] ), .S(\mult_19/SUMB[16][22] ) );
  FA_X1 \mult_19/S2_16_21  ( .A(\mult_19/ab[16][21] ), .B(
        \mult_19/CARRYB[15][21] ), .CI(\mult_19/SUMB[15][22] ), .CO(
        \mult_19/CARRYB[16][21] ), .S(\mult_19/SUMB[16][21] ) );
  FA_X1 \mult_19/S2_16_20  ( .A(\mult_19/ab[16][20] ), .B(
        \mult_19/CARRYB[15][20] ), .CI(\mult_19/SUMB[15][21] ), .CO(
        \mult_19/CARRYB[16][20] ), .S(\mult_19/SUMB[16][20] ) );
  FA_X1 \mult_19/S2_16_19  ( .A(\mult_19/ab[16][19] ), .B(
        \mult_19/CARRYB[15][19] ), .CI(\mult_19/SUMB[15][20] ), .CO(
        \mult_19/CARRYB[16][19] ), .S(\mult_19/SUMB[16][19] ) );
  FA_X1 \mult_19/S2_16_18  ( .A(\mult_19/ab[16][18] ), .B(
        \mult_19/CARRYB[15][18] ), .CI(\mult_19/SUMB[15][19] ), .CO(
        \mult_19/CARRYB[16][18] ), .S(\mult_19/SUMB[16][18] ) );
  FA_X1 \mult_19/S2_16_17  ( .A(\mult_19/ab[16][17] ), .B(
        \mult_19/CARRYB[15][17] ), .CI(\mult_19/SUMB[15][18] ), .CO(
        \mult_19/CARRYB[16][17] ), .S(\mult_19/SUMB[16][17] ) );
  FA_X1 \mult_19/S2_16_16  ( .A(\mult_19/ab[16][16] ), .B(
        \mult_19/CARRYB[15][16] ), .CI(\mult_19/SUMB[15][17] ), .CO(
        \mult_19/CARRYB[16][16] ), .S(\mult_19/SUMB[16][16] ) );
  FA_X1 \mult_19/S2_16_15  ( .A(\mult_19/ab[16][15] ), .B(
        \mult_19/CARRYB[15][15] ), .CI(\mult_19/SUMB[15][16] ), .CO(
        \mult_19/CARRYB[16][15] ), .S(\mult_19/SUMB[16][15] ) );
  FA_X1 \mult_19/S2_16_14  ( .A(\mult_19/ab[16][14] ), .B(
        \mult_19/CARRYB[15][14] ), .CI(\mult_19/SUMB[15][15] ), .CO(
        \mult_19/CARRYB[16][14] ), .S(\mult_19/SUMB[16][14] ) );
  FA_X1 \mult_19/S2_16_13  ( .A(\mult_19/ab[16][13] ), .B(
        \mult_19/CARRYB[15][13] ), .CI(\mult_19/SUMB[15][14] ), .CO(
        \mult_19/CARRYB[16][13] ), .S(\mult_19/SUMB[16][13] ) );
  FA_X1 \mult_19/S2_16_12  ( .A(\mult_19/ab[16][12] ), .B(
        \mult_19/CARRYB[15][12] ), .CI(\mult_19/SUMB[15][13] ), .CO(
        \mult_19/CARRYB[16][12] ), .S(\mult_19/SUMB[16][12] ) );
  FA_X1 \mult_19/S2_16_11  ( .A(\mult_19/ab[16][11] ), .B(
        \mult_19/CARRYB[15][11] ), .CI(\mult_19/SUMB[15][12] ), .CO(
        \mult_19/CARRYB[16][11] ), .S(\mult_19/SUMB[16][11] ) );
  FA_X1 \mult_19/S2_16_10  ( .A(\mult_19/ab[16][10] ), .B(
        \mult_19/CARRYB[15][10] ), .CI(\mult_19/SUMB[15][11] ), .CO(
        \mult_19/CARRYB[16][10] ), .S(\mult_19/SUMB[16][10] ) );
  FA_X1 \mult_19/S2_16_9  ( .A(\mult_19/ab[16][9] ), .B(
        \mult_19/CARRYB[15][9] ), .CI(\mult_19/SUMB[15][10] ), .CO(
        \mult_19/CARRYB[16][9] ), .S(\mult_19/SUMB[16][9] ) );
  FA_X1 \mult_19/S2_16_8  ( .A(\mult_19/ab[16][8] ), .B(
        \mult_19/CARRYB[15][8] ), .CI(\mult_19/SUMB[15][9] ), .CO(
        \mult_19/CARRYB[16][8] ), .S(\mult_19/SUMB[16][8] ) );
  FA_X1 \mult_19/S2_16_7  ( .A(\mult_19/ab[16][7] ), .B(
        \mult_19/CARRYB[15][7] ), .CI(\mult_19/SUMB[15][8] ), .CO(
        \mult_19/CARRYB[16][7] ), .S(\mult_19/SUMB[16][7] ) );
  FA_X1 \mult_19/S2_16_6  ( .A(\mult_19/ab[16][6] ), .B(
        \mult_19/CARRYB[15][6] ), .CI(\mult_19/SUMB[15][7] ), .CO(
        \mult_19/CARRYB[16][6] ), .S(\mult_19/SUMB[16][6] ) );
  FA_X1 \mult_19/S2_16_5  ( .A(\mult_19/ab[16][5] ), .B(
        \mult_19/CARRYB[15][5] ), .CI(\mult_19/SUMB[15][6] ), .CO(
        \mult_19/CARRYB[16][5] ), .S(\mult_19/SUMB[16][5] ) );
  FA_X1 \mult_19/S2_16_4  ( .A(\mult_19/ab[16][4] ), .B(
        \mult_19/CARRYB[15][4] ), .CI(\mult_19/SUMB[15][5] ), .CO(
        \mult_19/CARRYB[16][4] ), .S(\mult_19/SUMB[16][4] ) );
  FA_X1 \mult_19/S2_16_3  ( .A(\mult_19/ab[16][3] ), .B(
        \mult_19/CARRYB[15][3] ), .CI(\mult_19/SUMB[15][4] ), .CO(
        \mult_19/CARRYB[16][3] ), .S(\mult_19/SUMB[16][3] ) );
  FA_X1 \mult_19/S2_16_2  ( .A(\mult_19/ab[16][2] ), .B(
        \mult_19/CARRYB[15][2] ), .CI(\mult_19/SUMB[15][3] ), .CO(
        \mult_19/CARRYB[16][2] ), .S(\mult_19/SUMB[16][2] ) );
  FA_X1 \mult_19/S2_16_1  ( .A(\mult_19/ab[16][1] ), .B(
        \mult_19/CARRYB[15][1] ), .CI(\mult_19/SUMB[15][2] ), .CO(
        \mult_19/CARRYB[16][1] ), .S(\mult_19/SUMB[16][1] ) );
  FA_X1 \mult_19/S1_16_0  ( .A(\mult_19/ab[16][0] ), .B(
        \mult_19/CARRYB[15][0] ), .CI(\mult_19/SUMB[15][1] ), .CO(
        \mult_19/CARRYB[16][0] ), .S(N16) );
  FA_X1 \mult_19/S3_17_30  ( .A(\mult_19/ab[17][30] ), .B(
        \mult_19/CARRYB[16][30] ), .CI(\mult_19/ab[16][31] ), .CO(
        \mult_19/CARRYB[17][30] ), .S(\mult_19/SUMB[17][30] ) );
  FA_X1 \mult_19/S2_17_29  ( .A(\mult_19/ab[17][29] ), .B(
        \mult_19/CARRYB[16][29] ), .CI(\mult_19/SUMB[16][30] ), .CO(
        \mult_19/CARRYB[17][29] ), .S(\mult_19/SUMB[17][29] ) );
  FA_X1 \mult_19/S2_17_28  ( .A(\mult_19/ab[17][28] ), .B(
        \mult_19/CARRYB[16][28] ), .CI(\mult_19/SUMB[16][29] ), .CO(
        \mult_19/CARRYB[17][28] ), .S(\mult_19/SUMB[17][28] ) );
  FA_X1 \mult_19/S2_17_27  ( .A(\mult_19/ab[17][27] ), .B(
        \mult_19/CARRYB[16][27] ), .CI(\mult_19/SUMB[16][28] ), .CO(
        \mult_19/CARRYB[17][27] ), .S(\mult_19/SUMB[17][27] ) );
  FA_X1 \mult_19/S2_17_26  ( .A(\mult_19/ab[17][26] ), .B(
        \mult_19/CARRYB[16][26] ), .CI(\mult_19/SUMB[16][27] ), .CO(
        \mult_19/CARRYB[17][26] ), .S(\mult_19/SUMB[17][26] ) );
  FA_X1 \mult_19/S2_17_25  ( .A(\mult_19/ab[17][25] ), .B(
        \mult_19/CARRYB[16][25] ), .CI(\mult_19/SUMB[16][26] ), .CO(
        \mult_19/CARRYB[17][25] ), .S(\mult_19/SUMB[17][25] ) );
  FA_X1 \mult_19/S2_17_24  ( .A(\mult_19/ab[17][24] ), .B(
        \mult_19/CARRYB[16][24] ), .CI(\mult_19/SUMB[16][25] ), .CO(
        \mult_19/CARRYB[17][24] ), .S(\mult_19/SUMB[17][24] ) );
  FA_X1 \mult_19/S2_17_23  ( .A(\mult_19/ab[17][23] ), .B(
        \mult_19/CARRYB[16][23] ), .CI(\mult_19/SUMB[16][24] ), .CO(
        \mult_19/CARRYB[17][23] ), .S(\mult_19/SUMB[17][23] ) );
  FA_X1 \mult_19/S2_17_22  ( .A(\mult_19/ab[17][22] ), .B(
        \mult_19/CARRYB[16][22] ), .CI(\mult_19/SUMB[16][23] ), .CO(
        \mult_19/CARRYB[17][22] ), .S(\mult_19/SUMB[17][22] ) );
  FA_X1 \mult_19/S2_17_21  ( .A(\mult_19/ab[17][21] ), .B(
        \mult_19/CARRYB[16][21] ), .CI(\mult_19/SUMB[16][22] ), .CO(
        \mult_19/CARRYB[17][21] ), .S(\mult_19/SUMB[17][21] ) );
  FA_X1 \mult_19/S2_17_20  ( .A(\mult_19/ab[17][20] ), .B(
        \mult_19/CARRYB[16][20] ), .CI(\mult_19/SUMB[16][21] ), .CO(
        \mult_19/CARRYB[17][20] ), .S(\mult_19/SUMB[17][20] ) );
  FA_X1 \mult_19/S2_17_19  ( .A(\mult_19/ab[17][19] ), .B(
        \mult_19/CARRYB[16][19] ), .CI(\mult_19/SUMB[16][20] ), .CO(
        \mult_19/CARRYB[17][19] ), .S(\mult_19/SUMB[17][19] ) );
  FA_X1 \mult_19/S2_17_18  ( .A(\mult_19/ab[17][18] ), .B(
        \mult_19/CARRYB[16][18] ), .CI(\mult_19/SUMB[16][19] ), .CO(
        \mult_19/CARRYB[17][18] ), .S(\mult_19/SUMB[17][18] ) );
  FA_X1 \mult_19/S2_17_17  ( .A(\mult_19/ab[17][17] ), .B(
        \mult_19/CARRYB[16][17] ), .CI(\mult_19/SUMB[16][18] ), .CO(
        \mult_19/CARRYB[17][17] ), .S(\mult_19/SUMB[17][17] ) );
  FA_X1 \mult_19/S2_17_16  ( .A(\mult_19/ab[17][16] ), .B(
        \mult_19/CARRYB[16][16] ), .CI(\mult_19/SUMB[16][17] ), .CO(
        \mult_19/CARRYB[17][16] ), .S(\mult_19/SUMB[17][16] ) );
  FA_X1 \mult_19/S2_17_15  ( .A(\mult_19/ab[17][15] ), .B(
        \mult_19/CARRYB[16][15] ), .CI(\mult_19/SUMB[16][16] ), .CO(
        \mult_19/CARRYB[17][15] ), .S(\mult_19/SUMB[17][15] ) );
  FA_X1 \mult_19/S2_17_14  ( .A(\mult_19/ab[17][14] ), .B(
        \mult_19/CARRYB[16][14] ), .CI(\mult_19/SUMB[16][15] ), .CO(
        \mult_19/CARRYB[17][14] ), .S(\mult_19/SUMB[17][14] ) );
  FA_X1 \mult_19/S2_17_13  ( .A(\mult_19/ab[17][13] ), .B(
        \mult_19/CARRYB[16][13] ), .CI(\mult_19/SUMB[16][14] ), .CO(
        \mult_19/CARRYB[17][13] ), .S(\mult_19/SUMB[17][13] ) );
  FA_X1 \mult_19/S2_17_12  ( .A(\mult_19/ab[17][12] ), .B(
        \mult_19/CARRYB[16][12] ), .CI(\mult_19/SUMB[16][13] ), .CO(
        \mult_19/CARRYB[17][12] ), .S(\mult_19/SUMB[17][12] ) );
  FA_X1 \mult_19/S2_17_11  ( .A(\mult_19/ab[17][11] ), .B(
        \mult_19/CARRYB[16][11] ), .CI(\mult_19/SUMB[16][12] ), .CO(
        \mult_19/CARRYB[17][11] ), .S(\mult_19/SUMB[17][11] ) );
  FA_X1 \mult_19/S2_17_10  ( .A(\mult_19/ab[17][10] ), .B(
        \mult_19/CARRYB[16][10] ), .CI(\mult_19/SUMB[16][11] ), .CO(
        \mult_19/CARRYB[17][10] ), .S(\mult_19/SUMB[17][10] ) );
  FA_X1 \mult_19/S2_17_9  ( .A(\mult_19/ab[17][9] ), .B(
        \mult_19/CARRYB[16][9] ), .CI(\mult_19/SUMB[16][10] ), .CO(
        \mult_19/CARRYB[17][9] ), .S(\mult_19/SUMB[17][9] ) );
  FA_X1 \mult_19/S2_17_8  ( .A(\mult_19/ab[17][8] ), .B(
        \mult_19/CARRYB[16][8] ), .CI(\mult_19/SUMB[16][9] ), .CO(
        \mult_19/CARRYB[17][8] ), .S(\mult_19/SUMB[17][8] ) );
  FA_X1 \mult_19/S2_17_7  ( .A(\mult_19/ab[17][7] ), .B(
        \mult_19/CARRYB[16][7] ), .CI(\mult_19/SUMB[16][8] ), .CO(
        \mult_19/CARRYB[17][7] ), .S(\mult_19/SUMB[17][7] ) );
  FA_X1 \mult_19/S2_17_6  ( .A(\mult_19/ab[17][6] ), .B(
        \mult_19/CARRYB[16][6] ), .CI(\mult_19/SUMB[16][7] ), .CO(
        \mult_19/CARRYB[17][6] ), .S(\mult_19/SUMB[17][6] ) );
  FA_X1 \mult_19/S2_17_5  ( .A(\mult_19/ab[17][5] ), .B(
        \mult_19/CARRYB[16][5] ), .CI(\mult_19/SUMB[16][6] ), .CO(
        \mult_19/CARRYB[17][5] ), .S(\mult_19/SUMB[17][5] ) );
  FA_X1 \mult_19/S2_17_4  ( .A(\mult_19/ab[17][4] ), .B(
        \mult_19/CARRYB[16][4] ), .CI(\mult_19/SUMB[16][5] ), .CO(
        \mult_19/CARRYB[17][4] ), .S(\mult_19/SUMB[17][4] ) );
  FA_X1 \mult_19/S2_17_3  ( .A(\mult_19/ab[17][3] ), .B(
        \mult_19/CARRYB[16][3] ), .CI(\mult_19/SUMB[16][4] ), .CO(
        \mult_19/CARRYB[17][3] ), .S(\mult_19/SUMB[17][3] ) );
  FA_X1 \mult_19/S2_17_2  ( .A(\mult_19/ab[17][2] ), .B(
        \mult_19/CARRYB[16][2] ), .CI(\mult_19/SUMB[16][3] ), .CO(
        \mult_19/CARRYB[17][2] ), .S(\mult_19/SUMB[17][2] ) );
  FA_X1 \mult_19/S2_17_1  ( .A(\mult_19/ab[17][1] ), .B(
        \mult_19/CARRYB[16][1] ), .CI(\mult_19/SUMB[16][2] ), .CO(
        \mult_19/CARRYB[17][1] ), .S(\mult_19/SUMB[17][1] ) );
  FA_X1 \mult_19/S1_17_0  ( .A(\mult_19/ab[17][0] ), .B(
        \mult_19/CARRYB[16][0] ), .CI(\mult_19/SUMB[16][1] ), .CO(
        \mult_19/CARRYB[17][0] ), .S(N17) );
  FA_X1 \mult_19/S3_18_30  ( .A(\mult_19/ab[18][30] ), .B(
        \mult_19/CARRYB[17][30] ), .CI(\mult_19/ab[17][31] ), .CO(
        \mult_19/CARRYB[18][30] ), .S(\mult_19/SUMB[18][30] ) );
  FA_X1 \mult_19/S2_18_29  ( .A(\mult_19/ab[18][29] ), .B(
        \mult_19/CARRYB[17][29] ), .CI(\mult_19/SUMB[17][30] ), .CO(
        \mult_19/CARRYB[18][29] ), .S(\mult_19/SUMB[18][29] ) );
  FA_X1 \mult_19/S2_18_28  ( .A(\mult_19/ab[18][28] ), .B(
        \mult_19/CARRYB[17][28] ), .CI(\mult_19/SUMB[17][29] ), .CO(
        \mult_19/CARRYB[18][28] ), .S(\mult_19/SUMB[18][28] ) );
  FA_X1 \mult_19/S2_18_27  ( .A(\mult_19/ab[18][27] ), .B(
        \mult_19/CARRYB[17][27] ), .CI(\mult_19/SUMB[17][28] ), .CO(
        \mult_19/CARRYB[18][27] ), .S(\mult_19/SUMB[18][27] ) );
  FA_X1 \mult_19/S2_18_26  ( .A(\mult_19/ab[18][26] ), .B(
        \mult_19/CARRYB[17][26] ), .CI(\mult_19/SUMB[17][27] ), .CO(
        \mult_19/CARRYB[18][26] ), .S(\mult_19/SUMB[18][26] ) );
  FA_X1 \mult_19/S2_18_25  ( .A(\mult_19/ab[18][25] ), .B(
        \mult_19/CARRYB[17][25] ), .CI(\mult_19/SUMB[17][26] ), .CO(
        \mult_19/CARRYB[18][25] ), .S(\mult_19/SUMB[18][25] ) );
  FA_X1 \mult_19/S2_18_24  ( .A(\mult_19/ab[18][24] ), .B(
        \mult_19/CARRYB[17][24] ), .CI(\mult_19/SUMB[17][25] ), .CO(
        \mult_19/CARRYB[18][24] ), .S(\mult_19/SUMB[18][24] ) );
  FA_X1 \mult_19/S2_18_23  ( .A(\mult_19/ab[18][23] ), .B(
        \mult_19/CARRYB[17][23] ), .CI(\mult_19/SUMB[17][24] ), .CO(
        \mult_19/CARRYB[18][23] ), .S(\mult_19/SUMB[18][23] ) );
  FA_X1 \mult_19/S2_18_22  ( .A(\mult_19/ab[18][22] ), .B(
        \mult_19/CARRYB[17][22] ), .CI(\mult_19/SUMB[17][23] ), .CO(
        \mult_19/CARRYB[18][22] ), .S(\mult_19/SUMB[18][22] ) );
  FA_X1 \mult_19/S2_18_21  ( .A(\mult_19/ab[18][21] ), .B(
        \mult_19/CARRYB[17][21] ), .CI(\mult_19/SUMB[17][22] ), .CO(
        \mult_19/CARRYB[18][21] ), .S(\mult_19/SUMB[18][21] ) );
  FA_X1 \mult_19/S2_18_20  ( .A(\mult_19/ab[18][20] ), .B(
        \mult_19/CARRYB[17][20] ), .CI(\mult_19/SUMB[17][21] ), .CO(
        \mult_19/CARRYB[18][20] ), .S(\mult_19/SUMB[18][20] ) );
  FA_X1 \mult_19/S2_18_19  ( .A(\mult_19/ab[18][19] ), .B(
        \mult_19/CARRYB[17][19] ), .CI(\mult_19/SUMB[17][20] ), .CO(
        \mult_19/CARRYB[18][19] ), .S(\mult_19/SUMB[18][19] ) );
  FA_X1 \mult_19/S2_18_18  ( .A(\mult_19/ab[18][18] ), .B(
        \mult_19/CARRYB[17][18] ), .CI(\mult_19/SUMB[17][19] ), .CO(
        \mult_19/CARRYB[18][18] ), .S(\mult_19/SUMB[18][18] ) );
  FA_X1 \mult_19/S2_18_17  ( .A(\mult_19/ab[18][17] ), .B(
        \mult_19/CARRYB[17][17] ), .CI(\mult_19/SUMB[17][18] ), .CO(
        \mult_19/CARRYB[18][17] ), .S(\mult_19/SUMB[18][17] ) );
  FA_X1 \mult_19/S2_18_16  ( .A(\mult_19/ab[18][16] ), .B(
        \mult_19/CARRYB[17][16] ), .CI(\mult_19/SUMB[17][17] ), .CO(
        \mult_19/CARRYB[18][16] ), .S(\mult_19/SUMB[18][16] ) );
  FA_X1 \mult_19/S2_18_15  ( .A(\mult_19/ab[18][15] ), .B(
        \mult_19/CARRYB[17][15] ), .CI(\mult_19/SUMB[17][16] ), .CO(
        \mult_19/CARRYB[18][15] ), .S(\mult_19/SUMB[18][15] ) );
  FA_X1 \mult_19/S2_18_14  ( .A(\mult_19/ab[18][14] ), .B(
        \mult_19/CARRYB[17][14] ), .CI(\mult_19/SUMB[17][15] ), .CO(
        \mult_19/CARRYB[18][14] ), .S(\mult_19/SUMB[18][14] ) );
  FA_X1 \mult_19/S2_18_13  ( .A(\mult_19/ab[18][13] ), .B(
        \mult_19/CARRYB[17][13] ), .CI(\mult_19/SUMB[17][14] ), .CO(
        \mult_19/CARRYB[18][13] ), .S(\mult_19/SUMB[18][13] ) );
  FA_X1 \mult_19/S2_18_12  ( .A(\mult_19/ab[18][12] ), .B(
        \mult_19/CARRYB[17][12] ), .CI(\mult_19/SUMB[17][13] ), .CO(
        \mult_19/CARRYB[18][12] ), .S(\mult_19/SUMB[18][12] ) );
  FA_X1 \mult_19/S2_18_11  ( .A(\mult_19/ab[18][11] ), .B(
        \mult_19/CARRYB[17][11] ), .CI(\mult_19/SUMB[17][12] ), .CO(
        \mult_19/CARRYB[18][11] ), .S(\mult_19/SUMB[18][11] ) );
  FA_X1 \mult_19/S2_18_10  ( .A(\mult_19/ab[18][10] ), .B(
        \mult_19/CARRYB[17][10] ), .CI(\mult_19/SUMB[17][11] ), .CO(
        \mult_19/CARRYB[18][10] ), .S(\mult_19/SUMB[18][10] ) );
  FA_X1 \mult_19/S2_18_9  ( .A(\mult_19/ab[18][9] ), .B(
        \mult_19/CARRYB[17][9] ), .CI(\mult_19/SUMB[17][10] ), .CO(
        \mult_19/CARRYB[18][9] ), .S(\mult_19/SUMB[18][9] ) );
  FA_X1 \mult_19/S2_18_8  ( .A(\mult_19/ab[18][8] ), .B(
        \mult_19/CARRYB[17][8] ), .CI(\mult_19/SUMB[17][9] ), .CO(
        \mult_19/CARRYB[18][8] ), .S(\mult_19/SUMB[18][8] ) );
  FA_X1 \mult_19/S2_18_7  ( .A(\mult_19/ab[18][7] ), .B(
        \mult_19/CARRYB[17][7] ), .CI(\mult_19/SUMB[17][8] ), .CO(
        \mult_19/CARRYB[18][7] ), .S(\mult_19/SUMB[18][7] ) );
  FA_X1 \mult_19/S2_18_6  ( .A(\mult_19/ab[18][6] ), .B(
        \mult_19/CARRYB[17][6] ), .CI(\mult_19/SUMB[17][7] ), .CO(
        \mult_19/CARRYB[18][6] ), .S(\mult_19/SUMB[18][6] ) );
  FA_X1 \mult_19/S2_18_5  ( .A(\mult_19/ab[18][5] ), .B(
        \mult_19/CARRYB[17][5] ), .CI(\mult_19/SUMB[17][6] ), .CO(
        \mult_19/CARRYB[18][5] ), .S(\mult_19/SUMB[18][5] ) );
  FA_X1 \mult_19/S2_18_4  ( .A(\mult_19/ab[18][4] ), .B(
        \mult_19/CARRYB[17][4] ), .CI(\mult_19/SUMB[17][5] ), .CO(
        \mult_19/CARRYB[18][4] ), .S(\mult_19/SUMB[18][4] ) );
  FA_X1 \mult_19/S2_18_3  ( .A(\mult_19/ab[18][3] ), .B(
        \mult_19/CARRYB[17][3] ), .CI(\mult_19/SUMB[17][4] ), .CO(
        \mult_19/CARRYB[18][3] ), .S(\mult_19/SUMB[18][3] ) );
  FA_X1 \mult_19/S2_18_2  ( .A(\mult_19/ab[18][2] ), .B(
        \mult_19/CARRYB[17][2] ), .CI(\mult_19/SUMB[17][3] ), .CO(
        \mult_19/CARRYB[18][2] ), .S(\mult_19/SUMB[18][2] ) );
  FA_X1 \mult_19/S2_18_1  ( .A(\mult_19/ab[18][1] ), .B(
        \mult_19/CARRYB[17][1] ), .CI(\mult_19/SUMB[17][2] ), .CO(
        \mult_19/CARRYB[18][1] ), .S(\mult_19/SUMB[18][1] ) );
  FA_X1 \mult_19/S1_18_0  ( .A(\mult_19/ab[18][0] ), .B(
        \mult_19/CARRYB[17][0] ), .CI(\mult_19/SUMB[17][1] ), .CO(
        \mult_19/CARRYB[18][0] ), .S(N18) );
  FA_X1 \mult_19/S3_19_30  ( .A(\mult_19/ab[19][30] ), .B(
        \mult_19/CARRYB[18][30] ), .CI(\mult_19/ab[18][31] ), .CO(
        \mult_19/CARRYB[19][30] ), .S(\mult_19/SUMB[19][30] ) );
  FA_X1 \mult_19/S2_19_29  ( .A(\mult_19/ab[19][29] ), .B(
        \mult_19/CARRYB[18][29] ), .CI(\mult_19/SUMB[18][30] ), .CO(
        \mult_19/CARRYB[19][29] ), .S(\mult_19/SUMB[19][29] ) );
  FA_X1 \mult_19/S2_19_28  ( .A(\mult_19/ab[19][28] ), .B(
        \mult_19/CARRYB[18][28] ), .CI(\mult_19/SUMB[18][29] ), .CO(
        \mult_19/CARRYB[19][28] ), .S(\mult_19/SUMB[19][28] ) );
  FA_X1 \mult_19/S2_19_27  ( .A(\mult_19/ab[19][27] ), .B(
        \mult_19/CARRYB[18][27] ), .CI(\mult_19/SUMB[18][28] ), .CO(
        \mult_19/CARRYB[19][27] ), .S(\mult_19/SUMB[19][27] ) );
  FA_X1 \mult_19/S2_19_26  ( .A(\mult_19/ab[19][26] ), .B(
        \mult_19/CARRYB[18][26] ), .CI(\mult_19/SUMB[18][27] ), .CO(
        \mult_19/CARRYB[19][26] ), .S(\mult_19/SUMB[19][26] ) );
  FA_X1 \mult_19/S2_19_25  ( .A(\mult_19/ab[19][25] ), .B(
        \mult_19/CARRYB[18][25] ), .CI(\mult_19/SUMB[18][26] ), .CO(
        \mult_19/CARRYB[19][25] ), .S(\mult_19/SUMB[19][25] ) );
  FA_X1 \mult_19/S2_19_24  ( .A(\mult_19/ab[19][24] ), .B(
        \mult_19/CARRYB[18][24] ), .CI(\mult_19/SUMB[18][25] ), .CO(
        \mult_19/CARRYB[19][24] ), .S(\mult_19/SUMB[19][24] ) );
  FA_X1 \mult_19/S2_19_23  ( .A(\mult_19/ab[19][23] ), .B(
        \mult_19/CARRYB[18][23] ), .CI(\mult_19/SUMB[18][24] ), .CO(
        \mult_19/CARRYB[19][23] ), .S(\mult_19/SUMB[19][23] ) );
  FA_X1 \mult_19/S2_19_22  ( .A(\mult_19/ab[19][22] ), .B(
        \mult_19/CARRYB[18][22] ), .CI(\mult_19/SUMB[18][23] ), .CO(
        \mult_19/CARRYB[19][22] ), .S(\mult_19/SUMB[19][22] ) );
  FA_X1 \mult_19/S2_19_21  ( .A(\mult_19/ab[19][21] ), .B(
        \mult_19/CARRYB[18][21] ), .CI(\mult_19/SUMB[18][22] ), .CO(
        \mult_19/CARRYB[19][21] ), .S(\mult_19/SUMB[19][21] ) );
  FA_X1 \mult_19/S2_19_20  ( .A(\mult_19/ab[19][20] ), .B(
        \mult_19/CARRYB[18][20] ), .CI(\mult_19/SUMB[18][21] ), .CO(
        \mult_19/CARRYB[19][20] ), .S(\mult_19/SUMB[19][20] ) );
  FA_X1 \mult_19/S2_19_19  ( .A(\mult_19/ab[19][19] ), .B(
        \mult_19/CARRYB[18][19] ), .CI(\mult_19/SUMB[18][20] ), .CO(
        \mult_19/CARRYB[19][19] ), .S(\mult_19/SUMB[19][19] ) );
  FA_X1 \mult_19/S2_19_18  ( .A(\mult_19/ab[19][18] ), .B(
        \mult_19/CARRYB[18][18] ), .CI(\mult_19/SUMB[18][19] ), .CO(
        \mult_19/CARRYB[19][18] ), .S(\mult_19/SUMB[19][18] ) );
  FA_X1 \mult_19/S2_19_17  ( .A(\mult_19/ab[19][17] ), .B(
        \mult_19/CARRYB[18][17] ), .CI(\mult_19/SUMB[18][18] ), .CO(
        \mult_19/CARRYB[19][17] ), .S(\mult_19/SUMB[19][17] ) );
  FA_X1 \mult_19/S2_19_16  ( .A(\mult_19/ab[19][16] ), .B(
        \mult_19/CARRYB[18][16] ), .CI(\mult_19/SUMB[18][17] ), .CO(
        \mult_19/CARRYB[19][16] ), .S(\mult_19/SUMB[19][16] ) );
  FA_X1 \mult_19/S2_19_15  ( .A(\mult_19/ab[19][15] ), .B(
        \mult_19/CARRYB[18][15] ), .CI(\mult_19/SUMB[18][16] ), .CO(
        \mult_19/CARRYB[19][15] ), .S(\mult_19/SUMB[19][15] ) );
  FA_X1 \mult_19/S2_19_14  ( .A(\mult_19/ab[19][14] ), .B(
        \mult_19/CARRYB[18][14] ), .CI(\mult_19/SUMB[18][15] ), .CO(
        \mult_19/CARRYB[19][14] ), .S(\mult_19/SUMB[19][14] ) );
  FA_X1 \mult_19/S2_19_13  ( .A(\mult_19/ab[19][13] ), .B(
        \mult_19/CARRYB[18][13] ), .CI(\mult_19/SUMB[18][14] ), .CO(
        \mult_19/CARRYB[19][13] ), .S(\mult_19/SUMB[19][13] ) );
  FA_X1 \mult_19/S2_19_12  ( .A(\mult_19/ab[19][12] ), .B(
        \mult_19/CARRYB[18][12] ), .CI(\mult_19/SUMB[18][13] ), .CO(
        \mult_19/CARRYB[19][12] ), .S(\mult_19/SUMB[19][12] ) );
  FA_X1 \mult_19/S2_19_11  ( .A(\mult_19/ab[19][11] ), .B(
        \mult_19/CARRYB[18][11] ), .CI(\mult_19/SUMB[18][12] ), .CO(
        \mult_19/CARRYB[19][11] ), .S(\mult_19/SUMB[19][11] ) );
  FA_X1 \mult_19/S2_19_10  ( .A(\mult_19/ab[19][10] ), .B(
        \mult_19/CARRYB[18][10] ), .CI(\mult_19/SUMB[18][11] ), .CO(
        \mult_19/CARRYB[19][10] ), .S(\mult_19/SUMB[19][10] ) );
  FA_X1 \mult_19/S2_19_9  ( .A(\mult_19/ab[19][9] ), .B(
        \mult_19/CARRYB[18][9] ), .CI(\mult_19/SUMB[18][10] ), .CO(
        \mult_19/CARRYB[19][9] ), .S(\mult_19/SUMB[19][9] ) );
  FA_X1 \mult_19/S2_19_8  ( .A(\mult_19/ab[19][8] ), .B(
        \mult_19/CARRYB[18][8] ), .CI(\mult_19/SUMB[18][9] ), .CO(
        \mult_19/CARRYB[19][8] ), .S(\mult_19/SUMB[19][8] ) );
  FA_X1 \mult_19/S2_19_7  ( .A(\mult_19/ab[19][7] ), .B(
        \mult_19/CARRYB[18][7] ), .CI(\mult_19/SUMB[18][8] ), .CO(
        \mult_19/CARRYB[19][7] ), .S(\mult_19/SUMB[19][7] ) );
  FA_X1 \mult_19/S2_19_6  ( .A(\mult_19/ab[19][6] ), .B(
        \mult_19/CARRYB[18][6] ), .CI(\mult_19/SUMB[18][7] ), .CO(
        \mult_19/CARRYB[19][6] ), .S(\mult_19/SUMB[19][6] ) );
  FA_X1 \mult_19/S2_19_5  ( .A(\mult_19/ab[19][5] ), .B(
        \mult_19/CARRYB[18][5] ), .CI(\mult_19/SUMB[18][6] ), .CO(
        \mult_19/CARRYB[19][5] ), .S(\mult_19/SUMB[19][5] ) );
  FA_X1 \mult_19/S2_19_4  ( .A(\mult_19/ab[19][4] ), .B(
        \mult_19/CARRYB[18][4] ), .CI(\mult_19/SUMB[18][5] ), .CO(
        \mult_19/CARRYB[19][4] ), .S(\mult_19/SUMB[19][4] ) );
  FA_X1 \mult_19/S2_19_3  ( .A(\mult_19/ab[19][3] ), .B(
        \mult_19/CARRYB[18][3] ), .CI(\mult_19/SUMB[18][4] ), .CO(
        \mult_19/CARRYB[19][3] ), .S(\mult_19/SUMB[19][3] ) );
  FA_X1 \mult_19/S2_19_2  ( .A(\mult_19/ab[19][2] ), .B(
        \mult_19/CARRYB[18][2] ), .CI(\mult_19/SUMB[18][3] ), .CO(
        \mult_19/CARRYB[19][2] ), .S(\mult_19/SUMB[19][2] ) );
  FA_X1 \mult_19/S2_19_1  ( .A(\mult_19/ab[19][1] ), .B(
        \mult_19/CARRYB[18][1] ), .CI(\mult_19/SUMB[18][2] ), .CO(
        \mult_19/CARRYB[19][1] ), .S(\mult_19/SUMB[19][1] ) );
  FA_X1 \mult_19/S1_19_0  ( .A(\mult_19/ab[19][0] ), .B(
        \mult_19/CARRYB[18][0] ), .CI(\mult_19/SUMB[18][1] ), .CO(
        \mult_19/CARRYB[19][0] ), .S(N19) );
  FA_X1 \mult_19/S3_20_30  ( .A(\mult_19/ab[20][30] ), .B(
        \mult_19/CARRYB[19][30] ), .CI(\mult_19/ab[19][31] ), .CO(
        \mult_19/CARRYB[20][30] ), .S(\mult_19/SUMB[20][30] ) );
  FA_X1 \mult_19/S2_20_29  ( .A(\mult_19/ab[20][29] ), .B(
        \mult_19/CARRYB[19][29] ), .CI(\mult_19/SUMB[19][30] ), .CO(
        \mult_19/CARRYB[20][29] ), .S(\mult_19/SUMB[20][29] ) );
  FA_X1 \mult_19/S2_20_28  ( .A(\mult_19/ab[20][28] ), .B(
        \mult_19/CARRYB[19][28] ), .CI(\mult_19/SUMB[19][29] ), .CO(
        \mult_19/CARRYB[20][28] ), .S(\mult_19/SUMB[20][28] ) );
  FA_X1 \mult_19/S2_20_27  ( .A(\mult_19/ab[20][27] ), .B(
        \mult_19/CARRYB[19][27] ), .CI(\mult_19/SUMB[19][28] ), .CO(
        \mult_19/CARRYB[20][27] ), .S(\mult_19/SUMB[20][27] ) );
  FA_X1 \mult_19/S2_20_26  ( .A(\mult_19/ab[20][26] ), .B(
        \mult_19/CARRYB[19][26] ), .CI(\mult_19/SUMB[19][27] ), .CO(
        \mult_19/CARRYB[20][26] ), .S(\mult_19/SUMB[20][26] ) );
  FA_X1 \mult_19/S2_20_25  ( .A(\mult_19/ab[20][25] ), .B(
        \mult_19/CARRYB[19][25] ), .CI(\mult_19/SUMB[19][26] ), .CO(
        \mult_19/CARRYB[20][25] ), .S(\mult_19/SUMB[20][25] ) );
  FA_X1 \mult_19/S2_20_24  ( .A(\mult_19/ab[20][24] ), .B(
        \mult_19/CARRYB[19][24] ), .CI(\mult_19/SUMB[19][25] ), .CO(
        \mult_19/CARRYB[20][24] ), .S(\mult_19/SUMB[20][24] ) );
  FA_X1 \mult_19/S2_20_23  ( .A(\mult_19/ab[20][23] ), .B(
        \mult_19/CARRYB[19][23] ), .CI(\mult_19/SUMB[19][24] ), .CO(
        \mult_19/CARRYB[20][23] ), .S(\mult_19/SUMB[20][23] ) );
  FA_X1 \mult_19/S2_20_22  ( .A(\mult_19/ab[20][22] ), .B(
        \mult_19/CARRYB[19][22] ), .CI(\mult_19/SUMB[19][23] ), .CO(
        \mult_19/CARRYB[20][22] ), .S(\mult_19/SUMB[20][22] ) );
  FA_X1 \mult_19/S2_20_21  ( .A(\mult_19/ab[20][21] ), .B(
        \mult_19/CARRYB[19][21] ), .CI(\mult_19/SUMB[19][22] ), .CO(
        \mult_19/CARRYB[20][21] ), .S(\mult_19/SUMB[20][21] ) );
  FA_X1 \mult_19/S2_20_20  ( .A(\mult_19/ab[20][20] ), .B(
        \mult_19/CARRYB[19][20] ), .CI(\mult_19/SUMB[19][21] ), .CO(
        \mult_19/CARRYB[20][20] ), .S(\mult_19/SUMB[20][20] ) );
  FA_X1 \mult_19/S2_20_19  ( .A(\mult_19/ab[20][19] ), .B(
        \mult_19/CARRYB[19][19] ), .CI(\mult_19/SUMB[19][20] ), .CO(
        \mult_19/CARRYB[20][19] ), .S(\mult_19/SUMB[20][19] ) );
  FA_X1 \mult_19/S2_20_18  ( .A(\mult_19/ab[20][18] ), .B(
        \mult_19/CARRYB[19][18] ), .CI(\mult_19/SUMB[19][19] ), .CO(
        \mult_19/CARRYB[20][18] ), .S(\mult_19/SUMB[20][18] ) );
  FA_X1 \mult_19/S2_20_17  ( .A(\mult_19/ab[20][17] ), .B(
        \mult_19/CARRYB[19][17] ), .CI(\mult_19/SUMB[19][18] ), .CO(
        \mult_19/CARRYB[20][17] ), .S(\mult_19/SUMB[20][17] ) );
  FA_X1 \mult_19/S2_20_16  ( .A(\mult_19/ab[20][16] ), .B(
        \mult_19/CARRYB[19][16] ), .CI(\mult_19/SUMB[19][17] ), .CO(
        \mult_19/CARRYB[20][16] ), .S(\mult_19/SUMB[20][16] ) );
  FA_X1 \mult_19/S2_20_15  ( .A(\mult_19/ab[20][15] ), .B(
        \mult_19/CARRYB[19][15] ), .CI(\mult_19/SUMB[19][16] ), .CO(
        \mult_19/CARRYB[20][15] ), .S(\mult_19/SUMB[20][15] ) );
  FA_X1 \mult_19/S2_20_14  ( .A(\mult_19/ab[20][14] ), .B(
        \mult_19/CARRYB[19][14] ), .CI(\mult_19/SUMB[19][15] ), .CO(
        \mult_19/CARRYB[20][14] ), .S(\mult_19/SUMB[20][14] ) );
  FA_X1 \mult_19/S2_20_13  ( .A(\mult_19/ab[20][13] ), .B(
        \mult_19/CARRYB[19][13] ), .CI(\mult_19/SUMB[19][14] ), .CO(
        \mult_19/CARRYB[20][13] ), .S(\mult_19/SUMB[20][13] ) );
  FA_X1 \mult_19/S2_20_12  ( .A(\mult_19/ab[20][12] ), .B(
        \mult_19/CARRYB[19][12] ), .CI(\mult_19/SUMB[19][13] ), .CO(
        \mult_19/CARRYB[20][12] ), .S(\mult_19/SUMB[20][12] ) );
  FA_X1 \mult_19/S2_20_11  ( .A(\mult_19/ab[20][11] ), .B(
        \mult_19/CARRYB[19][11] ), .CI(\mult_19/SUMB[19][12] ), .CO(
        \mult_19/CARRYB[20][11] ), .S(\mult_19/SUMB[20][11] ) );
  FA_X1 \mult_19/S2_20_10  ( .A(\mult_19/ab[20][10] ), .B(
        \mult_19/CARRYB[19][10] ), .CI(\mult_19/SUMB[19][11] ), .CO(
        \mult_19/CARRYB[20][10] ), .S(\mult_19/SUMB[20][10] ) );
  FA_X1 \mult_19/S2_20_9  ( .A(\mult_19/ab[20][9] ), .B(
        \mult_19/CARRYB[19][9] ), .CI(\mult_19/SUMB[19][10] ), .CO(
        \mult_19/CARRYB[20][9] ), .S(\mult_19/SUMB[20][9] ) );
  FA_X1 \mult_19/S2_20_8  ( .A(\mult_19/ab[20][8] ), .B(
        \mult_19/CARRYB[19][8] ), .CI(\mult_19/SUMB[19][9] ), .CO(
        \mult_19/CARRYB[20][8] ), .S(\mult_19/SUMB[20][8] ) );
  FA_X1 \mult_19/S2_20_7  ( .A(\mult_19/ab[20][7] ), .B(
        \mult_19/CARRYB[19][7] ), .CI(\mult_19/SUMB[19][8] ), .CO(
        \mult_19/CARRYB[20][7] ), .S(\mult_19/SUMB[20][7] ) );
  FA_X1 \mult_19/S2_20_6  ( .A(\mult_19/ab[20][6] ), .B(
        \mult_19/CARRYB[19][6] ), .CI(\mult_19/SUMB[19][7] ), .CO(
        \mult_19/CARRYB[20][6] ), .S(\mult_19/SUMB[20][6] ) );
  FA_X1 \mult_19/S2_20_5  ( .A(\mult_19/ab[20][5] ), .B(
        \mult_19/CARRYB[19][5] ), .CI(\mult_19/SUMB[19][6] ), .CO(
        \mult_19/CARRYB[20][5] ), .S(\mult_19/SUMB[20][5] ) );
  FA_X1 \mult_19/S2_20_4  ( .A(\mult_19/ab[20][4] ), .B(
        \mult_19/CARRYB[19][4] ), .CI(\mult_19/SUMB[19][5] ), .CO(
        \mult_19/CARRYB[20][4] ), .S(\mult_19/SUMB[20][4] ) );
  FA_X1 \mult_19/S2_20_3  ( .A(\mult_19/ab[20][3] ), .B(
        \mult_19/CARRYB[19][3] ), .CI(\mult_19/SUMB[19][4] ), .CO(
        \mult_19/CARRYB[20][3] ), .S(\mult_19/SUMB[20][3] ) );
  FA_X1 \mult_19/S2_20_2  ( .A(\mult_19/ab[20][2] ), .B(
        \mult_19/CARRYB[19][2] ), .CI(\mult_19/SUMB[19][3] ), .CO(
        \mult_19/CARRYB[20][2] ), .S(\mult_19/SUMB[20][2] ) );
  FA_X1 \mult_19/S2_20_1  ( .A(\mult_19/ab[20][1] ), .B(
        \mult_19/CARRYB[19][1] ), .CI(\mult_19/SUMB[19][2] ), .CO(
        \mult_19/CARRYB[20][1] ), .S(\mult_19/SUMB[20][1] ) );
  FA_X1 \mult_19/S1_20_0  ( .A(\mult_19/ab[20][0] ), .B(
        \mult_19/CARRYB[19][0] ), .CI(\mult_19/SUMB[19][1] ), .CO(
        \mult_19/CARRYB[20][0] ), .S(N20) );
  FA_X1 \mult_19/S3_21_30  ( .A(\mult_19/ab[21][30] ), .B(
        \mult_19/CARRYB[20][30] ), .CI(\mult_19/ab[20][31] ), .CO(
        \mult_19/CARRYB[21][30] ), .S(\mult_19/SUMB[21][30] ) );
  FA_X1 \mult_19/S2_21_29  ( .A(\mult_19/ab[21][29] ), .B(
        \mult_19/CARRYB[20][29] ), .CI(\mult_19/SUMB[20][30] ), .CO(
        \mult_19/CARRYB[21][29] ), .S(\mult_19/SUMB[21][29] ) );
  FA_X1 \mult_19/S2_21_28  ( .A(\mult_19/ab[21][28] ), .B(
        \mult_19/CARRYB[20][28] ), .CI(\mult_19/SUMB[20][29] ), .CO(
        \mult_19/CARRYB[21][28] ), .S(\mult_19/SUMB[21][28] ) );
  FA_X1 \mult_19/S2_21_27  ( .A(\mult_19/ab[21][27] ), .B(
        \mult_19/CARRYB[20][27] ), .CI(\mult_19/SUMB[20][28] ), .CO(
        \mult_19/CARRYB[21][27] ), .S(\mult_19/SUMB[21][27] ) );
  FA_X1 \mult_19/S2_21_26  ( .A(\mult_19/ab[21][26] ), .B(
        \mult_19/CARRYB[20][26] ), .CI(\mult_19/SUMB[20][27] ), .CO(
        \mult_19/CARRYB[21][26] ), .S(\mult_19/SUMB[21][26] ) );
  FA_X1 \mult_19/S2_21_25  ( .A(\mult_19/ab[21][25] ), .B(
        \mult_19/CARRYB[20][25] ), .CI(\mult_19/SUMB[20][26] ), .CO(
        \mult_19/CARRYB[21][25] ), .S(\mult_19/SUMB[21][25] ) );
  FA_X1 \mult_19/S2_21_24  ( .A(\mult_19/ab[21][24] ), .B(
        \mult_19/CARRYB[20][24] ), .CI(\mult_19/SUMB[20][25] ), .CO(
        \mult_19/CARRYB[21][24] ), .S(\mult_19/SUMB[21][24] ) );
  FA_X1 \mult_19/S2_21_23  ( .A(\mult_19/ab[21][23] ), .B(
        \mult_19/CARRYB[20][23] ), .CI(\mult_19/SUMB[20][24] ), .CO(
        \mult_19/CARRYB[21][23] ), .S(\mult_19/SUMB[21][23] ) );
  FA_X1 \mult_19/S2_21_22  ( .A(\mult_19/ab[21][22] ), .B(
        \mult_19/CARRYB[20][22] ), .CI(\mult_19/SUMB[20][23] ), .CO(
        \mult_19/CARRYB[21][22] ), .S(\mult_19/SUMB[21][22] ) );
  FA_X1 \mult_19/S2_21_21  ( .A(\mult_19/ab[21][21] ), .B(
        \mult_19/CARRYB[20][21] ), .CI(\mult_19/SUMB[20][22] ), .CO(
        \mult_19/CARRYB[21][21] ), .S(\mult_19/SUMB[21][21] ) );
  FA_X1 \mult_19/S2_21_20  ( .A(\mult_19/ab[21][20] ), .B(
        \mult_19/CARRYB[20][20] ), .CI(\mult_19/SUMB[20][21] ), .CO(
        \mult_19/CARRYB[21][20] ), .S(\mult_19/SUMB[21][20] ) );
  FA_X1 \mult_19/S2_21_19  ( .A(\mult_19/ab[21][19] ), .B(
        \mult_19/CARRYB[20][19] ), .CI(\mult_19/SUMB[20][20] ), .CO(
        \mult_19/CARRYB[21][19] ), .S(\mult_19/SUMB[21][19] ) );
  FA_X1 \mult_19/S2_21_18  ( .A(\mult_19/ab[21][18] ), .B(
        \mult_19/CARRYB[20][18] ), .CI(\mult_19/SUMB[20][19] ), .CO(
        \mult_19/CARRYB[21][18] ), .S(\mult_19/SUMB[21][18] ) );
  FA_X1 \mult_19/S2_21_17  ( .A(\mult_19/ab[21][17] ), .B(
        \mult_19/CARRYB[20][17] ), .CI(\mult_19/SUMB[20][18] ), .CO(
        \mult_19/CARRYB[21][17] ), .S(\mult_19/SUMB[21][17] ) );
  FA_X1 \mult_19/S2_21_16  ( .A(\mult_19/ab[21][16] ), .B(
        \mult_19/CARRYB[20][16] ), .CI(\mult_19/SUMB[20][17] ), .CO(
        \mult_19/CARRYB[21][16] ), .S(\mult_19/SUMB[21][16] ) );
  FA_X1 \mult_19/S2_21_15  ( .A(\mult_19/ab[21][15] ), .B(
        \mult_19/CARRYB[20][15] ), .CI(\mult_19/SUMB[20][16] ), .CO(
        \mult_19/CARRYB[21][15] ), .S(\mult_19/SUMB[21][15] ) );
  FA_X1 \mult_19/S2_21_14  ( .A(\mult_19/ab[21][14] ), .B(
        \mult_19/CARRYB[20][14] ), .CI(\mult_19/SUMB[20][15] ), .CO(
        \mult_19/CARRYB[21][14] ), .S(\mult_19/SUMB[21][14] ) );
  FA_X1 \mult_19/S2_21_13  ( .A(\mult_19/ab[21][13] ), .B(
        \mult_19/CARRYB[20][13] ), .CI(\mult_19/SUMB[20][14] ), .CO(
        \mult_19/CARRYB[21][13] ), .S(\mult_19/SUMB[21][13] ) );
  FA_X1 \mult_19/S2_21_12  ( .A(\mult_19/ab[21][12] ), .B(
        \mult_19/CARRYB[20][12] ), .CI(\mult_19/SUMB[20][13] ), .CO(
        \mult_19/CARRYB[21][12] ), .S(\mult_19/SUMB[21][12] ) );
  FA_X1 \mult_19/S2_21_11  ( .A(\mult_19/ab[21][11] ), .B(
        \mult_19/CARRYB[20][11] ), .CI(\mult_19/SUMB[20][12] ), .CO(
        \mult_19/CARRYB[21][11] ), .S(\mult_19/SUMB[21][11] ) );
  FA_X1 \mult_19/S2_21_10  ( .A(\mult_19/ab[21][10] ), .B(
        \mult_19/CARRYB[20][10] ), .CI(\mult_19/SUMB[20][11] ), .CO(
        \mult_19/CARRYB[21][10] ), .S(\mult_19/SUMB[21][10] ) );
  FA_X1 \mult_19/S2_21_9  ( .A(\mult_19/ab[21][9] ), .B(
        \mult_19/CARRYB[20][9] ), .CI(\mult_19/SUMB[20][10] ), .CO(
        \mult_19/CARRYB[21][9] ), .S(\mult_19/SUMB[21][9] ) );
  FA_X1 \mult_19/S2_21_8  ( .A(\mult_19/ab[21][8] ), .B(
        \mult_19/CARRYB[20][8] ), .CI(\mult_19/SUMB[20][9] ), .CO(
        \mult_19/CARRYB[21][8] ), .S(\mult_19/SUMB[21][8] ) );
  FA_X1 \mult_19/S2_21_7  ( .A(\mult_19/ab[21][7] ), .B(
        \mult_19/CARRYB[20][7] ), .CI(\mult_19/SUMB[20][8] ), .CO(
        \mult_19/CARRYB[21][7] ), .S(\mult_19/SUMB[21][7] ) );
  FA_X1 \mult_19/S2_21_6  ( .A(\mult_19/ab[21][6] ), .B(
        \mult_19/CARRYB[20][6] ), .CI(\mult_19/SUMB[20][7] ), .CO(
        \mult_19/CARRYB[21][6] ), .S(\mult_19/SUMB[21][6] ) );
  FA_X1 \mult_19/S2_21_5  ( .A(\mult_19/ab[21][5] ), .B(
        \mult_19/CARRYB[20][5] ), .CI(\mult_19/SUMB[20][6] ), .CO(
        \mult_19/CARRYB[21][5] ), .S(\mult_19/SUMB[21][5] ) );
  FA_X1 \mult_19/S2_21_4  ( .A(\mult_19/ab[21][4] ), .B(
        \mult_19/CARRYB[20][4] ), .CI(\mult_19/SUMB[20][5] ), .CO(
        \mult_19/CARRYB[21][4] ), .S(\mult_19/SUMB[21][4] ) );
  FA_X1 \mult_19/S2_21_3  ( .A(\mult_19/ab[21][3] ), .B(
        \mult_19/CARRYB[20][3] ), .CI(\mult_19/SUMB[20][4] ), .CO(
        \mult_19/CARRYB[21][3] ), .S(\mult_19/SUMB[21][3] ) );
  FA_X1 \mult_19/S2_21_2  ( .A(\mult_19/ab[21][2] ), .B(
        \mult_19/CARRYB[20][2] ), .CI(\mult_19/SUMB[20][3] ), .CO(
        \mult_19/CARRYB[21][2] ), .S(\mult_19/SUMB[21][2] ) );
  FA_X1 \mult_19/S2_21_1  ( .A(\mult_19/ab[21][1] ), .B(
        \mult_19/CARRYB[20][1] ), .CI(\mult_19/SUMB[20][2] ), .CO(
        \mult_19/CARRYB[21][1] ), .S(\mult_19/SUMB[21][1] ) );
  FA_X1 \mult_19/S1_21_0  ( .A(\mult_19/ab[21][0] ), .B(
        \mult_19/CARRYB[20][0] ), .CI(\mult_19/SUMB[20][1] ), .CO(
        \mult_19/CARRYB[21][0] ), .S(N21) );
  FA_X1 \mult_19/S3_22_30  ( .A(\mult_19/ab[22][30] ), .B(
        \mult_19/CARRYB[21][30] ), .CI(\mult_19/ab[21][31] ), .CO(
        \mult_19/CARRYB[22][30] ), .S(\mult_19/SUMB[22][30] ) );
  FA_X1 \mult_19/S2_22_29  ( .A(\mult_19/ab[22][29] ), .B(
        \mult_19/CARRYB[21][29] ), .CI(\mult_19/SUMB[21][30] ), .CO(
        \mult_19/CARRYB[22][29] ), .S(\mult_19/SUMB[22][29] ) );
  FA_X1 \mult_19/S2_22_28  ( .A(\mult_19/ab[22][28] ), .B(
        \mult_19/CARRYB[21][28] ), .CI(\mult_19/SUMB[21][29] ), .CO(
        \mult_19/CARRYB[22][28] ), .S(\mult_19/SUMB[22][28] ) );
  FA_X1 \mult_19/S2_22_27  ( .A(\mult_19/ab[22][27] ), .B(
        \mult_19/CARRYB[21][27] ), .CI(\mult_19/SUMB[21][28] ), .CO(
        \mult_19/CARRYB[22][27] ), .S(\mult_19/SUMB[22][27] ) );
  FA_X1 \mult_19/S2_22_26  ( .A(\mult_19/ab[22][26] ), .B(
        \mult_19/CARRYB[21][26] ), .CI(\mult_19/SUMB[21][27] ), .CO(
        \mult_19/CARRYB[22][26] ), .S(\mult_19/SUMB[22][26] ) );
  FA_X1 \mult_19/S2_22_25  ( .A(\mult_19/ab[22][25] ), .B(
        \mult_19/CARRYB[21][25] ), .CI(\mult_19/SUMB[21][26] ), .CO(
        \mult_19/CARRYB[22][25] ), .S(\mult_19/SUMB[22][25] ) );
  FA_X1 \mult_19/S2_22_24  ( .A(\mult_19/ab[22][24] ), .B(
        \mult_19/CARRYB[21][24] ), .CI(\mult_19/SUMB[21][25] ), .CO(
        \mult_19/CARRYB[22][24] ), .S(\mult_19/SUMB[22][24] ) );
  FA_X1 \mult_19/S2_22_23  ( .A(\mult_19/ab[22][23] ), .B(
        \mult_19/CARRYB[21][23] ), .CI(\mult_19/SUMB[21][24] ), .CO(
        \mult_19/CARRYB[22][23] ), .S(\mult_19/SUMB[22][23] ) );
  FA_X1 \mult_19/S2_22_22  ( .A(\mult_19/ab[22][22] ), .B(
        \mult_19/CARRYB[21][22] ), .CI(\mult_19/SUMB[21][23] ), .CO(
        \mult_19/CARRYB[22][22] ), .S(\mult_19/SUMB[22][22] ) );
  FA_X1 \mult_19/S2_22_21  ( .A(\mult_19/ab[22][21] ), .B(
        \mult_19/CARRYB[21][21] ), .CI(\mult_19/SUMB[21][22] ), .CO(
        \mult_19/CARRYB[22][21] ), .S(\mult_19/SUMB[22][21] ) );
  FA_X1 \mult_19/S2_22_20  ( .A(\mult_19/ab[22][20] ), .B(
        \mult_19/CARRYB[21][20] ), .CI(\mult_19/SUMB[21][21] ), .CO(
        \mult_19/CARRYB[22][20] ), .S(\mult_19/SUMB[22][20] ) );
  FA_X1 \mult_19/S2_22_19  ( .A(\mult_19/ab[22][19] ), .B(
        \mult_19/CARRYB[21][19] ), .CI(\mult_19/SUMB[21][20] ), .CO(
        \mult_19/CARRYB[22][19] ), .S(\mult_19/SUMB[22][19] ) );
  FA_X1 \mult_19/S2_22_18  ( .A(\mult_19/ab[22][18] ), .B(
        \mult_19/CARRYB[21][18] ), .CI(\mult_19/SUMB[21][19] ), .CO(
        \mult_19/CARRYB[22][18] ), .S(\mult_19/SUMB[22][18] ) );
  FA_X1 \mult_19/S2_22_17  ( .A(\mult_19/ab[22][17] ), .B(
        \mult_19/CARRYB[21][17] ), .CI(\mult_19/SUMB[21][18] ), .CO(
        \mult_19/CARRYB[22][17] ), .S(\mult_19/SUMB[22][17] ) );
  FA_X1 \mult_19/S2_22_16  ( .A(\mult_19/ab[22][16] ), .B(
        \mult_19/CARRYB[21][16] ), .CI(\mult_19/SUMB[21][17] ), .CO(
        \mult_19/CARRYB[22][16] ), .S(\mult_19/SUMB[22][16] ) );
  FA_X1 \mult_19/S2_22_15  ( .A(\mult_19/ab[22][15] ), .B(
        \mult_19/CARRYB[21][15] ), .CI(\mult_19/SUMB[21][16] ), .CO(
        \mult_19/CARRYB[22][15] ), .S(\mult_19/SUMB[22][15] ) );
  FA_X1 \mult_19/S2_22_14  ( .A(\mult_19/ab[22][14] ), .B(
        \mult_19/CARRYB[21][14] ), .CI(\mult_19/SUMB[21][15] ), .CO(
        \mult_19/CARRYB[22][14] ), .S(\mult_19/SUMB[22][14] ) );
  FA_X1 \mult_19/S2_22_13  ( .A(\mult_19/ab[22][13] ), .B(
        \mult_19/CARRYB[21][13] ), .CI(\mult_19/SUMB[21][14] ), .CO(
        \mult_19/CARRYB[22][13] ), .S(\mult_19/SUMB[22][13] ) );
  FA_X1 \mult_19/S2_22_12  ( .A(\mult_19/ab[22][12] ), .B(
        \mult_19/CARRYB[21][12] ), .CI(\mult_19/SUMB[21][13] ), .CO(
        \mult_19/CARRYB[22][12] ), .S(\mult_19/SUMB[22][12] ) );
  FA_X1 \mult_19/S2_22_11  ( .A(\mult_19/ab[22][11] ), .B(
        \mult_19/CARRYB[21][11] ), .CI(\mult_19/SUMB[21][12] ), .CO(
        \mult_19/CARRYB[22][11] ), .S(\mult_19/SUMB[22][11] ) );
  FA_X1 \mult_19/S2_22_10  ( .A(\mult_19/ab[22][10] ), .B(
        \mult_19/CARRYB[21][10] ), .CI(\mult_19/SUMB[21][11] ), .CO(
        \mult_19/CARRYB[22][10] ), .S(\mult_19/SUMB[22][10] ) );
  FA_X1 \mult_19/S2_22_9  ( .A(\mult_19/ab[22][9] ), .B(
        \mult_19/CARRYB[21][9] ), .CI(\mult_19/SUMB[21][10] ), .CO(
        \mult_19/CARRYB[22][9] ), .S(\mult_19/SUMB[22][9] ) );
  FA_X1 \mult_19/S2_22_8  ( .A(\mult_19/ab[22][8] ), .B(
        \mult_19/CARRYB[21][8] ), .CI(\mult_19/SUMB[21][9] ), .CO(
        \mult_19/CARRYB[22][8] ), .S(\mult_19/SUMB[22][8] ) );
  FA_X1 \mult_19/S2_22_7  ( .A(\mult_19/ab[22][7] ), .B(
        \mult_19/CARRYB[21][7] ), .CI(\mult_19/SUMB[21][8] ), .CO(
        \mult_19/CARRYB[22][7] ), .S(\mult_19/SUMB[22][7] ) );
  FA_X1 \mult_19/S2_22_6  ( .A(\mult_19/ab[22][6] ), .B(
        \mult_19/CARRYB[21][6] ), .CI(\mult_19/SUMB[21][7] ), .CO(
        \mult_19/CARRYB[22][6] ), .S(\mult_19/SUMB[22][6] ) );
  FA_X1 \mult_19/S2_22_5  ( .A(\mult_19/ab[22][5] ), .B(
        \mult_19/CARRYB[21][5] ), .CI(\mult_19/SUMB[21][6] ), .CO(
        \mult_19/CARRYB[22][5] ), .S(\mult_19/SUMB[22][5] ) );
  FA_X1 \mult_19/S2_22_4  ( .A(\mult_19/ab[22][4] ), .B(
        \mult_19/CARRYB[21][4] ), .CI(\mult_19/SUMB[21][5] ), .CO(
        \mult_19/CARRYB[22][4] ), .S(\mult_19/SUMB[22][4] ) );
  FA_X1 \mult_19/S2_22_3  ( .A(\mult_19/ab[22][3] ), .B(
        \mult_19/CARRYB[21][3] ), .CI(\mult_19/SUMB[21][4] ), .CO(
        \mult_19/CARRYB[22][3] ), .S(\mult_19/SUMB[22][3] ) );
  FA_X1 \mult_19/S2_22_2  ( .A(\mult_19/ab[22][2] ), .B(
        \mult_19/CARRYB[21][2] ), .CI(\mult_19/SUMB[21][3] ), .CO(
        \mult_19/CARRYB[22][2] ), .S(\mult_19/SUMB[22][2] ) );
  FA_X1 \mult_19/S2_22_1  ( .A(\mult_19/ab[22][1] ), .B(
        \mult_19/CARRYB[21][1] ), .CI(\mult_19/SUMB[21][2] ), .CO(
        \mult_19/CARRYB[22][1] ), .S(\mult_19/SUMB[22][1] ) );
  FA_X1 \mult_19/S1_22_0  ( .A(\mult_19/ab[22][0] ), .B(
        \mult_19/CARRYB[21][0] ), .CI(\mult_19/SUMB[21][1] ), .CO(
        \mult_19/CARRYB[22][0] ), .S(N22) );
  FA_X1 \mult_19/S3_23_30  ( .A(\mult_19/ab[23][30] ), .B(
        \mult_19/CARRYB[22][30] ), .CI(\mult_19/ab[22][31] ), .CO(
        \mult_19/CARRYB[23][30] ), .S(\mult_19/SUMB[23][30] ) );
  FA_X1 \mult_19/S2_23_29  ( .A(\mult_19/ab[23][29] ), .B(
        \mult_19/CARRYB[22][29] ), .CI(\mult_19/SUMB[22][30] ), .CO(
        \mult_19/CARRYB[23][29] ), .S(\mult_19/SUMB[23][29] ) );
  FA_X1 \mult_19/S2_23_28  ( .A(\mult_19/ab[23][28] ), .B(
        \mult_19/CARRYB[22][28] ), .CI(\mult_19/SUMB[22][29] ), .CO(
        \mult_19/CARRYB[23][28] ), .S(\mult_19/SUMB[23][28] ) );
  FA_X1 \mult_19/S2_23_27  ( .A(\mult_19/ab[23][27] ), .B(
        \mult_19/CARRYB[22][27] ), .CI(\mult_19/SUMB[22][28] ), .CO(
        \mult_19/CARRYB[23][27] ), .S(\mult_19/SUMB[23][27] ) );
  FA_X1 \mult_19/S2_23_26  ( .A(\mult_19/ab[23][26] ), .B(
        \mult_19/CARRYB[22][26] ), .CI(\mult_19/SUMB[22][27] ), .CO(
        \mult_19/CARRYB[23][26] ), .S(\mult_19/SUMB[23][26] ) );
  FA_X1 \mult_19/S2_23_25  ( .A(\mult_19/ab[23][25] ), .B(
        \mult_19/CARRYB[22][25] ), .CI(\mult_19/SUMB[22][26] ), .CO(
        \mult_19/CARRYB[23][25] ), .S(\mult_19/SUMB[23][25] ) );
  FA_X1 \mult_19/S2_23_24  ( .A(\mult_19/ab[23][24] ), .B(
        \mult_19/CARRYB[22][24] ), .CI(\mult_19/SUMB[22][25] ), .CO(
        \mult_19/CARRYB[23][24] ), .S(\mult_19/SUMB[23][24] ) );
  FA_X1 \mult_19/S2_23_23  ( .A(\mult_19/ab[23][23] ), .B(
        \mult_19/CARRYB[22][23] ), .CI(\mult_19/SUMB[22][24] ), .CO(
        \mult_19/CARRYB[23][23] ), .S(\mult_19/SUMB[23][23] ) );
  FA_X1 \mult_19/S2_23_22  ( .A(\mult_19/ab[23][22] ), .B(
        \mult_19/CARRYB[22][22] ), .CI(\mult_19/SUMB[22][23] ), .CO(
        \mult_19/CARRYB[23][22] ), .S(\mult_19/SUMB[23][22] ) );
  FA_X1 \mult_19/S2_23_21  ( .A(\mult_19/ab[23][21] ), .B(
        \mult_19/CARRYB[22][21] ), .CI(\mult_19/SUMB[22][22] ), .CO(
        \mult_19/CARRYB[23][21] ), .S(\mult_19/SUMB[23][21] ) );
  FA_X1 \mult_19/S2_23_20  ( .A(\mult_19/ab[23][20] ), .B(
        \mult_19/CARRYB[22][20] ), .CI(\mult_19/SUMB[22][21] ), .CO(
        \mult_19/CARRYB[23][20] ), .S(\mult_19/SUMB[23][20] ) );
  FA_X1 \mult_19/S2_23_19  ( .A(\mult_19/ab[23][19] ), .B(
        \mult_19/CARRYB[22][19] ), .CI(\mult_19/SUMB[22][20] ), .CO(
        \mult_19/CARRYB[23][19] ), .S(\mult_19/SUMB[23][19] ) );
  FA_X1 \mult_19/S2_23_18  ( .A(\mult_19/ab[23][18] ), .B(
        \mult_19/CARRYB[22][18] ), .CI(\mult_19/SUMB[22][19] ), .CO(
        \mult_19/CARRYB[23][18] ), .S(\mult_19/SUMB[23][18] ) );
  FA_X1 \mult_19/S2_23_17  ( .A(\mult_19/ab[23][17] ), .B(
        \mult_19/CARRYB[22][17] ), .CI(\mult_19/SUMB[22][18] ), .CO(
        \mult_19/CARRYB[23][17] ), .S(\mult_19/SUMB[23][17] ) );
  FA_X1 \mult_19/S2_23_16  ( .A(\mult_19/ab[23][16] ), .B(
        \mult_19/CARRYB[22][16] ), .CI(\mult_19/SUMB[22][17] ), .CO(
        \mult_19/CARRYB[23][16] ), .S(\mult_19/SUMB[23][16] ) );
  FA_X1 \mult_19/S2_23_15  ( .A(\mult_19/ab[23][15] ), .B(
        \mult_19/CARRYB[22][15] ), .CI(\mult_19/SUMB[22][16] ), .CO(
        \mult_19/CARRYB[23][15] ), .S(\mult_19/SUMB[23][15] ) );
  FA_X1 \mult_19/S2_23_14  ( .A(\mult_19/ab[23][14] ), .B(
        \mult_19/CARRYB[22][14] ), .CI(\mult_19/SUMB[22][15] ), .CO(
        \mult_19/CARRYB[23][14] ), .S(\mult_19/SUMB[23][14] ) );
  FA_X1 \mult_19/S2_23_13  ( .A(\mult_19/ab[23][13] ), .B(
        \mult_19/CARRYB[22][13] ), .CI(\mult_19/SUMB[22][14] ), .CO(
        \mult_19/CARRYB[23][13] ), .S(\mult_19/SUMB[23][13] ) );
  FA_X1 \mult_19/S2_23_12  ( .A(\mult_19/ab[23][12] ), .B(
        \mult_19/CARRYB[22][12] ), .CI(\mult_19/SUMB[22][13] ), .CO(
        \mult_19/CARRYB[23][12] ), .S(\mult_19/SUMB[23][12] ) );
  FA_X1 \mult_19/S2_23_11  ( .A(\mult_19/ab[23][11] ), .B(
        \mult_19/CARRYB[22][11] ), .CI(\mult_19/SUMB[22][12] ), .CO(
        \mult_19/CARRYB[23][11] ), .S(\mult_19/SUMB[23][11] ) );
  FA_X1 \mult_19/S2_23_10  ( .A(\mult_19/ab[23][10] ), .B(
        \mult_19/CARRYB[22][10] ), .CI(\mult_19/SUMB[22][11] ), .CO(
        \mult_19/CARRYB[23][10] ), .S(\mult_19/SUMB[23][10] ) );
  FA_X1 \mult_19/S2_23_9  ( .A(\mult_19/ab[23][9] ), .B(
        \mult_19/CARRYB[22][9] ), .CI(\mult_19/SUMB[22][10] ), .CO(
        \mult_19/CARRYB[23][9] ), .S(\mult_19/SUMB[23][9] ) );
  FA_X1 \mult_19/S2_23_8  ( .A(\mult_19/ab[23][8] ), .B(
        \mult_19/CARRYB[22][8] ), .CI(\mult_19/SUMB[22][9] ), .CO(
        \mult_19/CARRYB[23][8] ), .S(\mult_19/SUMB[23][8] ) );
  FA_X1 \mult_19/S2_23_7  ( .A(\mult_19/ab[23][7] ), .B(
        \mult_19/CARRYB[22][7] ), .CI(\mult_19/SUMB[22][8] ), .CO(
        \mult_19/CARRYB[23][7] ), .S(\mult_19/SUMB[23][7] ) );
  FA_X1 \mult_19/S2_23_6  ( .A(\mult_19/ab[23][6] ), .B(
        \mult_19/CARRYB[22][6] ), .CI(\mult_19/SUMB[22][7] ), .CO(
        \mult_19/CARRYB[23][6] ), .S(\mult_19/SUMB[23][6] ) );
  FA_X1 \mult_19/S2_23_5  ( .A(\mult_19/ab[23][5] ), .B(
        \mult_19/CARRYB[22][5] ), .CI(\mult_19/SUMB[22][6] ), .CO(
        \mult_19/CARRYB[23][5] ), .S(\mult_19/SUMB[23][5] ) );
  FA_X1 \mult_19/S2_23_4  ( .A(\mult_19/ab[23][4] ), .B(
        \mult_19/CARRYB[22][4] ), .CI(\mult_19/SUMB[22][5] ), .CO(
        \mult_19/CARRYB[23][4] ), .S(\mult_19/SUMB[23][4] ) );
  FA_X1 \mult_19/S2_23_3  ( .A(\mult_19/ab[23][3] ), .B(
        \mult_19/CARRYB[22][3] ), .CI(\mult_19/SUMB[22][4] ), .CO(
        \mult_19/CARRYB[23][3] ), .S(\mult_19/SUMB[23][3] ) );
  FA_X1 \mult_19/S2_23_2  ( .A(\mult_19/ab[23][2] ), .B(
        \mult_19/CARRYB[22][2] ), .CI(\mult_19/SUMB[22][3] ), .CO(
        \mult_19/CARRYB[23][2] ), .S(\mult_19/SUMB[23][2] ) );
  FA_X1 \mult_19/S2_23_1  ( .A(\mult_19/ab[23][1] ), .B(
        \mult_19/CARRYB[22][1] ), .CI(\mult_19/SUMB[22][2] ), .CO(
        \mult_19/CARRYB[23][1] ), .S(\mult_19/SUMB[23][1] ) );
  FA_X1 \mult_19/S1_23_0  ( .A(\mult_19/ab[23][0] ), .B(
        \mult_19/CARRYB[22][0] ), .CI(\mult_19/SUMB[22][1] ), .CO(
        \mult_19/CARRYB[23][0] ), .S(N23) );
  FA_X1 \mult_19/S3_24_30  ( .A(\mult_19/ab[24][30] ), .B(
        \mult_19/CARRYB[23][30] ), .CI(\mult_19/ab[23][31] ), .CO(
        \mult_19/CARRYB[24][30] ), .S(\mult_19/SUMB[24][30] ) );
  FA_X1 \mult_19/S2_24_29  ( .A(\mult_19/ab[24][29] ), .B(
        \mult_19/CARRYB[23][29] ), .CI(\mult_19/SUMB[23][30] ), .CO(
        \mult_19/CARRYB[24][29] ), .S(\mult_19/SUMB[24][29] ) );
  FA_X1 \mult_19/S2_24_28  ( .A(\mult_19/ab[24][28] ), .B(
        \mult_19/CARRYB[23][28] ), .CI(\mult_19/SUMB[23][29] ), .CO(
        \mult_19/CARRYB[24][28] ), .S(\mult_19/SUMB[24][28] ) );
  FA_X1 \mult_19/S2_24_27  ( .A(\mult_19/ab[24][27] ), .B(
        \mult_19/CARRYB[23][27] ), .CI(\mult_19/SUMB[23][28] ), .CO(
        \mult_19/CARRYB[24][27] ), .S(\mult_19/SUMB[24][27] ) );
  FA_X1 \mult_19/S2_24_26  ( .A(\mult_19/ab[24][26] ), .B(
        \mult_19/CARRYB[23][26] ), .CI(\mult_19/SUMB[23][27] ), .CO(
        \mult_19/CARRYB[24][26] ), .S(\mult_19/SUMB[24][26] ) );
  FA_X1 \mult_19/S2_24_25  ( .A(\mult_19/ab[24][25] ), .B(
        \mult_19/CARRYB[23][25] ), .CI(\mult_19/SUMB[23][26] ), .CO(
        \mult_19/CARRYB[24][25] ), .S(\mult_19/SUMB[24][25] ) );
  FA_X1 \mult_19/S2_24_24  ( .A(\mult_19/ab[24][24] ), .B(
        \mult_19/CARRYB[23][24] ), .CI(\mult_19/SUMB[23][25] ), .CO(
        \mult_19/CARRYB[24][24] ), .S(\mult_19/SUMB[24][24] ) );
  FA_X1 \mult_19/S2_24_23  ( .A(\mult_19/ab[24][23] ), .B(
        \mult_19/CARRYB[23][23] ), .CI(\mult_19/SUMB[23][24] ), .CO(
        \mult_19/CARRYB[24][23] ), .S(\mult_19/SUMB[24][23] ) );
  FA_X1 \mult_19/S2_24_22  ( .A(\mult_19/ab[24][22] ), .B(
        \mult_19/CARRYB[23][22] ), .CI(\mult_19/SUMB[23][23] ), .CO(
        \mult_19/CARRYB[24][22] ), .S(\mult_19/SUMB[24][22] ) );
  FA_X1 \mult_19/S2_24_21  ( .A(\mult_19/ab[24][21] ), .B(
        \mult_19/CARRYB[23][21] ), .CI(\mult_19/SUMB[23][22] ), .CO(
        \mult_19/CARRYB[24][21] ), .S(\mult_19/SUMB[24][21] ) );
  FA_X1 \mult_19/S2_24_20  ( .A(\mult_19/ab[24][20] ), .B(
        \mult_19/CARRYB[23][20] ), .CI(\mult_19/SUMB[23][21] ), .CO(
        \mult_19/CARRYB[24][20] ), .S(\mult_19/SUMB[24][20] ) );
  FA_X1 \mult_19/S2_24_19  ( .A(\mult_19/ab[24][19] ), .B(
        \mult_19/CARRYB[23][19] ), .CI(\mult_19/SUMB[23][20] ), .CO(
        \mult_19/CARRYB[24][19] ), .S(\mult_19/SUMB[24][19] ) );
  FA_X1 \mult_19/S2_24_18  ( .A(\mult_19/ab[24][18] ), .B(
        \mult_19/CARRYB[23][18] ), .CI(\mult_19/SUMB[23][19] ), .CO(
        \mult_19/CARRYB[24][18] ), .S(\mult_19/SUMB[24][18] ) );
  FA_X1 \mult_19/S2_24_17  ( .A(\mult_19/ab[24][17] ), .B(
        \mult_19/CARRYB[23][17] ), .CI(\mult_19/SUMB[23][18] ), .CO(
        \mult_19/CARRYB[24][17] ), .S(\mult_19/SUMB[24][17] ) );
  FA_X1 \mult_19/S2_24_16  ( .A(\mult_19/ab[24][16] ), .B(
        \mult_19/CARRYB[23][16] ), .CI(\mult_19/SUMB[23][17] ), .CO(
        \mult_19/CARRYB[24][16] ), .S(\mult_19/SUMB[24][16] ) );
  FA_X1 \mult_19/S2_24_15  ( .A(\mult_19/ab[24][15] ), .B(
        \mult_19/CARRYB[23][15] ), .CI(\mult_19/SUMB[23][16] ), .CO(
        \mult_19/CARRYB[24][15] ), .S(\mult_19/SUMB[24][15] ) );
  FA_X1 \mult_19/S2_24_14  ( .A(\mult_19/ab[24][14] ), .B(
        \mult_19/CARRYB[23][14] ), .CI(\mult_19/SUMB[23][15] ), .CO(
        \mult_19/CARRYB[24][14] ), .S(\mult_19/SUMB[24][14] ) );
  FA_X1 \mult_19/S2_24_13  ( .A(\mult_19/ab[24][13] ), .B(
        \mult_19/CARRYB[23][13] ), .CI(\mult_19/SUMB[23][14] ), .CO(
        \mult_19/CARRYB[24][13] ), .S(\mult_19/SUMB[24][13] ) );
  FA_X1 \mult_19/S2_24_12  ( .A(\mult_19/ab[24][12] ), .B(
        \mult_19/CARRYB[23][12] ), .CI(\mult_19/SUMB[23][13] ), .CO(
        \mult_19/CARRYB[24][12] ), .S(\mult_19/SUMB[24][12] ) );
  FA_X1 \mult_19/S2_24_11  ( .A(\mult_19/ab[24][11] ), .B(
        \mult_19/CARRYB[23][11] ), .CI(\mult_19/SUMB[23][12] ), .CO(
        \mult_19/CARRYB[24][11] ), .S(\mult_19/SUMB[24][11] ) );
  FA_X1 \mult_19/S2_24_10  ( .A(\mult_19/ab[24][10] ), .B(
        \mult_19/CARRYB[23][10] ), .CI(\mult_19/SUMB[23][11] ), .CO(
        \mult_19/CARRYB[24][10] ), .S(\mult_19/SUMB[24][10] ) );
  FA_X1 \mult_19/S2_24_9  ( .A(\mult_19/ab[24][9] ), .B(
        \mult_19/CARRYB[23][9] ), .CI(\mult_19/SUMB[23][10] ), .CO(
        \mult_19/CARRYB[24][9] ), .S(\mult_19/SUMB[24][9] ) );
  FA_X1 \mult_19/S2_24_8  ( .A(\mult_19/ab[24][8] ), .B(
        \mult_19/CARRYB[23][8] ), .CI(\mult_19/SUMB[23][9] ), .CO(
        \mult_19/CARRYB[24][8] ), .S(\mult_19/SUMB[24][8] ) );
  FA_X1 \mult_19/S2_24_7  ( .A(\mult_19/ab[24][7] ), .B(
        \mult_19/CARRYB[23][7] ), .CI(\mult_19/SUMB[23][8] ), .CO(
        \mult_19/CARRYB[24][7] ), .S(\mult_19/SUMB[24][7] ) );
  FA_X1 \mult_19/S2_24_6  ( .A(\mult_19/ab[24][6] ), .B(
        \mult_19/CARRYB[23][6] ), .CI(\mult_19/SUMB[23][7] ), .CO(
        \mult_19/CARRYB[24][6] ), .S(\mult_19/SUMB[24][6] ) );
  FA_X1 \mult_19/S2_24_5  ( .A(\mult_19/ab[24][5] ), .B(
        \mult_19/CARRYB[23][5] ), .CI(\mult_19/SUMB[23][6] ), .CO(
        \mult_19/CARRYB[24][5] ), .S(\mult_19/SUMB[24][5] ) );
  FA_X1 \mult_19/S2_24_4  ( .A(\mult_19/ab[24][4] ), .B(
        \mult_19/CARRYB[23][4] ), .CI(\mult_19/SUMB[23][5] ), .CO(
        \mult_19/CARRYB[24][4] ), .S(\mult_19/SUMB[24][4] ) );
  FA_X1 \mult_19/S2_24_3  ( .A(\mult_19/ab[24][3] ), .B(
        \mult_19/CARRYB[23][3] ), .CI(\mult_19/SUMB[23][4] ), .CO(
        \mult_19/CARRYB[24][3] ), .S(\mult_19/SUMB[24][3] ) );
  FA_X1 \mult_19/S2_24_2  ( .A(\mult_19/ab[24][2] ), .B(
        \mult_19/CARRYB[23][2] ), .CI(\mult_19/SUMB[23][3] ), .CO(
        \mult_19/CARRYB[24][2] ), .S(\mult_19/SUMB[24][2] ) );
  FA_X1 \mult_19/S2_24_1  ( .A(\mult_19/ab[24][1] ), .B(
        \mult_19/CARRYB[23][1] ), .CI(\mult_19/SUMB[23][2] ), .CO(
        \mult_19/CARRYB[24][1] ), .S(\mult_19/SUMB[24][1] ) );
  FA_X1 \mult_19/S1_24_0  ( .A(\mult_19/ab[24][0] ), .B(
        \mult_19/CARRYB[23][0] ), .CI(\mult_19/SUMB[23][1] ), .CO(
        \mult_19/CARRYB[24][0] ), .S(N24) );
  FA_X1 \mult_19/S3_25_30  ( .A(\mult_19/ab[25][30] ), .B(
        \mult_19/CARRYB[24][30] ), .CI(\mult_19/ab[24][31] ), .CO(
        \mult_19/CARRYB[25][30] ), .S(\mult_19/SUMB[25][30] ) );
  FA_X1 \mult_19/S2_25_29  ( .A(\mult_19/ab[25][29] ), .B(
        \mult_19/CARRYB[24][29] ), .CI(\mult_19/SUMB[24][30] ), .CO(
        \mult_19/CARRYB[25][29] ), .S(\mult_19/SUMB[25][29] ) );
  FA_X1 \mult_19/S2_25_28  ( .A(\mult_19/ab[25][28] ), .B(
        \mult_19/CARRYB[24][28] ), .CI(\mult_19/SUMB[24][29] ), .CO(
        \mult_19/CARRYB[25][28] ), .S(\mult_19/SUMB[25][28] ) );
  FA_X1 \mult_19/S2_25_27  ( .A(\mult_19/ab[25][27] ), .B(
        \mult_19/CARRYB[24][27] ), .CI(\mult_19/SUMB[24][28] ), .CO(
        \mult_19/CARRYB[25][27] ), .S(\mult_19/SUMB[25][27] ) );
  FA_X1 \mult_19/S2_25_26  ( .A(\mult_19/ab[25][26] ), .B(
        \mult_19/CARRYB[24][26] ), .CI(\mult_19/SUMB[24][27] ), .CO(
        \mult_19/CARRYB[25][26] ), .S(\mult_19/SUMB[25][26] ) );
  FA_X1 \mult_19/S2_25_25  ( .A(\mult_19/ab[25][25] ), .B(
        \mult_19/CARRYB[24][25] ), .CI(\mult_19/SUMB[24][26] ), .CO(
        \mult_19/CARRYB[25][25] ), .S(\mult_19/SUMB[25][25] ) );
  FA_X1 \mult_19/S2_25_24  ( .A(\mult_19/ab[25][24] ), .B(
        \mult_19/CARRYB[24][24] ), .CI(\mult_19/SUMB[24][25] ), .CO(
        \mult_19/CARRYB[25][24] ), .S(\mult_19/SUMB[25][24] ) );
  FA_X1 \mult_19/S2_25_23  ( .A(\mult_19/ab[25][23] ), .B(
        \mult_19/CARRYB[24][23] ), .CI(\mult_19/SUMB[24][24] ), .CO(
        \mult_19/CARRYB[25][23] ), .S(\mult_19/SUMB[25][23] ) );
  FA_X1 \mult_19/S2_25_22  ( .A(\mult_19/ab[25][22] ), .B(
        \mult_19/CARRYB[24][22] ), .CI(\mult_19/SUMB[24][23] ), .CO(
        \mult_19/CARRYB[25][22] ), .S(\mult_19/SUMB[25][22] ) );
  FA_X1 \mult_19/S2_25_21  ( .A(\mult_19/ab[25][21] ), .B(
        \mult_19/CARRYB[24][21] ), .CI(\mult_19/SUMB[24][22] ), .CO(
        \mult_19/CARRYB[25][21] ), .S(\mult_19/SUMB[25][21] ) );
  FA_X1 \mult_19/S2_25_20  ( .A(\mult_19/ab[25][20] ), .B(
        \mult_19/CARRYB[24][20] ), .CI(\mult_19/SUMB[24][21] ), .CO(
        \mult_19/CARRYB[25][20] ), .S(\mult_19/SUMB[25][20] ) );
  FA_X1 \mult_19/S2_25_19  ( .A(\mult_19/ab[25][19] ), .B(
        \mult_19/CARRYB[24][19] ), .CI(\mult_19/SUMB[24][20] ), .CO(
        \mult_19/CARRYB[25][19] ), .S(\mult_19/SUMB[25][19] ) );
  FA_X1 \mult_19/S2_25_18  ( .A(\mult_19/ab[25][18] ), .B(
        \mult_19/CARRYB[24][18] ), .CI(\mult_19/SUMB[24][19] ), .CO(
        \mult_19/CARRYB[25][18] ), .S(\mult_19/SUMB[25][18] ) );
  FA_X1 \mult_19/S2_25_17  ( .A(\mult_19/ab[25][17] ), .B(
        \mult_19/CARRYB[24][17] ), .CI(\mult_19/SUMB[24][18] ), .CO(
        \mult_19/CARRYB[25][17] ), .S(\mult_19/SUMB[25][17] ) );
  FA_X1 \mult_19/S2_25_16  ( .A(\mult_19/ab[25][16] ), .B(
        \mult_19/CARRYB[24][16] ), .CI(\mult_19/SUMB[24][17] ), .CO(
        \mult_19/CARRYB[25][16] ), .S(\mult_19/SUMB[25][16] ) );
  FA_X1 \mult_19/S2_25_15  ( .A(\mult_19/ab[25][15] ), .B(
        \mult_19/CARRYB[24][15] ), .CI(\mult_19/SUMB[24][16] ), .CO(
        \mult_19/CARRYB[25][15] ), .S(\mult_19/SUMB[25][15] ) );
  FA_X1 \mult_19/S2_25_14  ( .A(\mult_19/ab[25][14] ), .B(
        \mult_19/CARRYB[24][14] ), .CI(\mult_19/SUMB[24][15] ), .CO(
        \mult_19/CARRYB[25][14] ), .S(\mult_19/SUMB[25][14] ) );
  FA_X1 \mult_19/S2_25_13  ( .A(\mult_19/ab[25][13] ), .B(
        \mult_19/CARRYB[24][13] ), .CI(\mult_19/SUMB[24][14] ), .CO(
        \mult_19/CARRYB[25][13] ), .S(\mult_19/SUMB[25][13] ) );
  FA_X1 \mult_19/S2_25_12  ( .A(\mult_19/ab[25][12] ), .B(
        \mult_19/CARRYB[24][12] ), .CI(\mult_19/SUMB[24][13] ), .CO(
        \mult_19/CARRYB[25][12] ), .S(\mult_19/SUMB[25][12] ) );
  FA_X1 \mult_19/S2_25_11  ( .A(\mult_19/ab[25][11] ), .B(
        \mult_19/CARRYB[24][11] ), .CI(\mult_19/SUMB[24][12] ), .CO(
        \mult_19/CARRYB[25][11] ), .S(\mult_19/SUMB[25][11] ) );
  FA_X1 \mult_19/S2_25_10  ( .A(\mult_19/ab[25][10] ), .B(
        \mult_19/CARRYB[24][10] ), .CI(\mult_19/SUMB[24][11] ), .CO(
        \mult_19/CARRYB[25][10] ), .S(\mult_19/SUMB[25][10] ) );
  FA_X1 \mult_19/S2_25_9  ( .A(\mult_19/ab[25][9] ), .B(
        \mult_19/CARRYB[24][9] ), .CI(\mult_19/SUMB[24][10] ), .CO(
        \mult_19/CARRYB[25][9] ), .S(\mult_19/SUMB[25][9] ) );
  FA_X1 \mult_19/S2_25_8  ( .A(\mult_19/ab[25][8] ), .B(
        \mult_19/CARRYB[24][8] ), .CI(\mult_19/SUMB[24][9] ), .CO(
        \mult_19/CARRYB[25][8] ), .S(\mult_19/SUMB[25][8] ) );
  FA_X1 \mult_19/S2_25_7  ( .A(\mult_19/ab[25][7] ), .B(
        \mult_19/CARRYB[24][7] ), .CI(\mult_19/SUMB[24][8] ), .CO(
        \mult_19/CARRYB[25][7] ), .S(\mult_19/SUMB[25][7] ) );
  FA_X1 \mult_19/S2_25_6  ( .A(\mult_19/ab[25][6] ), .B(
        \mult_19/CARRYB[24][6] ), .CI(\mult_19/SUMB[24][7] ), .CO(
        \mult_19/CARRYB[25][6] ), .S(\mult_19/SUMB[25][6] ) );
  FA_X1 \mult_19/S2_25_5  ( .A(\mult_19/ab[25][5] ), .B(
        \mult_19/CARRYB[24][5] ), .CI(\mult_19/SUMB[24][6] ), .CO(
        \mult_19/CARRYB[25][5] ), .S(\mult_19/SUMB[25][5] ) );
  FA_X1 \mult_19/S2_25_4  ( .A(\mult_19/ab[25][4] ), .B(
        \mult_19/CARRYB[24][4] ), .CI(\mult_19/SUMB[24][5] ), .CO(
        \mult_19/CARRYB[25][4] ), .S(\mult_19/SUMB[25][4] ) );
  FA_X1 \mult_19/S2_25_3  ( .A(\mult_19/ab[25][3] ), .B(
        \mult_19/CARRYB[24][3] ), .CI(\mult_19/SUMB[24][4] ), .CO(
        \mult_19/CARRYB[25][3] ), .S(\mult_19/SUMB[25][3] ) );
  FA_X1 \mult_19/S2_25_2  ( .A(\mult_19/ab[25][2] ), .B(
        \mult_19/CARRYB[24][2] ), .CI(\mult_19/SUMB[24][3] ), .CO(
        \mult_19/CARRYB[25][2] ), .S(\mult_19/SUMB[25][2] ) );
  FA_X1 \mult_19/S2_25_1  ( .A(\mult_19/ab[25][1] ), .B(
        \mult_19/CARRYB[24][1] ), .CI(\mult_19/SUMB[24][2] ), .CO(
        \mult_19/CARRYB[25][1] ), .S(\mult_19/SUMB[25][1] ) );
  FA_X1 \mult_19/S1_25_0  ( .A(\mult_19/ab[25][0] ), .B(
        \mult_19/CARRYB[24][0] ), .CI(\mult_19/SUMB[24][1] ), .CO(
        \mult_19/CARRYB[25][0] ), .S(N25) );
  FA_X1 \mult_19/S3_26_30  ( .A(\mult_19/ab[26][30] ), .B(
        \mult_19/CARRYB[25][30] ), .CI(\mult_19/ab[25][31] ), .CO(
        \mult_19/CARRYB[26][30] ), .S(\mult_19/SUMB[26][30] ) );
  FA_X1 \mult_19/S2_26_29  ( .A(\mult_19/ab[26][29] ), .B(
        \mult_19/CARRYB[25][29] ), .CI(\mult_19/SUMB[25][30] ), .CO(
        \mult_19/CARRYB[26][29] ), .S(\mult_19/SUMB[26][29] ) );
  FA_X1 \mult_19/S2_26_28  ( .A(\mult_19/ab[26][28] ), .B(
        \mult_19/CARRYB[25][28] ), .CI(\mult_19/SUMB[25][29] ), .CO(
        \mult_19/CARRYB[26][28] ), .S(\mult_19/SUMB[26][28] ) );
  FA_X1 \mult_19/S2_26_27  ( .A(\mult_19/ab[26][27] ), .B(
        \mult_19/CARRYB[25][27] ), .CI(\mult_19/SUMB[25][28] ), .CO(
        \mult_19/CARRYB[26][27] ), .S(\mult_19/SUMB[26][27] ) );
  FA_X1 \mult_19/S2_26_26  ( .A(\mult_19/ab[26][26] ), .B(
        \mult_19/CARRYB[25][26] ), .CI(\mult_19/SUMB[25][27] ), .CO(
        \mult_19/CARRYB[26][26] ), .S(\mult_19/SUMB[26][26] ) );
  FA_X1 \mult_19/S2_26_25  ( .A(\mult_19/ab[26][25] ), .B(
        \mult_19/CARRYB[25][25] ), .CI(\mult_19/SUMB[25][26] ), .CO(
        \mult_19/CARRYB[26][25] ), .S(\mult_19/SUMB[26][25] ) );
  FA_X1 \mult_19/S2_26_24  ( .A(\mult_19/ab[26][24] ), .B(
        \mult_19/CARRYB[25][24] ), .CI(\mult_19/SUMB[25][25] ), .CO(
        \mult_19/CARRYB[26][24] ), .S(\mult_19/SUMB[26][24] ) );
  FA_X1 \mult_19/S2_26_23  ( .A(\mult_19/ab[26][23] ), .B(
        \mult_19/CARRYB[25][23] ), .CI(\mult_19/SUMB[25][24] ), .CO(
        \mult_19/CARRYB[26][23] ), .S(\mult_19/SUMB[26][23] ) );
  FA_X1 \mult_19/S2_26_22  ( .A(\mult_19/ab[26][22] ), .B(
        \mult_19/CARRYB[25][22] ), .CI(\mult_19/SUMB[25][23] ), .CO(
        \mult_19/CARRYB[26][22] ), .S(\mult_19/SUMB[26][22] ) );
  FA_X1 \mult_19/S2_26_21  ( .A(\mult_19/ab[26][21] ), .B(
        \mult_19/CARRYB[25][21] ), .CI(\mult_19/SUMB[25][22] ), .CO(
        \mult_19/CARRYB[26][21] ), .S(\mult_19/SUMB[26][21] ) );
  FA_X1 \mult_19/S2_26_20  ( .A(\mult_19/ab[26][20] ), .B(
        \mult_19/CARRYB[25][20] ), .CI(\mult_19/SUMB[25][21] ), .CO(
        \mult_19/CARRYB[26][20] ), .S(\mult_19/SUMB[26][20] ) );
  FA_X1 \mult_19/S2_26_19  ( .A(\mult_19/ab[26][19] ), .B(
        \mult_19/CARRYB[25][19] ), .CI(\mult_19/SUMB[25][20] ), .CO(
        \mult_19/CARRYB[26][19] ), .S(\mult_19/SUMB[26][19] ) );
  FA_X1 \mult_19/S2_26_18  ( .A(\mult_19/ab[26][18] ), .B(
        \mult_19/CARRYB[25][18] ), .CI(\mult_19/SUMB[25][19] ), .CO(
        \mult_19/CARRYB[26][18] ), .S(\mult_19/SUMB[26][18] ) );
  FA_X1 \mult_19/S2_26_17  ( .A(\mult_19/ab[26][17] ), .B(
        \mult_19/CARRYB[25][17] ), .CI(\mult_19/SUMB[25][18] ), .CO(
        \mult_19/CARRYB[26][17] ), .S(\mult_19/SUMB[26][17] ) );
  FA_X1 \mult_19/S2_26_16  ( .A(\mult_19/ab[26][16] ), .B(
        \mult_19/CARRYB[25][16] ), .CI(\mult_19/SUMB[25][17] ), .CO(
        \mult_19/CARRYB[26][16] ), .S(\mult_19/SUMB[26][16] ) );
  FA_X1 \mult_19/S2_26_15  ( .A(\mult_19/ab[26][15] ), .B(
        \mult_19/CARRYB[25][15] ), .CI(\mult_19/SUMB[25][16] ), .CO(
        \mult_19/CARRYB[26][15] ), .S(\mult_19/SUMB[26][15] ) );
  FA_X1 \mult_19/S2_26_14  ( .A(\mult_19/ab[26][14] ), .B(
        \mult_19/CARRYB[25][14] ), .CI(\mult_19/SUMB[25][15] ), .CO(
        \mult_19/CARRYB[26][14] ), .S(\mult_19/SUMB[26][14] ) );
  FA_X1 \mult_19/S2_26_13  ( .A(\mult_19/ab[26][13] ), .B(
        \mult_19/CARRYB[25][13] ), .CI(\mult_19/SUMB[25][14] ), .CO(
        \mult_19/CARRYB[26][13] ), .S(\mult_19/SUMB[26][13] ) );
  FA_X1 \mult_19/S2_26_12  ( .A(\mult_19/ab[26][12] ), .B(
        \mult_19/CARRYB[25][12] ), .CI(\mult_19/SUMB[25][13] ), .CO(
        \mult_19/CARRYB[26][12] ), .S(\mult_19/SUMB[26][12] ) );
  FA_X1 \mult_19/S2_26_11  ( .A(\mult_19/ab[26][11] ), .B(
        \mult_19/CARRYB[25][11] ), .CI(\mult_19/SUMB[25][12] ), .CO(
        \mult_19/CARRYB[26][11] ), .S(\mult_19/SUMB[26][11] ) );
  FA_X1 \mult_19/S2_26_10  ( .A(\mult_19/ab[26][10] ), .B(
        \mult_19/CARRYB[25][10] ), .CI(\mult_19/SUMB[25][11] ), .CO(
        \mult_19/CARRYB[26][10] ), .S(\mult_19/SUMB[26][10] ) );
  FA_X1 \mult_19/S2_26_9  ( .A(\mult_19/ab[26][9] ), .B(
        \mult_19/CARRYB[25][9] ), .CI(\mult_19/SUMB[25][10] ), .CO(
        \mult_19/CARRYB[26][9] ), .S(\mult_19/SUMB[26][9] ) );
  FA_X1 \mult_19/S2_26_8  ( .A(\mult_19/ab[26][8] ), .B(
        \mult_19/CARRYB[25][8] ), .CI(\mult_19/SUMB[25][9] ), .CO(
        \mult_19/CARRYB[26][8] ), .S(\mult_19/SUMB[26][8] ) );
  FA_X1 \mult_19/S2_26_7  ( .A(\mult_19/ab[26][7] ), .B(
        \mult_19/CARRYB[25][7] ), .CI(\mult_19/SUMB[25][8] ), .CO(
        \mult_19/CARRYB[26][7] ), .S(\mult_19/SUMB[26][7] ) );
  FA_X1 \mult_19/S2_26_6  ( .A(\mult_19/ab[26][6] ), .B(
        \mult_19/CARRYB[25][6] ), .CI(\mult_19/SUMB[25][7] ), .CO(
        \mult_19/CARRYB[26][6] ), .S(\mult_19/SUMB[26][6] ) );
  FA_X1 \mult_19/S2_26_5  ( .A(\mult_19/ab[26][5] ), .B(
        \mult_19/CARRYB[25][5] ), .CI(\mult_19/SUMB[25][6] ), .CO(
        \mult_19/CARRYB[26][5] ), .S(\mult_19/SUMB[26][5] ) );
  FA_X1 \mult_19/S2_26_4  ( .A(\mult_19/ab[26][4] ), .B(
        \mult_19/CARRYB[25][4] ), .CI(\mult_19/SUMB[25][5] ), .CO(
        \mult_19/CARRYB[26][4] ), .S(\mult_19/SUMB[26][4] ) );
  FA_X1 \mult_19/S2_26_3  ( .A(\mult_19/ab[26][3] ), .B(
        \mult_19/CARRYB[25][3] ), .CI(\mult_19/SUMB[25][4] ), .CO(
        \mult_19/CARRYB[26][3] ), .S(\mult_19/SUMB[26][3] ) );
  FA_X1 \mult_19/S2_26_2  ( .A(\mult_19/ab[26][2] ), .B(
        \mult_19/CARRYB[25][2] ), .CI(\mult_19/SUMB[25][3] ), .CO(
        \mult_19/CARRYB[26][2] ), .S(\mult_19/SUMB[26][2] ) );
  FA_X1 \mult_19/S2_26_1  ( .A(\mult_19/ab[26][1] ), .B(
        \mult_19/CARRYB[25][1] ), .CI(\mult_19/SUMB[25][2] ), .CO(
        \mult_19/CARRYB[26][1] ), .S(\mult_19/SUMB[26][1] ) );
  FA_X1 \mult_19/S1_26_0  ( .A(\mult_19/ab[26][0] ), .B(
        \mult_19/CARRYB[25][0] ), .CI(\mult_19/SUMB[25][1] ), .CO(
        \mult_19/CARRYB[26][0] ), .S(N26) );
  FA_X1 \mult_19/S3_27_30  ( .A(\mult_19/ab[27][30] ), .B(
        \mult_19/CARRYB[26][30] ), .CI(\mult_19/ab[26][31] ), .CO(
        \mult_19/CARRYB[27][30] ), .S(\mult_19/SUMB[27][30] ) );
  FA_X1 \mult_19/S2_27_29  ( .A(\mult_19/ab[27][29] ), .B(
        \mult_19/CARRYB[26][29] ), .CI(\mult_19/SUMB[26][30] ), .CO(
        \mult_19/CARRYB[27][29] ), .S(\mult_19/SUMB[27][29] ) );
  FA_X1 \mult_19/S2_27_28  ( .A(\mult_19/ab[27][28] ), .B(
        \mult_19/CARRYB[26][28] ), .CI(\mult_19/SUMB[26][29] ), .CO(
        \mult_19/CARRYB[27][28] ), .S(\mult_19/SUMB[27][28] ) );
  FA_X1 \mult_19/S2_27_27  ( .A(\mult_19/ab[27][27] ), .B(
        \mult_19/CARRYB[26][27] ), .CI(\mult_19/SUMB[26][28] ), .CO(
        \mult_19/CARRYB[27][27] ), .S(\mult_19/SUMB[27][27] ) );
  FA_X1 \mult_19/S2_27_26  ( .A(\mult_19/ab[27][26] ), .B(
        \mult_19/CARRYB[26][26] ), .CI(\mult_19/SUMB[26][27] ), .CO(
        \mult_19/CARRYB[27][26] ), .S(\mult_19/SUMB[27][26] ) );
  FA_X1 \mult_19/S2_27_25  ( .A(\mult_19/ab[27][25] ), .B(
        \mult_19/CARRYB[26][25] ), .CI(\mult_19/SUMB[26][26] ), .CO(
        \mult_19/CARRYB[27][25] ), .S(\mult_19/SUMB[27][25] ) );
  FA_X1 \mult_19/S2_27_24  ( .A(\mult_19/ab[27][24] ), .B(
        \mult_19/CARRYB[26][24] ), .CI(\mult_19/SUMB[26][25] ), .CO(
        \mult_19/CARRYB[27][24] ), .S(\mult_19/SUMB[27][24] ) );
  FA_X1 \mult_19/S2_27_23  ( .A(\mult_19/ab[27][23] ), .B(
        \mult_19/CARRYB[26][23] ), .CI(\mult_19/SUMB[26][24] ), .CO(
        \mult_19/CARRYB[27][23] ), .S(\mult_19/SUMB[27][23] ) );
  FA_X1 \mult_19/S2_27_22  ( .A(\mult_19/ab[27][22] ), .B(
        \mult_19/CARRYB[26][22] ), .CI(\mult_19/SUMB[26][23] ), .CO(
        \mult_19/CARRYB[27][22] ), .S(\mult_19/SUMB[27][22] ) );
  FA_X1 \mult_19/S2_27_21  ( .A(\mult_19/ab[27][21] ), .B(
        \mult_19/CARRYB[26][21] ), .CI(\mult_19/SUMB[26][22] ), .CO(
        \mult_19/CARRYB[27][21] ), .S(\mult_19/SUMB[27][21] ) );
  FA_X1 \mult_19/S2_27_20  ( .A(\mult_19/ab[27][20] ), .B(
        \mult_19/CARRYB[26][20] ), .CI(\mult_19/SUMB[26][21] ), .CO(
        \mult_19/CARRYB[27][20] ), .S(\mult_19/SUMB[27][20] ) );
  FA_X1 \mult_19/S2_27_19  ( .A(\mult_19/ab[27][19] ), .B(
        \mult_19/CARRYB[26][19] ), .CI(\mult_19/SUMB[26][20] ), .CO(
        \mult_19/CARRYB[27][19] ), .S(\mult_19/SUMB[27][19] ) );
  FA_X1 \mult_19/S2_27_18  ( .A(\mult_19/ab[27][18] ), .B(
        \mult_19/CARRYB[26][18] ), .CI(\mult_19/SUMB[26][19] ), .CO(
        \mult_19/CARRYB[27][18] ), .S(\mult_19/SUMB[27][18] ) );
  FA_X1 \mult_19/S2_27_17  ( .A(\mult_19/ab[27][17] ), .B(
        \mult_19/CARRYB[26][17] ), .CI(\mult_19/SUMB[26][18] ), .CO(
        \mult_19/CARRYB[27][17] ), .S(\mult_19/SUMB[27][17] ) );
  FA_X1 \mult_19/S2_27_16  ( .A(\mult_19/ab[27][16] ), .B(
        \mult_19/CARRYB[26][16] ), .CI(\mult_19/SUMB[26][17] ), .CO(
        \mult_19/CARRYB[27][16] ), .S(\mult_19/SUMB[27][16] ) );
  FA_X1 \mult_19/S2_27_15  ( .A(\mult_19/ab[27][15] ), .B(
        \mult_19/CARRYB[26][15] ), .CI(\mult_19/SUMB[26][16] ), .CO(
        \mult_19/CARRYB[27][15] ), .S(\mult_19/SUMB[27][15] ) );
  FA_X1 \mult_19/S2_27_14  ( .A(\mult_19/ab[27][14] ), .B(
        \mult_19/CARRYB[26][14] ), .CI(\mult_19/SUMB[26][15] ), .CO(
        \mult_19/CARRYB[27][14] ), .S(\mult_19/SUMB[27][14] ) );
  FA_X1 \mult_19/S2_27_13  ( .A(\mult_19/ab[27][13] ), .B(
        \mult_19/CARRYB[26][13] ), .CI(\mult_19/SUMB[26][14] ), .CO(
        \mult_19/CARRYB[27][13] ), .S(\mult_19/SUMB[27][13] ) );
  FA_X1 \mult_19/S2_27_12  ( .A(\mult_19/ab[27][12] ), .B(
        \mult_19/CARRYB[26][12] ), .CI(\mult_19/SUMB[26][13] ), .CO(
        \mult_19/CARRYB[27][12] ), .S(\mult_19/SUMB[27][12] ) );
  FA_X1 \mult_19/S2_27_11  ( .A(\mult_19/ab[27][11] ), .B(
        \mult_19/CARRYB[26][11] ), .CI(\mult_19/SUMB[26][12] ), .CO(
        \mult_19/CARRYB[27][11] ), .S(\mult_19/SUMB[27][11] ) );
  FA_X1 \mult_19/S2_27_10  ( .A(\mult_19/ab[27][10] ), .B(
        \mult_19/CARRYB[26][10] ), .CI(\mult_19/SUMB[26][11] ), .CO(
        \mult_19/CARRYB[27][10] ), .S(\mult_19/SUMB[27][10] ) );
  FA_X1 \mult_19/S2_27_9  ( .A(\mult_19/ab[27][9] ), .B(
        \mult_19/CARRYB[26][9] ), .CI(\mult_19/SUMB[26][10] ), .CO(
        \mult_19/CARRYB[27][9] ), .S(\mult_19/SUMB[27][9] ) );
  FA_X1 \mult_19/S2_27_8  ( .A(\mult_19/ab[27][8] ), .B(
        \mult_19/CARRYB[26][8] ), .CI(\mult_19/SUMB[26][9] ), .CO(
        \mult_19/CARRYB[27][8] ), .S(\mult_19/SUMB[27][8] ) );
  FA_X1 \mult_19/S2_27_7  ( .A(\mult_19/ab[27][7] ), .B(
        \mult_19/CARRYB[26][7] ), .CI(\mult_19/SUMB[26][8] ), .CO(
        \mult_19/CARRYB[27][7] ), .S(\mult_19/SUMB[27][7] ) );
  FA_X1 \mult_19/S2_27_6  ( .A(\mult_19/ab[27][6] ), .B(
        \mult_19/CARRYB[26][6] ), .CI(\mult_19/SUMB[26][7] ), .CO(
        \mult_19/CARRYB[27][6] ), .S(\mult_19/SUMB[27][6] ) );
  FA_X1 \mult_19/S2_27_5  ( .A(\mult_19/ab[27][5] ), .B(
        \mult_19/CARRYB[26][5] ), .CI(\mult_19/SUMB[26][6] ), .CO(
        \mult_19/CARRYB[27][5] ), .S(\mult_19/SUMB[27][5] ) );
  FA_X1 \mult_19/S2_27_4  ( .A(\mult_19/ab[27][4] ), .B(
        \mult_19/CARRYB[26][4] ), .CI(\mult_19/SUMB[26][5] ), .CO(
        \mult_19/CARRYB[27][4] ), .S(\mult_19/SUMB[27][4] ) );
  FA_X1 \mult_19/S2_27_3  ( .A(\mult_19/ab[27][3] ), .B(
        \mult_19/CARRYB[26][3] ), .CI(\mult_19/SUMB[26][4] ), .CO(
        \mult_19/CARRYB[27][3] ), .S(\mult_19/SUMB[27][3] ) );
  FA_X1 \mult_19/S2_27_2  ( .A(\mult_19/ab[27][2] ), .B(
        \mult_19/CARRYB[26][2] ), .CI(\mult_19/SUMB[26][3] ), .CO(
        \mult_19/CARRYB[27][2] ), .S(\mult_19/SUMB[27][2] ) );
  FA_X1 \mult_19/S2_27_1  ( .A(\mult_19/ab[27][1] ), .B(
        \mult_19/CARRYB[26][1] ), .CI(\mult_19/SUMB[26][2] ), .CO(
        \mult_19/CARRYB[27][1] ), .S(\mult_19/SUMB[27][1] ) );
  FA_X1 \mult_19/S1_27_0  ( .A(\mult_19/ab[27][0] ), .B(
        \mult_19/CARRYB[26][0] ), .CI(\mult_19/SUMB[26][1] ), .CO(
        \mult_19/CARRYB[27][0] ), .S(N27) );
  FA_X1 \mult_19/S3_28_30  ( .A(\mult_19/ab[28][30] ), .B(
        \mult_19/CARRYB[27][30] ), .CI(\mult_19/ab[27][31] ), .CO(
        \mult_19/CARRYB[28][30] ), .S(\mult_19/SUMB[28][30] ) );
  FA_X1 \mult_19/S2_28_29  ( .A(\mult_19/ab[28][29] ), .B(
        \mult_19/CARRYB[27][29] ), .CI(\mult_19/SUMB[27][30] ), .CO(
        \mult_19/CARRYB[28][29] ), .S(\mult_19/SUMB[28][29] ) );
  FA_X1 \mult_19/S2_28_28  ( .A(\mult_19/ab[28][28] ), .B(
        \mult_19/CARRYB[27][28] ), .CI(\mult_19/SUMB[27][29] ), .CO(
        \mult_19/CARRYB[28][28] ), .S(\mult_19/SUMB[28][28] ) );
  FA_X1 \mult_19/S2_28_27  ( .A(\mult_19/ab[28][27] ), .B(
        \mult_19/CARRYB[27][27] ), .CI(\mult_19/SUMB[27][28] ), .CO(
        \mult_19/CARRYB[28][27] ), .S(\mult_19/SUMB[28][27] ) );
  FA_X1 \mult_19/S2_28_26  ( .A(\mult_19/ab[28][26] ), .B(
        \mult_19/CARRYB[27][26] ), .CI(\mult_19/SUMB[27][27] ), .CO(
        \mult_19/CARRYB[28][26] ), .S(\mult_19/SUMB[28][26] ) );
  FA_X1 \mult_19/S2_28_25  ( .A(\mult_19/ab[28][25] ), .B(
        \mult_19/CARRYB[27][25] ), .CI(\mult_19/SUMB[27][26] ), .CO(
        \mult_19/CARRYB[28][25] ), .S(\mult_19/SUMB[28][25] ) );
  FA_X1 \mult_19/S2_28_24  ( .A(\mult_19/ab[28][24] ), .B(
        \mult_19/CARRYB[27][24] ), .CI(\mult_19/SUMB[27][25] ), .CO(
        \mult_19/CARRYB[28][24] ), .S(\mult_19/SUMB[28][24] ) );
  FA_X1 \mult_19/S2_28_23  ( .A(\mult_19/ab[28][23] ), .B(
        \mult_19/CARRYB[27][23] ), .CI(\mult_19/SUMB[27][24] ), .CO(
        \mult_19/CARRYB[28][23] ), .S(\mult_19/SUMB[28][23] ) );
  FA_X1 \mult_19/S2_28_22  ( .A(\mult_19/ab[28][22] ), .B(
        \mult_19/CARRYB[27][22] ), .CI(\mult_19/SUMB[27][23] ), .CO(
        \mult_19/CARRYB[28][22] ), .S(\mult_19/SUMB[28][22] ) );
  FA_X1 \mult_19/S2_28_21  ( .A(\mult_19/ab[28][21] ), .B(
        \mult_19/CARRYB[27][21] ), .CI(\mult_19/SUMB[27][22] ), .CO(
        \mult_19/CARRYB[28][21] ), .S(\mult_19/SUMB[28][21] ) );
  FA_X1 \mult_19/S2_28_20  ( .A(\mult_19/ab[28][20] ), .B(
        \mult_19/CARRYB[27][20] ), .CI(\mult_19/SUMB[27][21] ), .CO(
        \mult_19/CARRYB[28][20] ), .S(\mult_19/SUMB[28][20] ) );
  FA_X1 \mult_19/S2_28_19  ( .A(\mult_19/ab[28][19] ), .B(
        \mult_19/CARRYB[27][19] ), .CI(\mult_19/SUMB[27][20] ), .CO(
        \mult_19/CARRYB[28][19] ), .S(\mult_19/SUMB[28][19] ) );
  FA_X1 \mult_19/S2_28_18  ( .A(\mult_19/ab[28][18] ), .B(
        \mult_19/CARRYB[27][18] ), .CI(\mult_19/SUMB[27][19] ), .CO(
        \mult_19/CARRYB[28][18] ), .S(\mult_19/SUMB[28][18] ) );
  FA_X1 \mult_19/S2_28_17  ( .A(\mult_19/ab[28][17] ), .B(
        \mult_19/CARRYB[27][17] ), .CI(\mult_19/SUMB[27][18] ), .CO(
        \mult_19/CARRYB[28][17] ), .S(\mult_19/SUMB[28][17] ) );
  FA_X1 \mult_19/S2_28_16  ( .A(\mult_19/ab[28][16] ), .B(
        \mult_19/CARRYB[27][16] ), .CI(\mult_19/SUMB[27][17] ), .CO(
        \mult_19/CARRYB[28][16] ), .S(\mult_19/SUMB[28][16] ) );
  FA_X1 \mult_19/S2_28_15  ( .A(\mult_19/ab[28][15] ), .B(
        \mult_19/CARRYB[27][15] ), .CI(\mult_19/SUMB[27][16] ), .CO(
        \mult_19/CARRYB[28][15] ), .S(\mult_19/SUMB[28][15] ) );
  FA_X1 \mult_19/S2_28_14  ( .A(\mult_19/ab[28][14] ), .B(
        \mult_19/CARRYB[27][14] ), .CI(\mult_19/SUMB[27][15] ), .CO(
        \mult_19/CARRYB[28][14] ), .S(\mult_19/SUMB[28][14] ) );
  FA_X1 \mult_19/S2_28_13  ( .A(\mult_19/ab[28][13] ), .B(
        \mult_19/CARRYB[27][13] ), .CI(\mult_19/SUMB[27][14] ), .CO(
        \mult_19/CARRYB[28][13] ), .S(\mult_19/SUMB[28][13] ) );
  FA_X1 \mult_19/S2_28_12  ( .A(\mult_19/ab[28][12] ), .B(
        \mult_19/CARRYB[27][12] ), .CI(\mult_19/SUMB[27][13] ), .CO(
        \mult_19/CARRYB[28][12] ), .S(\mult_19/SUMB[28][12] ) );
  FA_X1 \mult_19/S2_28_11  ( .A(\mult_19/ab[28][11] ), .B(
        \mult_19/CARRYB[27][11] ), .CI(\mult_19/SUMB[27][12] ), .CO(
        \mult_19/CARRYB[28][11] ), .S(\mult_19/SUMB[28][11] ) );
  FA_X1 \mult_19/S2_28_10  ( .A(\mult_19/ab[28][10] ), .B(
        \mult_19/CARRYB[27][10] ), .CI(\mult_19/SUMB[27][11] ), .CO(
        \mult_19/CARRYB[28][10] ), .S(\mult_19/SUMB[28][10] ) );
  FA_X1 \mult_19/S2_28_9  ( .A(\mult_19/ab[28][9] ), .B(
        \mult_19/CARRYB[27][9] ), .CI(\mult_19/SUMB[27][10] ), .CO(
        \mult_19/CARRYB[28][9] ), .S(\mult_19/SUMB[28][9] ) );
  FA_X1 \mult_19/S2_28_8  ( .A(\mult_19/ab[28][8] ), .B(
        \mult_19/CARRYB[27][8] ), .CI(\mult_19/SUMB[27][9] ), .CO(
        \mult_19/CARRYB[28][8] ), .S(\mult_19/SUMB[28][8] ) );
  FA_X1 \mult_19/S2_28_7  ( .A(\mult_19/ab[28][7] ), .B(
        \mult_19/CARRYB[27][7] ), .CI(\mult_19/SUMB[27][8] ), .CO(
        \mult_19/CARRYB[28][7] ), .S(\mult_19/SUMB[28][7] ) );
  FA_X1 \mult_19/S2_28_6  ( .A(\mult_19/ab[28][6] ), .B(
        \mult_19/CARRYB[27][6] ), .CI(\mult_19/SUMB[27][7] ), .CO(
        \mult_19/CARRYB[28][6] ), .S(\mult_19/SUMB[28][6] ) );
  FA_X1 \mult_19/S2_28_5  ( .A(\mult_19/ab[28][5] ), .B(
        \mult_19/CARRYB[27][5] ), .CI(\mult_19/SUMB[27][6] ), .CO(
        \mult_19/CARRYB[28][5] ), .S(\mult_19/SUMB[28][5] ) );
  FA_X1 \mult_19/S2_28_4  ( .A(\mult_19/ab[28][4] ), .B(
        \mult_19/CARRYB[27][4] ), .CI(\mult_19/SUMB[27][5] ), .CO(
        \mult_19/CARRYB[28][4] ), .S(\mult_19/SUMB[28][4] ) );
  FA_X1 \mult_19/S2_28_3  ( .A(\mult_19/ab[28][3] ), .B(
        \mult_19/CARRYB[27][3] ), .CI(\mult_19/SUMB[27][4] ), .CO(
        \mult_19/CARRYB[28][3] ), .S(\mult_19/SUMB[28][3] ) );
  FA_X1 \mult_19/S2_28_2  ( .A(\mult_19/ab[28][2] ), .B(
        \mult_19/CARRYB[27][2] ), .CI(\mult_19/SUMB[27][3] ), .CO(
        \mult_19/CARRYB[28][2] ), .S(\mult_19/SUMB[28][2] ) );
  FA_X1 \mult_19/S2_28_1  ( .A(\mult_19/ab[28][1] ), .B(
        \mult_19/CARRYB[27][1] ), .CI(\mult_19/SUMB[27][2] ), .CO(
        \mult_19/CARRYB[28][1] ), .S(\mult_19/SUMB[28][1] ) );
  FA_X1 \mult_19/S1_28_0  ( .A(\mult_19/ab[28][0] ), .B(
        \mult_19/CARRYB[27][0] ), .CI(\mult_19/SUMB[27][1] ), .CO(
        \mult_19/CARRYB[28][0] ), .S(N28) );
  FA_X1 \mult_19/S3_29_30  ( .A(\mult_19/ab[29][30] ), .B(
        \mult_19/CARRYB[28][30] ), .CI(\mult_19/ab[28][31] ), .CO(
        \mult_19/CARRYB[29][30] ), .S(\mult_19/SUMB[29][30] ) );
  FA_X1 \mult_19/S2_29_29  ( .A(\mult_19/ab[29][29] ), .B(
        \mult_19/CARRYB[28][29] ), .CI(\mult_19/SUMB[28][30] ), .CO(
        \mult_19/CARRYB[29][29] ), .S(\mult_19/SUMB[29][29] ) );
  FA_X1 \mult_19/S2_29_28  ( .A(\mult_19/ab[29][28] ), .B(
        \mult_19/CARRYB[28][28] ), .CI(\mult_19/SUMB[28][29] ), .CO(
        \mult_19/CARRYB[29][28] ), .S(\mult_19/SUMB[29][28] ) );
  FA_X1 \mult_19/S2_29_27  ( .A(\mult_19/ab[29][27] ), .B(
        \mult_19/CARRYB[28][27] ), .CI(\mult_19/SUMB[28][28] ), .CO(
        \mult_19/CARRYB[29][27] ), .S(\mult_19/SUMB[29][27] ) );
  FA_X1 \mult_19/S2_29_26  ( .A(\mult_19/ab[29][26] ), .B(
        \mult_19/CARRYB[28][26] ), .CI(\mult_19/SUMB[28][27] ), .CO(
        \mult_19/CARRYB[29][26] ), .S(\mult_19/SUMB[29][26] ) );
  FA_X1 \mult_19/S2_29_25  ( .A(\mult_19/ab[29][25] ), .B(
        \mult_19/CARRYB[28][25] ), .CI(\mult_19/SUMB[28][26] ), .CO(
        \mult_19/CARRYB[29][25] ), .S(\mult_19/SUMB[29][25] ) );
  FA_X1 \mult_19/S2_29_24  ( .A(\mult_19/ab[29][24] ), .B(
        \mult_19/CARRYB[28][24] ), .CI(\mult_19/SUMB[28][25] ), .CO(
        \mult_19/CARRYB[29][24] ), .S(\mult_19/SUMB[29][24] ) );
  FA_X1 \mult_19/S2_29_23  ( .A(\mult_19/ab[29][23] ), .B(
        \mult_19/CARRYB[28][23] ), .CI(\mult_19/SUMB[28][24] ), .CO(
        \mult_19/CARRYB[29][23] ), .S(\mult_19/SUMB[29][23] ) );
  FA_X1 \mult_19/S2_29_22  ( .A(\mult_19/ab[29][22] ), .B(
        \mult_19/CARRYB[28][22] ), .CI(\mult_19/SUMB[28][23] ), .CO(
        \mult_19/CARRYB[29][22] ), .S(\mult_19/SUMB[29][22] ) );
  FA_X1 \mult_19/S2_29_21  ( .A(\mult_19/ab[29][21] ), .B(
        \mult_19/CARRYB[28][21] ), .CI(\mult_19/SUMB[28][22] ), .CO(
        \mult_19/CARRYB[29][21] ), .S(\mult_19/SUMB[29][21] ) );
  FA_X1 \mult_19/S2_29_20  ( .A(\mult_19/ab[29][20] ), .B(
        \mult_19/CARRYB[28][20] ), .CI(\mult_19/SUMB[28][21] ), .CO(
        \mult_19/CARRYB[29][20] ), .S(\mult_19/SUMB[29][20] ) );
  FA_X1 \mult_19/S2_29_19  ( .A(\mult_19/ab[29][19] ), .B(
        \mult_19/CARRYB[28][19] ), .CI(\mult_19/SUMB[28][20] ), .CO(
        \mult_19/CARRYB[29][19] ), .S(\mult_19/SUMB[29][19] ) );
  FA_X1 \mult_19/S2_29_18  ( .A(\mult_19/ab[29][18] ), .B(
        \mult_19/CARRYB[28][18] ), .CI(\mult_19/SUMB[28][19] ), .CO(
        \mult_19/CARRYB[29][18] ), .S(\mult_19/SUMB[29][18] ) );
  FA_X1 \mult_19/S2_29_17  ( .A(\mult_19/ab[29][17] ), .B(
        \mult_19/CARRYB[28][17] ), .CI(\mult_19/SUMB[28][18] ), .CO(
        \mult_19/CARRYB[29][17] ), .S(\mult_19/SUMB[29][17] ) );
  FA_X1 \mult_19/S2_29_16  ( .A(\mult_19/ab[29][16] ), .B(
        \mult_19/CARRYB[28][16] ), .CI(\mult_19/SUMB[28][17] ), .CO(
        \mult_19/CARRYB[29][16] ), .S(\mult_19/SUMB[29][16] ) );
  FA_X1 \mult_19/S2_29_15  ( .A(\mult_19/ab[29][15] ), .B(
        \mult_19/CARRYB[28][15] ), .CI(\mult_19/SUMB[28][16] ), .CO(
        \mult_19/CARRYB[29][15] ), .S(\mult_19/SUMB[29][15] ) );
  FA_X1 \mult_19/S2_29_14  ( .A(\mult_19/ab[29][14] ), .B(
        \mult_19/CARRYB[28][14] ), .CI(\mult_19/SUMB[28][15] ), .CO(
        \mult_19/CARRYB[29][14] ), .S(\mult_19/SUMB[29][14] ) );
  FA_X1 \mult_19/S2_29_13  ( .A(\mult_19/ab[29][13] ), .B(
        \mult_19/CARRYB[28][13] ), .CI(\mult_19/SUMB[28][14] ), .CO(
        \mult_19/CARRYB[29][13] ), .S(\mult_19/SUMB[29][13] ) );
  FA_X1 \mult_19/S2_29_12  ( .A(\mult_19/ab[29][12] ), .B(
        \mult_19/CARRYB[28][12] ), .CI(\mult_19/SUMB[28][13] ), .CO(
        \mult_19/CARRYB[29][12] ), .S(\mult_19/SUMB[29][12] ) );
  FA_X1 \mult_19/S2_29_11  ( .A(\mult_19/ab[29][11] ), .B(
        \mult_19/CARRYB[28][11] ), .CI(\mult_19/SUMB[28][12] ), .CO(
        \mult_19/CARRYB[29][11] ), .S(\mult_19/SUMB[29][11] ) );
  FA_X1 \mult_19/S2_29_10  ( .A(\mult_19/ab[29][10] ), .B(
        \mult_19/CARRYB[28][10] ), .CI(\mult_19/SUMB[28][11] ), .CO(
        \mult_19/CARRYB[29][10] ), .S(\mult_19/SUMB[29][10] ) );
  FA_X1 \mult_19/S2_29_9  ( .A(\mult_19/ab[29][9] ), .B(
        \mult_19/CARRYB[28][9] ), .CI(\mult_19/SUMB[28][10] ), .CO(
        \mult_19/CARRYB[29][9] ), .S(\mult_19/SUMB[29][9] ) );
  FA_X1 \mult_19/S2_29_8  ( .A(\mult_19/ab[29][8] ), .B(
        \mult_19/CARRYB[28][8] ), .CI(\mult_19/SUMB[28][9] ), .CO(
        \mult_19/CARRYB[29][8] ), .S(\mult_19/SUMB[29][8] ) );
  FA_X1 \mult_19/S2_29_7  ( .A(\mult_19/ab[29][7] ), .B(
        \mult_19/CARRYB[28][7] ), .CI(\mult_19/SUMB[28][8] ), .CO(
        \mult_19/CARRYB[29][7] ), .S(\mult_19/SUMB[29][7] ) );
  FA_X1 \mult_19/S2_29_6  ( .A(\mult_19/ab[29][6] ), .B(
        \mult_19/CARRYB[28][6] ), .CI(\mult_19/SUMB[28][7] ), .CO(
        \mult_19/CARRYB[29][6] ), .S(\mult_19/SUMB[29][6] ) );
  FA_X1 \mult_19/S2_29_5  ( .A(\mult_19/ab[29][5] ), .B(
        \mult_19/CARRYB[28][5] ), .CI(\mult_19/SUMB[28][6] ), .CO(
        \mult_19/CARRYB[29][5] ), .S(\mult_19/SUMB[29][5] ) );
  FA_X1 \mult_19/S2_29_4  ( .A(\mult_19/ab[29][4] ), .B(
        \mult_19/CARRYB[28][4] ), .CI(\mult_19/SUMB[28][5] ), .CO(
        \mult_19/CARRYB[29][4] ), .S(\mult_19/SUMB[29][4] ) );
  FA_X1 \mult_19/S2_29_3  ( .A(\mult_19/ab[29][3] ), .B(
        \mult_19/CARRYB[28][3] ), .CI(\mult_19/SUMB[28][4] ), .CO(
        \mult_19/CARRYB[29][3] ), .S(\mult_19/SUMB[29][3] ) );
  FA_X1 \mult_19/S2_29_2  ( .A(\mult_19/ab[29][2] ), .B(
        \mult_19/CARRYB[28][2] ), .CI(\mult_19/SUMB[28][3] ), .CO(
        \mult_19/CARRYB[29][2] ), .S(\mult_19/SUMB[29][2] ) );
  FA_X1 \mult_19/S2_29_1  ( .A(\mult_19/ab[29][1] ), .B(
        \mult_19/CARRYB[28][1] ), .CI(\mult_19/SUMB[28][2] ), .CO(
        \mult_19/CARRYB[29][1] ), .S(\mult_19/SUMB[29][1] ) );
  FA_X1 \mult_19/S1_29_0  ( .A(\mult_19/ab[29][0] ), .B(
        \mult_19/CARRYB[28][0] ), .CI(\mult_19/SUMB[28][1] ), .CO(
        \mult_19/CARRYB[29][0] ), .S(N29) );
  FA_X1 \mult_19/S3_30_30  ( .A(\mult_19/ab[30][30] ), .B(
        \mult_19/CARRYB[29][30] ), .CI(\mult_19/ab[29][31] ), .CO(
        \mult_19/CARRYB[30][30] ), .S(\mult_19/SUMB[30][30] ) );
  FA_X1 \mult_19/S2_30_29  ( .A(\mult_19/ab[30][29] ), .B(
        \mult_19/CARRYB[29][29] ), .CI(\mult_19/SUMB[29][30] ), .CO(
        \mult_19/CARRYB[30][29] ), .S(\mult_19/SUMB[30][29] ) );
  FA_X1 \mult_19/S2_30_28  ( .A(\mult_19/ab[30][28] ), .B(
        \mult_19/CARRYB[29][28] ), .CI(\mult_19/SUMB[29][29] ), .CO(
        \mult_19/CARRYB[30][28] ), .S(\mult_19/SUMB[30][28] ) );
  FA_X1 \mult_19/S2_30_27  ( .A(\mult_19/ab[30][27] ), .B(
        \mult_19/CARRYB[29][27] ), .CI(\mult_19/SUMB[29][28] ), .CO(
        \mult_19/CARRYB[30][27] ), .S(\mult_19/SUMB[30][27] ) );
  FA_X1 \mult_19/S2_30_26  ( .A(\mult_19/ab[30][26] ), .B(
        \mult_19/CARRYB[29][26] ), .CI(\mult_19/SUMB[29][27] ), .CO(
        \mult_19/CARRYB[30][26] ), .S(\mult_19/SUMB[30][26] ) );
  FA_X1 \mult_19/S2_30_25  ( .A(\mult_19/ab[30][25] ), .B(
        \mult_19/CARRYB[29][25] ), .CI(\mult_19/SUMB[29][26] ), .CO(
        \mult_19/CARRYB[30][25] ), .S(\mult_19/SUMB[30][25] ) );
  FA_X1 \mult_19/S2_30_24  ( .A(\mult_19/ab[30][24] ), .B(
        \mult_19/CARRYB[29][24] ), .CI(\mult_19/SUMB[29][25] ), .CO(
        \mult_19/CARRYB[30][24] ), .S(\mult_19/SUMB[30][24] ) );
  FA_X1 \mult_19/S2_30_23  ( .A(\mult_19/ab[30][23] ), .B(
        \mult_19/CARRYB[29][23] ), .CI(\mult_19/SUMB[29][24] ), .CO(
        \mult_19/CARRYB[30][23] ), .S(\mult_19/SUMB[30][23] ) );
  FA_X1 \mult_19/S2_30_22  ( .A(\mult_19/ab[30][22] ), .B(
        \mult_19/CARRYB[29][22] ), .CI(\mult_19/SUMB[29][23] ), .CO(
        \mult_19/CARRYB[30][22] ), .S(\mult_19/SUMB[30][22] ) );
  FA_X1 \mult_19/S2_30_21  ( .A(\mult_19/ab[30][21] ), .B(
        \mult_19/CARRYB[29][21] ), .CI(\mult_19/SUMB[29][22] ), .CO(
        \mult_19/CARRYB[30][21] ), .S(\mult_19/SUMB[30][21] ) );
  FA_X1 \mult_19/S2_30_20  ( .A(\mult_19/ab[30][20] ), .B(
        \mult_19/CARRYB[29][20] ), .CI(\mult_19/SUMB[29][21] ), .CO(
        \mult_19/CARRYB[30][20] ), .S(\mult_19/SUMB[30][20] ) );
  FA_X1 \mult_19/S2_30_19  ( .A(\mult_19/ab[30][19] ), .B(
        \mult_19/CARRYB[29][19] ), .CI(\mult_19/SUMB[29][20] ), .CO(
        \mult_19/CARRYB[30][19] ), .S(\mult_19/SUMB[30][19] ) );
  FA_X1 \mult_19/S2_30_18  ( .A(\mult_19/ab[30][18] ), .B(
        \mult_19/CARRYB[29][18] ), .CI(\mult_19/SUMB[29][19] ), .CO(
        \mult_19/CARRYB[30][18] ), .S(\mult_19/SUMB[30][18] ) );
  FA_X1 \mult_19/S2_30_17  ( .A(\mult_19/ab[30][17] ), .B(
        \mult_19/CARRYB[29][17] ), .CI(\mult_19/SUMB[29][18] ), .CO(
        \mult_19/CARRYB[30][17] ), .S(\mult_19/SUMB[30][17] ) );
  FA_X1 \mult_19/S2_30_16  ( .A(\mult_19/ab[30][16] ), .B(
        \mult_19/CARRYB[29][16] ), .CI(\mult_19/SUMB[29][17] ), .CO(
        \mult_19/CARRYB[30][16] ), .S(\mult_19/SUMB[30][16] ) );
  FA_X1 \mult_19/S2_30_15  ( .A(\mult_19/ab[30][15] ), .B(
        \mult_19/CARRYB[29][15] ), .CI(\mult_19/SUMB[29][16] ), .CO(
        \mult_19/CARRYB[30][15] ), .S(\mult_19/SUMB[30][15] ) );
  FA_X1 \mult_19/S2_30_14  ( .A(\mult_19/ab[30][14] ), .B(
        \mult_19/CARRYB[29][14] ), .CI(\mult_19/SUMB[29][15] ), .CO(
        \mult_19/CARRYB[30][14] ), .S(\mult_19/SUMB[30][14] ) );
  FA_X1 \mult_19/S2_30_13  ( .A(\mult_19/ab[30][13] ), .B(
        \mult_19/CARRYB[29][13] ), .CI(\mult_19/SUMB[29][14] ), .CO(
        \mult_19/CARRYB[30][13] ), .S(\mult_19/SUMB[30][13] ) );
  FA_X1 \mult_19/S2_30_12  ( .A(\mult_19/ab[30][12] ), .B(
        \mult_19/CARRYB[29][12] ), .CI(\mult_19/SUMB[29][13] ), .CO(
        \mult_19/CARRYB[30][12] ), .S(\mult_19/SUMB[30][12] ) );
  FA_X1 \mult_19/S2_30_11  ( .A(\mult_19/ab[30][11] ), .B(
        \mult_19/CARRYB[29][11] ), .CI(\mult_19/SUMB[29][12] ), .CO(
        \mult_19/CARRYB[30][11] ), .S(\mult_19/SUMB[30][11] ) );
  FA_X1 \mult_19/S2_30_10  ( .A(\mult_19/ab[30][10] ), .B(
        \mult_19/CARRYB[29][10] ), .CI(\mult_19/SUMB[29][11] ), .CO(
        \mult_19/CARRYB[30][10] ), .S(\mult_19/SUMB[30][10] ) );
  FA_X1 \mult_19/S2_30_9  ( .A(\mult_19/ab[30][9] ), .B(
        \mult_19/CARRYB[29][9] ), .CI(\mult_19/SUMB[29][10] ), .CO(
        \mult_19/CARRYB[30][9] ), .S(\mult_19/SUMB[30][9] ) );
  FA_X1 \mult_19/S2_30_8  ( .A(\mult_19/ab[30][8] ), .B(
        \mult_19/CARRYB[29][8] ), .CI(\mult_19/SUMB[29][9] ), .CO(
        \mult_19/CARRYB[30][8] ), .S(\mult_19/SUMB[30][8] ) );
  FA_X1 \mult_19/S2_30_7  ( .A(\mult_19/ab[30][7] ), .B(
        \mult_19/CARRYB[29][7] ), .CI(\mult_19/SUMB[29][8] ), .CO(
        \mult_19/CARRYB[30][7] ), .S(\mult_19/SUMB[30][7] ) );
  FA_X1 \mult_19/S2_30_6  ( .A(\mult_19/ab[30][6] ), .B(
        \mult_19/CARRYB[29][6] ), .CI(\mult_19/SUMB[29][7] ), .CO(
        \mult_19/CARRYB[30][6] ), .S(\mult_19/SUMB[30][6] ) );
  FA_X1 \mult_19/S2_30_5  ( .A(\mult_19/ab[30][5] ), .B(
        \mult_19/CARRYB[29][5] ), .CI(\mult_19/SUMB[29][6] ), .CO(
        \mult_19/CARRYB[30][5] ), .S(\mult_19/SUMB[30][5] ) );
  FA_X1 \mult_19/S2_30_4  ( .A(\mult_19/ab[30][4] ), .B(
        \mult_19/CARRYB[29][4] ), .CI(\mult_19/SUMB[29][5] ), .CO(
        \mult_19/CARRYB[30][4] ), .S(\mult_19/SUMB[30][4] ) );
  FA_X1 \mult_19/S2_30_3  ( .A(\mult_19/ab[30][3] ), .B(
        \mult_19/CARRYB[29][3] ), .CI(\mult_19/SUMB[29][4] ), .CO(
        \mult_19/CARRYB[30][3] ), .S(\mult_19/SUMB[30][3] ) );
  FA_X1 \mult_19/S2_30_2  ( .A(\mult_19/ab[30][2] ), .B(
        \mult_19/CARRYB[29][2] ), .CI(\mult_19/SUMB[29][3] ), .CO(
        \mult_19/CARRYB[30][2] ), .S(\mult_19/SUMB[30][2] ) );
  FA_X1 \mult_19/S2_30_1  ( .A(\mult_19/ab[30][1] ), .B(
        \mult_19/CARRYB[29][1] ), .CI(\mult_19/SUMB[29][2] ), .CO(
        \mult_19/CARRYB[30][1] ), .S(\mult_19/SUMB[30][1] ) );
  FA_X1 \mult_19/S1_30_0  ( .A(\mult_19/ab[30][0] ), .B(
        \mult_19/CARRYB[29][0] ), .CI(\mult_19/SUMB[29][1] ), .CO(
        \mult_19/CARRYB[30][0] ), .S(N30) );
  FA_X1 \mult_19/S5_30  ( .A(\mult_19/ab[31][30] ), .B(
        \mult_19/CARRYB[30][30] ), .CI(\mult_19/ab[30][31] ), .CO(
        \mult_19/CARRYB[31][30] ), .S(\mult_19/SUMB[31][30] ) );
  FA_X1 \mult_19/S4_29  ( .A(\mult_19/ab[31][29] ), .B(
        \mult_19/CARRYB[30][29] ), .CI(\mult_19/SUMB[30][30] ), .CO(
        \mult_19/CARRYB[31][29] ), .S(\mult_19/SUMB[31][29] ) );
  FA_X1 \mult_19/S4_28  ( .A(\mult_19/ab[31][28] ), .B(
        \mult_19/CARRYB[30][28] ), .CI(\mult_19/SUMB[30][29] ), .CO(
        \mult_19/CARRYB[31][28] ), .S(\mult_19/SUMB[31][28] ) );
  FA_X1 \mult_19/S4_27  ( .A(\mult_19/ab[31][27] ), .B(
        \mult_19/CARRYB[30][27] ), .CI(\mult_19/SUMB[30][28] ), .CO(
        \mult_19/CARRYB[31][27] ), .S(\mult_19/SUMB[31][27] ) );
  FA_X1 \mult_19/S4_26  ( .A(\mult_19/ab[31][26] ), .B(
        \mult_19/CARRYB[30][26] ), .CI(\mult_19/SUMB[30][27] ), .CO(
        \mult_19/CARRYB[31][26] ), .S(\mult_19/SUMB[31][26] ) );
  FA_X1 \mult_19/S4_25  ( .A(\mult_19/ab[31][25] ), .B(
        \mult_19/CARRYB[30][25] ), .CI(\mult_19/SUMB[30][26] ), .CO(
        \mult_19/CARRYB[31][25] ), .S(\mult_19/SUMB[31][25] ) );
  FA_X1 \mult_19/S4_24  ( .A(\mult_19/ab[31][24] ), .B(
        \mult_19/CARRYB[30][24] ), .CI(\mult_19/SUMB[30][25] ), .CO(
        \mult_19/CARRYB[31][24] ), .S(\mult_19/SUMB[31][24] ) );
  FA_X1 \mult_19/S4_23  ( .A(\mult_19/ab[31][23] ), .B(
        \mult_19/CARRYB[30][23] ), .CI(\mult_19/SUMB[30][24] ), .CO(
        \mult_19/CARRYB[31][23] ), .S(\mult_19/SUMB[31][23] ) );
  FA_X1 \mult_19/S4_22  ( .A(\mult_19/ab[31][22] ), .B(
        \mult_19/CARRYB[30][22] ), .CI(\mult_19/SUMB[30][23] ), .CO(
        \mult_19/CARRYB[31][22] ), .S(\mult_19/SUMB[31][22] ) );
  FA_X1 \mult_19/S4_21  ( .A(\mult_19/ab[31][21] ), .B(
        \mult_19/CARRYB[30][21] ), .CI(\mult_19/SUMB[30][22] ), .CO(
        \mult_19/CARRYB[31][21] ), .S(\mult_19/SUMB[31][21] ) );
  FA_X1 \mult_19/S4_20  ( .A(\mult_19/ab[31][20] ), .B(
        \mult_19/CARRYB[30][20] ), .CI(\mult_19/SUMB[30][21] ), .CO(
        \mult_19/CARRYB[31][20] ), .S(\mult_19/SUMB[31][20] ) );
  FA_X1 \mult_19/S4_19  ( .A(\mult_19/ab[31][19] ), .B(
        \mult_19/CARRYB[30][19] ), .CI(\mult_19/SUMB[30][20] ), .CO(
        \mult_19/CARRYB[31][19] ), .S(\mult_19/SUMB[31][19] ) );
  FA_X1 \mult_19/S4_18  ( .A(\mult_19/ab[31][18] ), .B(
        \mult_19/CARRYB[30][18] ), .CI(\mult_19/SUMB[30][19] ), .CO(
        \mult_19/CARRYB[31][18] ), .S(\mult_19/SUMB[31][18] ) );
  FA_X1 \mult_19/S4_17  ( .A(\mult_19/ab[31][17] ), .B(
        \mult_19/CARRYB[30][17] ), .CI(\mult_19/SUMB[30][18] ), .CO(
        \mult_19/CARRYB[31][17] ), .S(\mult_19/SUMB[31][17] ) );
  FA_X1 \mult_19/S4_16  ( .A(\mult_19/ab[31][16] ), .B(
        \mult_19/CARRYB[30][16] ), .CI(\mult_19/SUMB[30][17] ), .CO(
        \mult_19/CARRYB[31][16] ), .S(\mult_19/SUMB[31][16] ) );
  FA_X1 \mult_19/S4_15  ( .A(\mult_19/ab[31][15] ), .B(
        \mult_19/CARRYB[30][15] ), .CI(\mult_19/SUMB[30][16] ), .CO(
        \mult_19/CARRYB[31][15] ), .S(\mult_19/SUMB[31][15] ) );
  FA_X1 \mult_19/S4_14  ( .A(\mult_19/ab[31][14] ), .B(
        \mult_19/CARRYB[30][14] ), .CI(\mult_19/SUMB[30][15] ), .CO(
        \mult_19/CARRYB[31][14] ), .S(\mult_19/SUMB[31][14] ) );
  FA_X1 \mult_19/S4_13  ( .A(\mult_19/ab[31][13] ), .B(
        \mult_19/CARRYB[30][13] ), .CI(\mult_19/SUMB[30][14] ), .CO(
        \mult_19/CARRYB[31][13] ), .S(\mult_19/SUMB[31][13] ) );
  FA_X1 \mult_19/S4_12  ( .A(\mult_19/ab[31][12] ), .B(
        \mult_19/CARRYB[30][12] ), .CI(\mult_19/SUMB[30][13] ), .CO(
        \mult_19/CARRYB[31][12] ), .S(\mult_19/SUMB[31][12] ) );
  FA_X1 \mult_19/S4_11  ( .A(\mult_19/ab[31][11] ), .B(
        \mult_19/CARRYB[30][11] ), .CI(\mult_19/SUMB[30][12] ), .CO(
        \mult_19/CARRYB[31][11] ), .S(\mult_19/SUMB[31][11] ) );
  FA_X1 \mult_19/S4_10  ( .A(\mult_19/ab[31][10] ), .B(
        \mult_19/CARRYB[30][10] ), .CI(\mult_19/SUMB[30][11] ), .CO(
        \mult_19/CARRYB[31][10] ), .S(\mult_19/SUMB[31][10] ) );
  FA_X1 \mult_19/S4_9  ( .A(\mult_19/ab[31][9] ), .B(\mult_19/CARRYB[30][9] ), 
        .CI(\mult_19/SUMB[30][10] ), .CO(\mult_19/CARRYB[31][9] ), .S(
        \mult_19/SUMB[31][9] ) );
  FA_X1 \mult_19/S4_8  ( .A(\mult_19/ab[31][8] ), .B(\mult_19/CARRYB[30][8] ), 
        .CI(\mult_19/SUMB[30][9] ), .CO(\mult_19/CARRYB[31][8] ), .S(
        \mult_19/SUMB[31][8] ) );
  FA_X1 \mult_19/S4_7  ( .A(\mult_19/ab[31][7] ), .B(\mult_19/CARRYB[30][7] ), 
        .CI(\mult_19/SUMB[30][8] ), .CO(\mult_19/CARRYB[31][7] ), .S(
        \mult_19/SUMB[31][7] ) );
  FA_X1 \mult_19/S4_6  ( .A(\mult_19/ab[31][6] ), .B(\mult_19/CARRYB[30][6] ), 
        .CI(\mult_19/SUMB[30][7] ), .CO(\mult_19/CARRYB[31][6] ), .S(
        \mult_19/SUMB[31][6] ) );
  FA_X1 \mult_19/S4_5  ( .A(\mult_19/ab[31][5] ), .B(\mult_19/CARRYB[30][5] ), 
        .CI(\mult_19/SUMB[30][6] ), .CO(\mult_19/CARRYB[31][5] ), .S(
        \mult_19/SUMB[31][5] ) );
  FA_X1 \mult_19/S4_4  ( .A(\mult_19/ab[31][4] ), .B(\mult_19/CARRYB[30][4] ), 
        .CI(\mult_19/SUMB[30][5] ), .CO(\mult_19/CARRYB[31][4] ), .S(
        \mult_19/SUMB[31][4] ) );
  FA_X1 \mult_19/S4_3  ( .A(\mult_19/ab[31][3] ), .B(\mult_19/CARRYB[30][3] ), 
        .CI(\mult_19/SUMB[30][4] ), .CO(\mult_19/CARRYB[31][3] ), .S(
        \mult_19/SUMB[31][3] ) );
  FA_X1 \mult_19/S4_2  ( .A(\mult_19/ab[31][2] ), .B(\mult_19/CARRYB[30][2] ), 
        .CI(\mult_19/SUMB[30][3] ), .CO(\mult_19/CARRYB[31][2] ), .S(
        \mult_19/SUMB[31][2] ) );
  FA_X1 \mult_19/S4_1  ( .A(\mult_19/ab[31][1] ), .B(\mult_19/CARRYB[30][1] ), 
        .CI(\mult_19/SUMB[30][2] ), .CO(\mult_19/CARRYB[31][1] ), .S(
        \mult_19/SUMB[31][1] ) );
  FA_X1 \mult_19/S4_0  ( .A(\mult_19/ab[31][0] ), .B(\mult_19/CARRYB[30][0] ), 
        .CI(\mult_19/SUMB[30][1] ), .CO(\mult_19/CARRYB[31][0] ), .S(N31) );
  FA_X1 \mult_22/S3_2_62  ( .A(\mult_22/ab[2][62] ), .B(\mult_22/n181 ), .CI(
        \mult_22/ab[1][63] ), .CO(\mult_22/CARRYB[2][62] ), .S(
        \mult_22/SUMB[2][62] ) );
  FA_X1 \mult_22/S2_2_61  ( .A(n1800), .B(\mult_22/ab[2][61] ), .CI(
        \mult_22/n325 ), .CO(\mult_22/CARRYB[2][61] ), .S(
        \mult_22/SUMB[2][61] ) );
  FA_X1 \mult_22/S2_2_60  ( .A(\mult_22/n323 ), .B(\mult_22/ab[2][60] ), .CI(
        \mult_22/SUMB[1][61] ), .CO(\mult_22/CARRYB[2][60] ), .S(
        \mult_22/SUMB[2][60] ) );
  FA_X1 \mult_22/S2_2_59  ( .A(\mult_22/ab[2][59] ), .B(\mult_22/n163 ), .CI(
        \mult_22/n196 ), .CO(\mult_22/CARRYB[2][59] ), .S(
        \mult_22/SUMB[2][59] ) );
  FA_X1 \mult_22/S2_2_58  ( .A(\mult_22/ab[2][58] ), .B(
        \mult_22/CARRYB[1][58] ), .CI(\mult_22/n195 ), .CO(
        \mult_22/CARRYB[2][58] ), .S(\mult_22/SUMB[2][58] ) );
  FA_X1 \mult_22/S2_2_57  ( .A(\mult_22/ab[2][57] ), .B(\mult_22/n60 ), .CI(
        \mult_22/n194 ), .CO(\mult_22/CARRYB[2][57] ), .S(
        \mult_22/SUMB[2][57] ) );
  FA_X1 \mult_22/S2_2_55  ( .A(\mult_22/ab[2][55] ), .B(
        \mult_22/CARRYB[1][55] ), .CI(\mult_22/n322 ), .CO(
        \mult_22/CARRYB[2][55] ), .S(\mult_22/SUMB[2][55] ) );
  FA_X1 \mult_22/S2_2_54  ( .A(\mult_22/ab[2][54] ), .B(\mult_22/n324 ), .CI(
        \mult_22/SUMB[1][55] ), .CO(\mult_22/CARRYB[2][54] ), .S(
        \mult_22/SUMB[2][54] ) );
  FA_X1 \mult_22/S2_2_53  ( .A(\mult_22/ab[2][53] ), .B(\mult_22/n6 ), .CI(
        \mult_22/n66 ), .CO(\mult_22/CARRYB[2][53] ), .S(\mult_22/SUMB[2][53] ) );
  FA_X1 \mult_22/S2_2_52  ( .A(\mult_22/ab[2][52] ), .B(\mult_22/n7 ), .CI(
        \mult_22/n61 ), .CO(\mult_22/CARRYB[2][52] ), .S(\mult_22/SUMB[2][52] ) );
  FA_X1 \mult_22/S2_2_51  ( .A(\mult_22/ab[2][51] ), .B(\mult_22/n10 ), .CI(
        \mult_22/n62 ), .CO(\mult_22/CARRYB[2][51] ), .S(\mult_22/SUMB[2][51] ) );
  FA_X1 \mult_22/S2_2_50  ( .A(\mult_22/ab[2][50] ), .B(\mult_22/n8 ), .CI(
        \mult_22/n64 ), .CO(\mult_22/CARRYB[2][50] ), .S(\mult_22/SUMB[2][50] ) );
  FA_X1 \mult_22/S2_2_49  ( .A(\mult_22/ab[2][49] ), .B(\mult_22/n9 ), .CI(
        \mult_22/n63 ), .CO(\mult_22/CARRYB[2][49] ), .S(\mult_22/SUMB[2][49] ) );
  FA_X1 \mult_22/S2_2_48  ( .A(\mult_22/ab[2][48] ), .B(\mult_22/n67 ), .CI(
        \mult_22/n13 ), .CO(\mult_22/CARRYB[2][48] ), .S(\mult_22/SUMB[2][48] ) );
  FA_X1 \mult_22/S2_2_47  ( .A(\mult_22/ab[2][47] ), .B(\mult_22/n11 ), .CI(
        \mult_22/n90 ), .CO(\mult_22/CARRYB[2][47] ), .S(\mult_22/SUMB[2][47] ) );
  FA_X1 \mult_22/S2_2_46  ( .A(\mult_22/ab[2][46] ), .B(\mult_22/n5 ), .CI(
        \mult_22/n65 ), .CO(\mult_22/CARRYB[2][46] ), .S(\mult_22/SUMB[2][46] ) );
  FA_X1 \mult_22/S2_2_45  ( .A(\mult_22/ab[2][45] ), .B(\mult_22/n68 ), .CI(
        \mult_22/n12 ), .CO(\mult_22/CARRYB[2][45] ), .S(\mult_22/SUMB[2][45] ) );
  FA_X1 \mult_22/S2_2_44  ( .A(\mult_22/ab[2][44] ), .B(\mult_22/n22 ), .CI(
        \mult_22/n113 ), .CO(\mult_22/CARRYB[2][44] ), .S(
        \mult_22/SUMB[2][44] ) );
  FA_X1 \mult_22/S2_2_43  ( .A(\mult_22/ab[2][43] ), .B(\mult_22/n57 ), .CI(
        \mult_22/n91 ), .CO(\mult_22/CARRYB[2][43] ), .S(\mult_22/SUMB[2][43] ) );
  FA_X1 \mult_22/S2_2_42  ( .A(\mult_22/ab[2][42] ), .B(\mult_22/n23 ), .CI(
        \mult_22/n112 ), .CO(\mult_22/CARRYB[2][42] ), .S(
        \mult_22/SUMB[2][42] ) );
  FA_X1 \mult_22/S2_2_41  ( .A(\mult_22/ab[2][41] ), .B(\mult_22/n58 ), .CI(
        \mult_22/n92 ), .CO(\mult_22/CARRYB[2][41] ), .S(\mult_22/SUMB[2][41] ) );
  FA_X1 \mult_22/S2_2_40  ( .A(\mult_22/ab[2][40] ), .B(\mult_22/n14 ), .CI(
        \mult_22/n114 ), .CO(\mult_22/CARRYB[2][40] ), .S(
        \mult_22/SUMB[2][40] ) );
  FA_X1 \mult_22/S2_2_39  ( .A(\mult_22/ab[2][39] ), .B(\mult_22/n24 ), .CI(
        \mult_22/n69 ), .CO(\mult_22/CARRYB[2][39] ), .S(\mult_22/SUMB[2][39] ) );
  FA_X1 \mult_22/S2_2_38  ( .A(\mult_22/ab[2][38] ), .B(\mult_22/n25 ), .CI(
        \mult_22/n93 ), .CO(\mult_22/CARRYB[2][38] ), .S(\mult_22/SUMB[2][38] ) );
  FA_X1 \mult_22/S2_2_37  ( .A(\mult_22/ab[2][37] ), .B(\mult_22/n26 ), .CI(
        \mult_22/n94 ), .CO(\mult_22/CARRYB[2][37] ), .S(\mult_22/SUMB[2][37] ) );
  FA_X1 \mult_22/S2_2_36  ( .A(\mult_22/ab[2][36] ), .B(\mult_22/n27 ), .CI(
        \mult_22/n95 ), .CO(\mult_22/CARRYB[2][36] ), .S(\mult_22/SUMB[2][36] ) );
  FA_X1 \mult_22/S2_2_35  ( .A(\mult_22/ab[2][35] ), .B(\mult_22/n28 ), .CI(
        \mult_22/n96 ), .CO(\mult_22/CARRYB[2][35] ), .S(\mult_22/SUMB[2][35] ) );
  FA_X1 \mult_22/S2_2_34  ( .A(\mult_22/ab[2][34] ), .B(\mult_22/n29 ), .CI(
        \mult_22/n97 ), .CO(\mult_22/CARRYB[2][34] ), .S(\mult_22/SUMB[2][34] ) );
  FA_X1 \mult_22/S2_2_33  ( .A(\mult_22/ab[2][33] ), .B(\mult_22/n30 ), .CI(
        \mult_22/n98 ), .CO(\mult_22/CARRYB[2][33] ), .S(\mult_22/SUMB[2][33] ) );
  FA_X1 \mult_22/S2_2_32  ( .A(\mult_22/ab[2][32] ), .B(\mult_22/n31 ), .CI(
        \mult_22/n99 ), .CO(\mult_22/CARRYB[2][32] ), .S(\mult_22/SUMB[2][32] ) );
  FA_X1 \mult_22/S2_2_31  ( .A(\mult_22/ab[2][31] ), .B(\mult_22/n15 ), .CI(
        \mult_22/n100 ), .CO(\mult_22/CARRYB[2][31] ), .S(
        \mult_22/SUMB[2][31] ) );
  FA_X1 \mult_22/S2_2_30  ( .A(\mult_22/ab[2][30] ), .B(\mult_22/n32 ), .CI(
        \mult_22/n70 ), .CO(\mult_22/CARRYB[2][30] ), .S(\mult_22/SUMB[2][30] ) );
  FA_X1 \mult_22/S2_2_29  ( .A(\mult_22/ab[2][29] ), .B(\mult_22/n33 ), .CI(
        \mult_22/n101 ), .CO(\mult_22/CARRYB[2][29] ), .S(
        \mult_22/SUMB[2][29] ) );
  FA_X1 \mult_22/S2_2_28  ( .A(\mult_22/ab[2][28] ), .B(\mult_22/n34 ), .CI(
        \mult_22/n102 ), .CO(\mult_22/CARRYB[2][28] ), .S(
        \mult_22/SUMB[2][28] ) );
  FA_X1 \mult_22/S2_2_27  ( .A(\mult_22/ab[2][27] ), .B(\mult_22/n35 ), .CI(
        \mult_22/n103 ), .CO(\mult_22/CARRYB[2][27] ), .S(
        \mult_22/SUMB[2][27] ) );
  FA_X1 \mult_22/S2_2_26  ( .A(\mult_22/ab[2][26] ), .B(\mult_22/n36 ), .CI(
        \mult_22/n104 ), .CO(\mult_22/CARRYB[2][26] ), .S(
        \mult_22/SUMB[2][26] ) );
  FA_X1 \mult_22/S2_2_25  ( .A(\mult_22/ab[2][25] ), .B(\mult_22/n37 ), .CI(
        \mult_22/n105 ), .CO(\mult_22/CARRYB[2][25] ), .S(
        \mult_22/SUMB[2][25] ) );
  FA_X1 \mult_22/S2_2_24  ( .A(\mult_22/ab[2][24] ), .B(\mult_22/n38 ), .CI(
        \mult_22/n106 ), .CO(\mult_22/CARRYB[2][24] ), .S(
        \mult_22/SUMB[2][24] ) );
  FA_X1 \mult_22/S2_2_23  ( .A(\mult_22/ab[2][23] ), .B(\mult_22/n39 ), .CI(
        \mult_22/n107 ), .CO(\mult_22/CARRYB[2][23] ), .S(
        \mult_22/SUMB[2][23] ) );
  FA_X1 \mult_22/S2_2_22  ( .A(\mult_22/ab[2][22] ), .B(\mult_22/n40 ), .CI(
        \mult_22/n76 ), .CO(\mult_22/CARRYB[2][22] ), .S(\mult_22/SUMB[2][22] ) );
  FA_X1 \mult_22/S2_2_21  ( .A(\mult_22/ab[2][21] ), .B(\mult_22/n41 ), .CI(
        \mult_22/n77 ), .CO(\mult_22/CARRYB[2][21] ), .S(\mult_22/SUMB[2][21] ) );
  FA_X1 \mult_22/S2_2_20  ( .A(\mult_22/ab[2][20] ), .B(\mult_22/n42 ), .CI(
        \mult_22/n78 ), .CO(\mult_22/CARRYB[2][20] ), .S(\mult_22/SUMB[2][20] ) );
  FA_X1 \mult_22/S2_2_19  ( .A(\mult_22/ab[2][19] ), .B(\mult_22/n16 ), .CI(
        \mult_22/n79 ), .CO(\mult_22/CARRYB[2][19] ), .S(\mult_22/SUMB[2][19] ) );
  FA_X1 \mult_22/S2_2_18  ( .A(\mult_22/ab[2][18] ), .B(\mult_22/n43 ), .CI(
        \mult_22/n71 ), .CO(\mult_22/CARRYB[2][18] ), .S(\mult_22/SUMB[2][18] ) );
  FA_X1 \mult_22/S2_2_17  ( .A(\mult_22/ab[2][17] ), .B(\mult_22/n44 ), .CI(
        \mult_22/n80 ), .CO(\mult_22/CARRYB[2][17] ), .S(\mult_22/SUMB[2][17] ) );
  FA_X1 \mult_22/S2_2_16  ( .A(\mult_22/ab[2][16] ), .B(\mult_22/n45 ), .CI(
        \mult_22/n81 ), .CO(\mult_22/CARRYB[2][16] ), .S(\mult_22/SUMB[2][16] ) );
  FA_X1 \mult_22/S2_2_15  ( .A(\mult_22/ab[2][15] ), .B(\mult_22/n46 ), .CI(
        \mult_22/n82 ), .CO(\mult_22/CARRYB[2][15] ), .S(\mult_22/SUMB[2][15] ) );
  FA_X1 \mult_22/S2_2_14  ( .A(\mult_22/ab[2][14] ), .B(\mult_22/n17 ), .CI(
        \mult_22/n83 ), .CO(\mult_22/CARRYB[2][14] ), .S(\mult_22/SUMB[2][14] ) );
  FA_X1 \mult_22/S2_2_13  ( .A(\mult_22/ab[2][13] ), .B(\mult_22/n47 ), .CI(
        \mult_22/n72 ), .CO(\mult_22/CARRYB[2][13] ), .S(\mult_22/SUMB[2][13] ) );
  FA_X1 \mult_22/S2_2_12  ( .A(\mult_22/ab[2][12] ), .B(\mult_22/n48 ), .CI(
        \mult_22/n84 ), .CO(\mult_22/CARRYB[2][12] ), .S(\mult_22/SUMB[2][12] ) );
  FA_X1 \mult_22/S2_2_11  ( .A(\mult_22/ab[2][11] ), .B(\mult_22/n49 ), .CI(
        \mult_22/n108 ), .CO(\mult_22/CARRYB[2][11] ), .S(
        \mult_22/SUMB[2][11] ) );
  FA_X1 \mult_22/S2_2_10  ( .A(\mult_22/ab[2][10] ), .B(\mult_22/n50 ), .CI(
        \mult_22/n109 ), .CO(\mult_22/CARRYB[2][10] ), .S(
        \mult_22/SUMB[2][10] ) );
  FA_X1 \mult_22/S2_2_9  ( .A(\mult_22/ab[2][9] ), .B(\mult_22/n51 ), .CI(
        \mult_22/n110 ), .CO(\mult_22/CARRYB[2][9] ), .S(\mult_22/SUMB[2][9] )
         );
  FA_X1 \mult_22/S2_2_8  ( .A(\mult_22/ab[2][8] ), .B(\mult_22/n52 ), .CI(
        \mult_22/n85 ), .CO(\mult_22/CARRYB[2][8] ), .S(\mult_22/SUMB[2][8] )
         );
  FA_X1 \mult_22/S2_2_7  ( .A(\mult_22/ab[2][7] ), .B(\mult_22/n53 ), .CI(
        \mult_22/n86 ), .CO(\mult_22/CARRYB[2][7] ), .S(\mult_22/SUMB[2][7] )
         );
  FA_X1 \mult_22/S2_2_6  ( .A(\mult_22/ab[2][6] ), .B(\mult_22/n18 ), .CI(
        \mult_22/n87 ), .CO(\mult_22/CARRYB[2][6] ), .S(\mult_22/SUMB[2][6] )
         );
  FA_X1 \mult_22/S2_2_5  ( .A(\mult_22/ab[2][5] ), .B(\mult_22/n54 ), .CI(
        \mult_22/n73 ), .CO(\mult_22/CARRYB[2][5] ), .S(\mult_22/SUMB[2][5] )
         );
  FA_X1 \mult_22/S2_2_4  ( .A(\mult_22/ab[2][4] ), .B(\mult_22/n55 ), .CI(
        \mult_22/n88 ), .CO(\mult_22/CARRYB[2][4] ), .S(\mult_22/SUMB[2][4] )
         );
  FA_X1 \mult_22/S2_2_3  ( .A(\mult_22/ab[2][3] ), .B(\mult_22/n19 ), .CI(
        \mult_22/n111 ), .CO(\mult_22/CARRYB[2][3] ), .S(\mult_22/SUMB[2][3] )
         );
  FA_X1 \mult_22/S2_2_2  ( .A(\mult_22/ab[2][2] ), .B(\mult_22/n20 ), .CI(
        \mult_22/n74 ), .CO(\mult_22/CARRYB[2][2] ), .S(\mult_22/SUMB[2][2] )
         );
  FA_X1 \mult_22/S2_2_1  ( .A(\mult_22/ab[2][1] ), .B(\mult_22/n56 ), .CI(
        \mult_22/n75 ), .CO(\mult_22/CARRYB[2][1] ), .S(\mult_22/SUMB[2][1] )
         );
  FA_X1 \mult_22/S1_2_0  ( .A(\mult_22/ab[2][0] ), .B(\mult_22/n21 ), .CI(
        \mult_22/n89 ), .CO(\mult_22/CARRYB[2][0] ), .S(N130) );
  FA_X1 \mult_22/S2_3_60  ( .A(\mult_22/ab[3][60] ), .B(
        \mult_22/CARRYB[2][60] ), .CI(\mult_22/SUMB[2][61] ), .CO(
        \mult_22/CARRYB[3][60] ), .S(\mult_22/SUMB[3][60] ) );
  FA_X1 \mult_22/S2_3_59  ( .A(\mult_22/CARRYB[2][59] ), .B(
        \mult_22/ab[3][59] ), .CI(\mult_22/SUMB[2][60] ), .CO(
        \mult_22/CARRYB[3][59] ), .S(\mult_22/SUMB[3][59] ) );
  FA_X1 \mult_22/S2_3_58  ( .A(\mult_22/ab[3][58] ), .B(
        \mult_22/CARRYB[2][58] ), .CI(\mult_22/SUMB[2][59] ), .CO(
        \mult_22/CARRYB[3][58] ), .S(\mult_22/SUMB[3][58] ) );
  FA_X1 \mult_22/S2_3_57  ( .A(\mult_22/ab[3][57] ), .B(
        \mult_22/CARRYB[2][57] ), .CI(\mult_22/SUMB[2][58] ), .CO(
        \mult_22/CARRYB[3][57] ), .S(\mult_22/SUMB[3][57] ) );
  FA_X1 \mult_22/S2_3_54  ( .A(\mult_22/ab[3][54] ), .B(
        \mult_22/CARRYB[2][54] ), .CI(\mult_22/SUMB[2][55] ), .CO(
        \mult_22/CARRYB[3][54] ), .S(\mult_22/SUMB[3][54] ) );
  FA_X1 \mult_22/S2_3_53  ( .A(\mult_22/ab[3][53] ), .B(
        \mult_22/CARRYB[2][53] ), .CI(\mult_22/SUMB[2][54] ), .CO(
        \mult_22/CARRYB[3][53] ), .S(\mult_22/SUMB[3][53] ) );
  FA_X1 \mult_22/S2_3_52  ( .A(\mult_22/ab[3][52] ), .B(
        \mult_22/CARRYB[2][52] ), .CI(\mult_22/SUMB[2][53] ), .CO(
        \mult_22/CARRYB[3][52] ), .S(\mult_22/SUMB[3][52] ) );
  FA_X1 \mult_22/S2_3_51  ( .A(\mult_22/ab[3][51] ), .B(
        \mult_22/CARRYB[2][51] ), .CI(\mult_22/SUMB[2][52] ), .CO(
        \mult_22/CARRYB[3][51] ), .S(\mult_22/SUMB[3][51] ) );
  FA_X1 \mult_22/S2_3_50  ( .A(\mult_22/ab[3][50] ), .B(
        \mult_22/CARRYB[2][50] ), .CI(\mult_22/SUMB[2][51] ), .CO(
        \mult_22/CARRYB[3][50] ), .S(\mult_22/SUMB[3][50] ) );
  FA_X1 \mult_22/S2_3_49  ( .A(\mult_22/ab[3][49] ), .B(
        \mult_22/CARRYB[2][49] ), .CI(\mult_22/SUMB[2][50] ), .CO(
        \mult_22/CARRYB[3][49] ), .S(\mult_22/SUMB[3][49] ) );
  FA_X1 \mult_22/S2_3_48  ( .A(\mult_22/ab[3][48] ), .B(
        \mult_22/CARRYB[2][48] ), .CI(\mult_22/SUMB[2][49] ), .CO(
        \mult_22/CARRYB[3][48] ), .S(\mult_22/SUMB[3][48] ) );
  FA_X1 \mult_22/S2_3_47  ( .A(\mult_22/ab[3][47] ), .B(
        \mult_22/CARRYB[2][47] ), .CI(\mult_22/SUMB[2][48] ), .CO(
        \mult_22/CARRYB[3][47] ), .S(\mult_22/SUMB[3][47] ) );
  FA_X1 \mult_22/S2_3_46  ( .A(\mult_22/ab[3][46] ), .B(
        \mult_22/CARRYB[2][46] ), .CI(\mult_22/SUMB[2][47] ), .CO(
        \mult_22/CARRYB[3][46] ), .S(\mult_22/SUMB[3][46] ) );
  FA_X1 \mult_22/S2_3_45  ( .A(\mult_22/ab[3][45] ), .B(
        \mult_22/CARRYB[2][45] ), .CI(\mult_22/SUMB[2][46] ), .CO(
        \mult_22/CARRYB[3][45] ), .S(\mult_22/SUMB[3][45] ) );
  FA_X1 \mult_22/S2_3_44  ( .A(\mult_22/ab[3][44] ), .B(
        \mult_22/CARRYB[2][44] ), .CI(\mult_22/SUMB[2][45] ), .CO(
        \mult_22/CARRYB[3][44] ), .S(\mult_22/SUMB[3][44] ) );
  FA_X1 \mult_22/S2_3_43  ( .A(\mult_22/ab[3][43] ), .B(
        \mult_22/CARRYB[2][43] ), .CI(\mult_22/SUMB[2][44] ), .CO(
        \mult_22/CARRYB[3][43] ), .S(\mult_22/SUMB[3][43] ) );
  FA_X1 \mult_22/S2_3_42  ( .A(\mult_22/ab[3][42] ), .B(
        \mult_22/CARRYB[2][42] ), .CI(\mult_22/SUMB[2][43] ), .CO(
        \mult_22/CARRYB[3][42] ), .S(\mult_22/SUMB[3][42] ) );
  FA_X1 \mult_22/S2_3_41  ( .A(\mult_22/ab[3][41] ), .B(
        \mult_22/CARRYB[2][41] ), .CI(\mult_22/SUMB[2][42] ), .CO(
        \mult_22/CARRYB[3][41] ), .S(\mult_22/SUMB[3][41] ) );
  FA_X1 \mult_22/S2_3_40  ( .A(\mult_22/ab[3][40] ), .B(
        \mult_22/CARRYB[2][40] ), .CI(\mult_22/SUMB[2][41] ), .CO(
        \mult_22/CARRYB[3][40] ), .S(\mult_22/SUMB[3][40] ) );
  FA_X1 \mult_22/S2_3_39  ( .A(\mult_22/ab[3][39] ), .B(
        \mult_22/CARRYB[2][39] ), .CI(\mult_22/SUMB[2][40] ), .CO(
        \mult_22/CARRYB[3][39] ), .S(\mult_22/SUMB[3][39] ) );
  FA_X1 \mult_22/S2_3_38  ( .A(\mult_22/ab[3][38] ), .B(
        \mult_22/CARRYB[2][38] ), .CI(\mult_22/SUMB[2][39] ), .CO(
        \mult_22/CARRYB[3][38] ), .S(\mult_22/SUMB[3][38] ) );
  FA_X1 \mult_22/S2_3_37  ( .A(\mult_22/ab[3][37] ), .B(
        \mult_22/CARRYB[2][37] ), .CI(\mult_22/SUMB[2][38] ), .CO(
        \mult_22/CARRYB[3][37] ), .S(\mult_22/SUMB[3][37] ) );
  FA_X1 \mult_22/S2_3_36  ( .A(\mult_22/ab[3][36] ), .B(
        \mult_22/CARRYB[2][36] ), .CI(\mult_22/SUMB[2][37] ), .CO(
        \mult_22/CARRYB[3][36] ), .S(\mult_22/SUMB[3][36] ) );
  FA_X1 \mult_22/S2_3_35  ( .A(\mult_22/ab[3][35] ), .B(
        \mult_22/CARRYB[2][35] ), .CI(\mult_22/SUMB[2][36] ), .CO(
        \mult_22/CARRYB[3][35] ), .S(\mult_22/SUMB[3][35] ) );
  FA_X1 \mult_22/S2_3_34  ( .A(\mult_22/ab[3][34] ), .B(
        \mult_22/CARRYB[2][34] ), .CI(\mult_22/SUMB[2][35] ), .CO(
        \mult_22/CARRYB[3][34] ), .S(\mult_22/SUMB[3][34] ) );
  FA_X1 \mult_22/S2_3_33  ( .A(\mult_22/ab[3][33] ), .B(
        \mult_22/CARRYB[2][33] ), .CI(\mult_22/SUMB[2][34] ), .CO(
        \mult_22/CARRYB[3][33] ), .S(\mult_22/SUMB[3][33] ) );
  FA_X1 \mult_22/S2_3_32  ( .A(\mult_22/ab[3][32] ), .B(
        \mult_22/CARRYB[2][32] ), .CI(\mult_22/SUMB[2][33] ), .CO(
        \mult_22/CARRYB[3][32] ), .S(\mult_22/SUMB[3][32] ) );
  FA_X1 \mult_22/S2_3_31  ( .A(\mult_22/ab[3][31] ), .B(
        \mult_22/CARRYB[2][31] ), .CI(\mult_22/SUMB[2][32] ), .CO(
        \mult_22/CARRYB[3][31] ), .S(\mult_22/SUMB[3][31] ) );
  FA_X1 \mult_22/S2_3_30  ( .A(\mult_22/ab[3][30] ), .B(
        \mult_22/CARRYB[2][30] ), .CI(\mult_22/SUMB[2][31] ), .CO(
        \mult_22/CARRYB[3][30] ), .S(\mult_22/SUMB[3][30] ) );
  FA_X1 \mult_22/S2_3_29  ( .A(\mult_22/ab[3][29] ), .B(
        \mult_22/CARRYB[2][29] ), .CI(\mult_22/SUMB[2][30] ), .CO(
        \mult_22/CARRYB[3][29] ), .S(\mult_22/SUMB[3][29] ) );
  FA_X1 \mult_22/S2_3_28  ( .A(\mult_22/ab[3][28] ), .B(
        \mult_22/CARRYB[2][28] ), .CI(\mult_22/SUMB[2][29] ), .CO(
        \mult_22/CARRYB[3][28] ), .S(\mult_22/SUMB[3][28] ) );
  FA_X1 \mult_22/S2_3_27  ( .A(\mult_22/ab[3][27] ), .B(
        \mult_22/CARRYB[2][27] ), .CI(\mult_22/SUMB[2][28] ), .CO(
        \mult_22/CARRYB[3][27] ), .S(\mult_22/SUMB[3][27] ) );
  FA_X1 \mult_22/S2_3_26  ( .A(\mult_22/ab[3][26] ), .B(
        \mult_22/CARRYB[2][26] ), .CI(\mult_22/SUMB[2][27] ), .CO(
        \mult_22/CARRYB[3][26] ), .S(\mult_22/SUMB[3][26] ) );
  FA_X1 \mult_22/S2_3_25  ( .A(\mult_22/ab[3][25] ), .B(
        \mult_22/CARRYB[2][25] ), .CI(\mult_22/SUMB[2][26] ), .CO(
        \mult_22/CARRYB[3][25] ), .S(\mult_22/SUMB[3][25] ) );
  FA_X1 \mult_22/S2_3_24  ( .A(\mult_22/ab[3][24] ), .B(
        \mult_22/CARRYB[2][24] ), .CI(\mult_22/SUMB[2][25] ), .CO(
        \mult_22/CARRYB[3][24] ), .S(\mult_22/SUMB[3][24] ) );
  FA_X1 \mult_22/S2_3_23  ( .A(\mult_22/ab[3][23] ), .B(
        \mult_22/CARRYB[2][23] ), .CI(\mult_22/SUMB[2][24] ), .CO(
        \mult_22/CARRYB[3][23] ), .S(\mult_22/SUMB[3][23] ) );
  FA_X1 \mult_22/S2_3_22  ( .A(\mult_22/ab[3][22] ), .B(
        \mult_22/CARRYB[2][22] ), .CI(\mult_22/SUMB[2][23] ), .CO(
        \mult_22/CARRYB[3][22] ), .S(\mult_22/SUMB[3][22] ) );
  FA_X1 \mult_22/S2_3_21  ( .A(\mult_22/ab[3][21] ), .B(
        \mult_22/CARRYB[2][21] ), .CI(\mult_22/SUMB[2][22] ), .CO(
        \mult_22/CARRYB[3][21] ), .S(\mult_22/SUMB[3][21] ) );
  FA_X1 \mult_22/S2_3_20  ( .A(\mult_22/ab[3][20] ), .B(
        \mult_22/CARRYB[2][20] ), .CI(\mult_22/SUMB[2][21] ), .CO(
        \mult_22/CARRYB[3][20] ), .S(\mult_22/SUMB[3][20] ) );
  FA_X1 \mult_22/S2_3_19  ( .A(\mult_22/ab[3][19] ), .B(
        \mult_22/CARRYB[2][19] ), .CI(\mult_22/SUMB[2][20] ), .CO(
        \mult_22/CARRYB[3][19] ), .S(\mult_22/SUMB[3][19] ) );
  FA_X1 \mult_22/S2_3_18  ( .A(\mult_22/ab[3][18] ), .B(
        \mult_22/CARRYB[2][18] ), .CI(\mult_22/SUMB[2][19] ), .CO(
        \mult_22/CARRYB[3][18] ), .S(\mult_22/SUMB[3][18] ) );
  FA_X1 \mult_22/S2_3_17  ( .A(\mult_22/ab[3][17] ), .B(
        \mult_22/CARRYB[2][17] ), .CI(\mult_22/SUMB[2][18] ), .CO(
        \mult_22/CARRYB[3][17] ), .S(\mult_22/SUMB[3][17] ) );
  FA_X1 \mult_22/S2_3_16  ( .A(\mult_22/ab[3][16] ), .B(
        \mult_22/CARRYB[2][16] ), .CI(\mult_22/SUMB[2][17] ), .CO(
        \mult_22/CARRYB[3][16] ), .S(\mult_22/SUMB[3][16] ) );
  FA_X1 \mult_22/S2_3_15  ( .A(\mult_22/ab[3][15] ), .B(
        \mult_22/CARRYB[2][15] ), .CI(\mult_22/SUMB[2][16] ), .CO(
        \mult_22/CARRYB[3][15] ), .S(\mult_22/SUMB[3][15] ) );
  FA_X1 \mult_22/S2_3_14  ( .A(\mult_22/ab[3][14] ), .B(
        \mult_22/CARRYB[2][14] ), .CI(\mult_22/SUMB[2][15] ), .CO(
        \mult_22/CARRYB[3][14] ), .S(\mult_22/SUMB[3][14] ) );
  FA_X1 \mult_22/S2_3_13  ( .A(\mult_22/ab[3][13] ), .B(
        \mult_22/CARRYB[2][13] ), .CI(\mult_22/SUMB[2][14] ), .CO(
        \mult_22/CARRYB[3][13] ), .S(\mult_22/SUMB[3][13] ) );
  FA_X1 \mult_22/S2_3_12  ( .A(\mult_22/ab[3][12] ), .B(
        \mult_22/CARRYB[2][12] ), .CI(\mult_22/SUMB[2][13] ), .CO(
        \mult_22/CARRYB[3][12] ), .S(\mult_22/SUMB[3][12] ) );
  FA_X1 \mult_22/S2_3_11  ( .A(\mult_22/ab[3][11] ), .B(
        \mult_22/CARRYB[2][11] ), .CI(\mult_22/SUMB[2][12] ), .CO(
        \mult_22/CARRYB[3][11] ), .S(\mult_22/SUMB[3][11] ) );
  FA_X1 \mult_22/S2_3_10  ( .A(\mult_22/ab[3][10] ), .B(
        \mult_22/CARRYB[2][10] ), .CI(\mult_22/SUMB[2][11] ), .CO(
        \mult_22/CARRYB[3][10] ), .S(\mult_22/SUMB[3][10] ) );
  FA_X1 \mult_22/S2_3_9  ( .A(\mult_22/ab[3][9] ), .B(\mult_22/CARRYB[2][9] ), 
        .CI(\mult_22/SUMB[2][10] ), .CO(\mult_22/CARRYB[3][9] ), .S(
        \mult_22/SUMB[3][9] ) );
  FA_X1 \mult_22/S2_3_8  ( .A(\mult_22/ab[3][8] ), .B(\mult_22/CARRYB[2][8] ), 
        .CI(\mult_22/SUMB[2][9] ), .CO(\mult_22/CARRYB[3][8] ), .S(
        \mult_22/SUMB[3][8] ) );
  FA_X1 \mult_22/S2_3_7  ( .A(\mult_22/ab[3][7] ), .B(\mult_22/CARRYB[2][7] ), 
        .CI(\mult_22/SUMB[2][8] ), .CO(\mult_22/CARRYB[3][7] ), .S(
        \mult_22/SUMB[3][7] ) );
  FA_X1 \mult_22/S2_3_6  ( .A(\mult_22/ab[3][6] ), .B(\mult_22/CARRYB[2][6] ), 
        .CI(\mult_22/SUMB[2][7] ), .CO(\mult_22/CARRYB[3][6] ), .S(
        \mult_22/SUMB[3][6] ) );
  FA_X1 \mult_22/S2_3_5  ( .A(\mult_22/ab[3][5] ), .B(\mult_22/CARRYB[2][5] ), 
        .CI(\mult_22/SUMB[2][6] ), .CO(\mult_22/CARRYB[3][5] ), .S(
        \mult_22/SUMB[3][5] ) );
  FA_X1 \mult_22/S2_3_4  ( .A(\mult_22/ab[3][4] ), .B(\mult_22/CARRYB[2][4] ), 
        .CI(\mult_22/SUMB[2][5] ), .CO(\mult_22/CARRYB[3][4] ), .S(
        \mult_22/SUMB[3][4] ) );
  FA_X1 \mult_22/S2_3_3  ( .A(\mult_22/ab[3][3] ), .B(\mult_22/CARRYB[2][3] ), 
        .CI(\mult_22/SUMB[2][4] ), .CO(\mult_22/CARRYB[3][3] ), .S(
        \mult_22/SUMB[3][3] ) );
  FA_X1 \mult_22/S2_3_2  ( .A(\mult_22/ab[3][2] ), .B(\mult_22/CARRYB[2][2] ), 
        .CI(\mult_22/SUMB[2][3] ), .CO(\mult_22/CARRYB[3][2] ), .S(
        \mult_22/SUMB[3][2] ) );
  FA_X1 \mult_22/S2_3_1  ( .A(\mult_22/ab[3][1] ), .B(\mult_22/CARRYB[2][1] ), 
        .CI(\mult_22/SUMB[2][2] ), .CO(\mult_22/CARRYB[3][1] ), .S(
        \mult_22/SUMB[3][1] ) );
  FA_X1 \mult_22/S1_3_0  ( .A(\mult_22/ab[3][0] ), .B(\mult_22/CARRYB[2][0] ), 
        .CI(\mult_22/SUMB[2][1] ), .CO(\mult_22/CARRYB[3][0] ), .S(N131) );
  FA_X1 \mult_22/S2_4_59  ( .A(\mult_22/ab[4][59] ), .B(
        \mult_22/CARRYB[3][59] ), .CI(\mult_22/SUMB[3][60] ), .CO(
        \mult_22/CARRYB[4][59] ), .S(\mult_22/SUMB[4][59] ) );
  FA_X1 \mult_22/S2_4_58  ( .A(\mult_22/ab[4][58] ), .B(
        \mult_22/CARRYB[3][58] ), .CI(\mult_22/SUMB[3][59] ), .CO(
        \mult_22/CARRYB[4][58] ), .S(\mult_22/SUMB[4][58] ) );
  FA_X1 \mult_22/S2_4_57  ( .A(\mult_22/CARRYB[3][57] ), .B(
        \mult_22/ab[4][57] ), .CI(\mult_22/SUMB[3][58] ), .CO(
        \mult_22/CARRYB[4][57] ), .S(\mult_22/SUMB[4][57] ) );
  FA_X1 \mult_22/S2_4_56  ( .A(\mult_22/ab[4][56] ), .B(
        \mult_22/CARRYB[3][56] ), .CI(\mult_22/SUMB[3][57] ), .CO(
        \mult_22/CARRYB[4][56] ), .S(\mult_22/SUMB[4][56] ) );
  FA_X1 \mult_22/S2_4_54  ( .A(\mult_22/ab[4][54] ), .B(
        \mult_22/CARRYB[3][54] ), .CI(\mult_22/SUMB[3][55] ), .CO(
        \mult_22/CARRYB[4][54] ), .S(\mult_22/SUMB[4][54] ) );
  FA_X1 \mult_22/S2_4_53  ( .A(\mult_22/ab[4][53] ), .B(
        \mult_22/CARRYB[3][53] ), .CI(\mult_22/SUMB[3][54] ), .CO(
        \mult_22/CARRYB[4][53] ), .S(\mult_22/SUMB[4][53] ) );
  FA_X1 \mult_22/S2_4_51  ( .A(\mult_22/ab[4][51] ), .B(
        \mult_22/CARRYB[3][51] ), .CI(\mult_22/SUMB[3][52] ), .CO(
        \mult_22/CARRYB[4][51] ), .S(\mult_22/SUMB[4][51] ) );
  FA_X1 \mult_22/S2_4_50  ( .A(\mult_22/ab[4][50] ), .B(
        \mult_22/CARRYB[3][50] ), .CI(\mult_22/SUMB[3][51] ), .CO(
        \mult_22/CARRYB[4][50] ), .S(\mult_22/SUMB[4][50] ) );
  FA_X1 \mult_22/S2_4_49  ( .A(\mult_22/ab[4][49] ), .B(
        \mult_22/CARRYB[3][49] ), .CI(\mult_22/SUMB[3][50] ), .CO(
        \mult_22/CARRYB[4][49] ), .S(\mult_22/SUMB[4][49] ) );
  FA_X1 \mult_22/S2_4_48  ( .A(\mult_22/ab[4][48] ), .B(
        \mult_22/CARRYB[3][48] ), .CI(\mult_22/SUMB[3][49] ), .CO(
        \mult_22/CARRYB[4][48] ), .S(\mult_22/SUMB[4][48] ) );
  FA_X1 \mult_22/S2_4_47  ( .A(\mult_22/ab[4][47] ), .B(
        \mult_22/CARRYB[3][47] ), .CI(\mult_22/SUMB[3][48] ), .CO(
        \mult_22/CARRYB[4][47] ), .S(\mult_22/SUMB[4][47] ) );
  FA_X1 \mult_22/S2_4_46  ( .A(\mult_22/ab[4][46] ), .B(
        \mult_22/CARRYB[3][46] ), .CI(\mult_22/SUMB[3][47] ), .CO(
        \mult_22/CARRYB[4][46] ), .S(\mult_22/SUMB[4][46] ) );
  FA_X1 \mult_22/S2_4_45  ( .A(\mult_22/ab[4][45] ), .B(
        \mult_22/CARRYB[3][45] ), .CI(\mult_22/SUMB[3][46] ), .CO(
        \mult_22/CARRYB[4][45] ), .S(\mult_22/SUMB[4][45] ) );
  FA_X1 \mult_22/S2_4_44  ( .A(\mult_22/ab[4][44] ), .B(
        \mult_22/CARRYB[3][44] ), .CI(\mult_22/SUMB[3][45] ), .CO(
        \mult_22/CARRYB[4][44] ), .S(\mult_22/SUMB[4][44] ) );
  FA_X1 \mult_22/S2_4_43  ( .A(\mult_22/ab[4][43] ), .B(
        \mult_22/CARRYB[3][43] ), .CI(\mult_22/SUMB[3][44] ), .CO(
        \mult_22/CARRYB[4][43] ), .S(\mult_22/SUMB[4][43] ) );
  FA_X1 \mult_22/S2_4_42  ( .A(\mult_22/ab[4][42] ), .B(
        \mult_22/CARRYB[3][42] ), .CI(\mult_22/SUMB[3][43] ), .CO(
        \mult_22/CARRYB[4][42] ), .S(\mult_22/SUMB[4][42] ) );
  FA_X1 \mult_22/S2_4_41  ( .A(\mult_22/ab[4][41] ), .B(
        \mult_22/CARRYB[3][41] ), .CI(\mult_22/SUMB[3][42] ), .CO(
        \mult_22/CARRYB[4][41] ), .S(\mult_22/SUMB[4][41] ) );
  FA_X1 \mult_22/S2_4_40  ( .A(\mult_22/ab[4][40] ), .B(
        \mult_22/CARRYB[3][40] ), .CI(\mult_22/SUMB[3][41] ), .CO(
        \mult_22/CARRYB[4][40] ), .S(\mult_22/SUMB[4][40] ) );
  FA_X1 \mult_22/S2_4_39  ( .A(\mult_22/ab[4][39] ), .B(
        \mult_22/CARRYB[3][39] ), .CI(\mult_22/SUMB[3][40] ), .CO(
        \mult_22/CARRYB[4][39] ), .S(\mult_22/SUMB[4][39] ) );
  FA_X1 \mult_22/S2_4_38  ( .A(\mult_22/ab[4][38] ), .B(
        \mult_22/CARRYB[3][38] ), .CI(\mult_22/SUMB[3][39] ), .CO(
        \mult_22/CARRYB[4][38] ), .S(\mult_22/SUMB[4][38] ) );
  FA_X1 \mult_22/S2_4_37  ( .A(\mult_22/ab[4][37] ), .B(
        \mult_22/CARRYB[3][37] ), .CI(\mult_22/SUMB[3][38] ), .CO(
        \mult_22/CARRYB[4][37] ), .S(\mult_22/SUMB[4][37] ) );
  FA_X1 \mult_22/S2_4_36  ( .A(\mult_22/ab[4][36] ), .B(
        \mult_22/CARRYB[3][36] ), .CI(\mult_22/SUMB[3][37] ), .CO(
        \mult_22/CARRYB[4][36] ), .S(\mult_22/SUMB[4][36] ) );
  FA_X1 \mult_22/S2_4_35  ( .A(\mult_22/ab[4][35] ), .B(
        \mult_22/CARRYB[3][35] ), .CI(\mult_22/SUMB[3][36] ), .CO(
        \mult_22/CARRYB[4][35] ), .S(\mult_22/SUMB[4][35] ) );
  FA_X1 \mult_22/S2_4_34  ( .A(\mult_22/ab[4][34] ), .B(
        \mult_22/CARRYB[3][34] ), .CI(\mult_22/SUMB[3][35] ), .CO(
        \mult_22/CARRYB[4][34] ), .S(\mult_22/SUMB[4][34] ) );
  FA_X1 \mult_22/S2_4_33  ( .A(\mult_22/ab[4][33] ), .B(
        \mult_22/CARRYB[3][33] ), .CI(\mult_22/SUMB[3][34] ), .CO(
        \mult_22/CARRYB[4][33] ), .S(\mult_22/SUMB[4][33] ) );
  FA_X1 \mult_22/S2_4_32  ( .A(\mult_22/ab[4][32] ), .B(
        \mult_22/CARRYB[3][32] ), .CI(\mult_22/SUMB[3][33] ), .CO(
        \mult_22/CARRYB[4][32] ), .S(\mult_22/SUMB[4][32] ) );
  FA_X1 \mult_22/S2_4_31  ( .A(\mult_22/ab[4][31] ), .B(
        \mult_22/CARRYB[3][31] ), .CI(\mult_22/SUMB[3][32] ), .CO(
        \mult_22/CARRYB[4][31] ), .S(\mult_22/SUMB[4][31] ) );
  FA_X1 \mult_22/S2_4_30  ( .A(\mult_22/ab[4][30] ), .B(
        \mult_22/CARRYB[3][30] ), .CI(\mult_22/SUMB[3][31] ), .CO(
        \mult_22/CARRYB[4][30] ), .S(\mult_22/SUMB[4][30] ) );
  FA_X1 \mult_22/S2_4_29  ( .A(\mult_22/ab[4][29] ), .B(
        \mult_22/CARRYB[3][29] ), .CI(\mult_22/SUMB[3][30] ), .CO(
        \mult_22/CARRYB[4][29] ), .S(\mult_22/SUMB[4][29] ) );
  FA_X1 \mult_22/S2_4_28  ( .A(\mult_22/ab[4][28] ), .B(
        \mult_22/CARRYB[3][28] ), .CI(\mult_22/SUMB[3][29] ), .CO(
        \mult_22/CARRYB[4][28] ), .S(\mult_22/SUMB[4][28] ) );
  FA_X1 \mult_22/S2_4_27  ( .A(\mult_22/ab[4][27] ), .B(
        \mult_22/CARRYB[3][27] ), .CI(\mult_22/SUMB[3][28] ), .CO(
        \mult_22/CARRYB[4][27] ), .S(\mult_22/SUMB[4][27] ) );
  FA_X1 \mult_22/S2_4_26  ( .A(\mult_22/ab[4][26] ), .B(
        \mult_22/CARRYB[3][26] ), .CI(\mult_22/SUMB[3][27] ), .CO(
        \mult_22/CARRYB[4][26] ), .S(\mult_22/SUMB[4][26] ) );
  FA_X1 \mult_22/S2_4_25  ( .A(\mult_22/ab[4][25] ), .B(
        \mult_22/CARRYB[3][25] ), .CI(\mult_22/SUMB[3][26] ), .CO(
        \mult_22/CARRYB[4][25] ), .S(\mult_22/SUMB[4][25] ) );
  FA_X1 \mult_22/S2_4_24  ( .A(\mult_22/ab[4][24] ), .B(
        \mult_22/CARRYB[3][24] ), .CI(\mult_22/SUMB[3][25] ), .CO(
        \mult_22/CARRYB[4][24] ), .S(\mult_22/SUMB[4][24] ) );
  FA_X1 \mult_22/S2_4_23  ( .A(\mult_22/ab[4][23] ), .B(
        \mult_22/CARRYB[3][23] ), .CI(\mult_22/SUMB[3][24] ), .CO(
        \mult_22/CARRYB[4][23] ), .S(\mult_22/SUMB[4][23] ) );
  FA_X1 \mult_22/S2_4_22  ( .A(\mult_22/ab[4][22] ), .B(
        \mult_22/CARRYB[3][22] ), .CI(\mult_22/SUMB[3][23] ), .CO(
        \mult_22/CARRYB[4][22] ), .S(\mult_22/SUMB[4][22] ) );
  FA_X1 \mult_22/S2_4_21  ( .A(\mult_22/ab[4][21] ), .B(
        \mult_22/CARRYB[3][21] ), .CI(\mult_22/SUMB[3][22] ), .CO(
        \mult_22/CARRYB[4][21] ), .S(\mult_22/SUMB[4][21] ) );
  FA_X1 \mult_22/S2_4_20  ( .A(\mult_22/ab[4][20] ), .B(
        \mult_22/CARRYB[3][20] ), .CI(\mult_22/SUMB[3][21] ), .CO(
        \mult_22/CARRYB[4][20] ), .S(\mult_22/SUMB[4][20] ) );
  FA_X1 \mult_22/S2_4_19  ( .A(\mult_22/ab[4][19] ), .B(
        \mult_22/CARRYB[3][19] ), .CI(\mult_22/SUMB[3][20] ), .CO(
        \mult_22/CARRYB[4][19] ), .S(\mult_22/SUMB[4][19] ) );
  FA_X1 \mult_22/S2_4_18  ( .A(\mult_22/ab[4][18] ), .B(
        \mult_22/CARRYB[3][18] ), .CI(\mult_22/SUMB[3][19] ), .CO(
        \mult_22/CARRYB[4][18] ), .S(\mult_22/SUMB[4][18] ) );
  FA_X1 \mult_22/S2_4_17  ( .A(\mult_22/ab[4][17] ), .B(
        \mult_22/CARRYB[3][17] ), .CI(\mult_22/SUMB[3][18] ), .CO(
        \mult_22/CARRYB[4][17] ), .S(\mult_22/SUMB[4][17] ) );
  FA_X1 \mult_22/S2_4_16  ( .A(\mult_22/ab[4][16] ), .B(
        \mult_22/CARRYB[3][16] ), .CI(\mult_22/SUMB[3][17] ), .CO(
        \mult_22/CARRYB[4][16] ), .S(\mult_22/SUMB[4][16] ) );
  FA_X1 \mult_22/S2_4_15  ( .A(\mult_22/ab[4][15] ), .B(
        \mult_22/CARRYB[3][15] ), .CI(\mult_22/SUMB[3][16] ), .CO(
        \mult_22/CARRYB[4][15] ), .S(\mult_22/SUMB[4][15] ) );
  FA_X1 \mult_22/S2_4_14  ( .A(\mult_22/ab[4][14] ), .B(
        \mult_22/CARRYB[3][14] ), .CI(\mult_22/SUMB[3][15] ), .CO(
        \mult_22/CARRYB[4][14] ), .S(\mult_22/SUMB[4][14] ) );
  FA_X1 \mult_22/S2_4_13  ( .A(\mult_22/ab[4][13] ), .B(
        \mult_22/CARRYB[3][13] ), .CI(\mult_22/SUMB[3][14] ), .CO(
        \mult_22/CARRYB[4][13] ), .S(\mult_22/SUMB[4][13] ) );
  FA_X1 \mult_22/S2_4_12  ( .A(\mult_22/ab[4][12] ), .B(
        \mult_22/CARRYB[3][12] ), .CI(\mult_22/SUMB[3][13] ), .CO(
        \mult_22/CARRYB[4][12] ), .S(\mult_22/SUMB[4][12] ) );
  FA_X1 \mult_22/S2_4_11  ( .A(\mult_22/ab[4][11] ), .B(
        \mult_22/CARRYB[3][11] ), .CI(\mult_22/SUMB[3][12] ), .CO(
        \mult_22/CARRYB[4][11] ), .S(\mult_22/SUMB[4][11] ) );
  FA_X1 \mult_22/S2_4_10  ( .A(\mult_22/ab[4][10] ), .B(
        \mult_22/CARRYB[3][10] ), .CI(\mult_22/SUMB[3][11] ), .CO(
        \mult_22/CARRYB[4][10] ), .S(\mult_22/SUMB[4][10] ) );
  FA_X1 \mult_22/S2_4_9  ( .A(\mult_22/ab[4][9] ), .B(\mult_22/CARRYB[3][9] ), 
        .CI(\mult_22/SUMB[3][10] ), .CO(\mult_22/CARRYB[4][9] ), .S(
        \mult_22/SUMB[4][9] ) );
  FA_X1 \mult_22/S2_4_8  ( .A(\mult_22/ab[4][8] ), .B(\mult_22/CARRYB[3][8] ), 
        .CI(\mult_22/SUMB[3][9] ), .CO(\mult_22/CARRYB[4][8] ), .S(
        \mult_22/SUMB[4][8] ) );
  FA_X1 \mult_22/S2_4_7  ( .A(\mult_22/ab[4][7] ), .B(\mult_22/CARRYB[3][7] ), 
        .CI(\mult_22/SUMB[3][8] ), .CO(\mult_22/CARRYB[4][7] ), .S(
        \mult_22/SUMB[4][7] ) );
  FA_X1 \mult_22/S2_4_6  ( .A(\mult_22/ab[4][6] ), .B(\mult_22/CARRYB[3][6] ), 
        .CI(\mult_22/SUMB[3][7] ), .CO(\mult_22/CARRYB[4][6] ), .S(
        \mult_22/SUMB[4][6] ) );
  FA_X1 \mult_22/S2_4_5  ( .A(\mult_22/ab[4][5] ), .B(\mult_22/CARRYB[3][5] ), 
        .CI(\mult_22/SUMB[3][6] ), .CO(\mult_22/CARRYB[4][5] ), .S(
        \mult_22/SUMB[4][5] ) );
  FA_X1 \mult_22/S2_4_4  ( .A(\mult_22/ab[4][4] ), .B(\mult_22/CARRYB[3][4] ), 
        .CI(\mult_22/SUMB[3][5] ), .CO(\mult_22/CARRYB[4][4] ), .S(
        \mult_22/SUMB[4][4] ) );
  FA_X1 \mult_22/S2_4_3  ( .A(\mult_22/ab[4][3] ), .B(\mult_22/CARRYB[3][3] ), 
        .CI(\mult_22/SUMB[3][4] ), .CO(\mult_22/CARRYB[4][3] ), .S(
        \mult_22/SUMB[4][3] ) );
  FA_X1 \mult_22/S2_4_2  ( .A(\mult_22/ab[4][2] ), .B(\mult_22/CARRYB[3][2] ), 
        .CI(\mult_22/SUMB[3][3] ), .CO(\mult_22/CARRYB[4][2] ), .S(
        \mult_22/SUMB[4][2] ) );
  FA_X1 \mult_22/S2_4_1  ( .A(\mult_22/ab[4][1] ), .B(\mult_22/CARRYB[3][1] ), 
        .CI(\mult_22/SUMB[3][2] ), .CO(\mult_22/CARRYB[4][1] ), .S(
        \mult_22/SUMB[4][1] ) );
  FA_X1 \mult_22/S1_4_0  ( .A(\mult_22/ab[4][0] ), .B(\mult_22/CARRYB[3][0] ), 
        .CI(\mult_22/SUMB[3][1] ), .CO(\mult_22/CARRYB[4][0] ), .S(N132) );
  FA_X1 \mult_22/S3_5_62  ( .A(\mult_22/ab[5][62] ), .B(
        \mult_22/CARRYB[4][62] ), .CI(\mult_22/ab[4][63] ), .CO(
        \mult_22/CARRYB[5][62] ), .S(\mult_22/SUMB[5][62] ) );
  FA_X1 \mult_22/S2_5_59  ( .A(\mult_22/CARRYB[4][59] ), .B(
        \mult_22/ab[5][59] ), .CI(\mult_22/SUMB[4][60] ), .CO(
        \mult_22/CARRYB[5][59] ), .S(\mult_22/SUMB[5][59] ) );
  FA_X1 \mult_22/S2_5_58  ( .A(\mult_22/ab[5][58] ), .B(
        \mult_22/CARRYB[4][58] ), .CI(\mult_22/SUMB[4][59] ), .CO(
        \mult_22/CARRYB[5][58] ), .S(\mult_22/SUMB[5][58] ) );
  FA_X1 \mult_22/S2_5_57  ( .A(\mult_22/ab[5][57] ), .B(
        \mult_22/CARRYB[4][57] ), .CI(\mult_22/SUMB[4][58] ), .CO(
        \mult_22/CARRYB[5][57] ), .S(\mult_22/SUMB[5][57] ) );
  FA_X1 \mult_22/S2_5_56  ( .A(\mult_22/CARRYB[4][56] ), .B(
        \mult_22/ab[5][56] ), .CI(\mult_22/SUMB[4][57] ), .CO(
        \mult_22/CARRYB[5][56] ), .S(\mult_22/SUMB[5][56] ) );
  FA_X1 \mult_22/S2_5_55  ( .A(\mult_22/ab[5][55] ), .B(
        \mult_22/CARRYB[4][55] ), .CI(\mult_22/SUMB[4][56] ), .CO(
        \mult_22/CARRYB[5][55] ), .S(\mult_22/SUMB[5][55] ) );
  FA_X1 \mult_22/S2_5_53  ( .A(\mult_22/ab[5][53] ), .B(
        \mult_22/CARRYB[4][53] ), .CI(\mult_22/SUMB[4][54] ), .CO(
        \mult_22/CARRYB[5][53] ), .S(\mult_22/SUMB[5][53] ) );
  FA_X1 \mult_22/S2_5_52  ( .A(\mult_22/CARRYB[4][52] ), .B(
        \mult_22/ab[5][52] ), .CI(\mult_22/SUMB[4][53] ), .CO(
        \mult_22/CARRYB[5][52] ), .S(\mult_22/SUMB[5][52] ) );
  FA_X1 \mult_22/S2_5_51  ( .A(\mult_22/ab[5][51] ), .B(
        \mult_22/CARRYB[4][51] ), .CI(\mult_22/SUMB[4][52] ), .CO(
        \mult_22/CARRYB[5][51] ), .S(\mult_22/SUMB[5][51] ) );
  FA_X1 \mult_22/S2_5_50  ( .A(\mult_22/ab[5][50] ), .B(
        \mult_22/CARRYB[4][50] ), .CI(\mult_22/SUMB[4][51] ), .CO(
        \mult_22/CARRYB[5][50] ), .S(\mult_22/SUMB[5][50] ) );
  FA_X1 \mult_22/S2_5_49  ( .A(\mult_22/ab[5][49] ), .B(
        \mult_22/CARRYB[4][49] ), .CI(\mult_22/SUMB[4][50] ), .CO(
        \mult_22/CARRYB[5][49] ), .S(\mult_22/SUMB[5][49] ) );
  FA_X1 \mult_22/S2_5_48  ( .A(\mult_22/ab[5][48] ), .B(
        \mult_22/CARRYB[4][48] ), .CI(\mult_22/SUMB[4][49] ), .CO(
        \mult_22/CARRYB[5][48] ), .S(\mult_22/SUMB[5][48] ) );
  FA_X1 \mult_22/S2_5_47  ( .A(\mult_22/ab[5][47] ), .B(
        \mult_22/CARRYB[4][47] ), .CI(\mult_22/SUMB[4][48] ), .CO(
        \mult_22/CARRYB[5][47] ), .S(\mult_22/SUMB[5][47] ) );
  FA_X1 \mult_22/S2_5_46  ( .A(\mult_22/ab[5][46] ), .B(
        \mult_22/CARRYB[4][46] ), .CI(\mult_22/SUMB[4][47] ), .CO(
        \mult_22/CARRYB[5][46] ), .S(\mult_22/SUMB[5][46] ) );
  FA_X1 \mult_22/S2_5_45  ( .A(\mult_22/ab[5][45] ), .B(
        \mult_22/CARRYB[4][45] ), .CI(\mult_22/SUMB[4][46] ), .CO(
        \mult_22/CARRYB[5][45] ), .S(\mult_22/SUMB[5][45] ) );
  FA_X1 \mult_22/S2_5_44  ( .A(\mult_22/ab[5][44] ), .B(
        \mult_22/CARRYB[4][44] ), .CI(\mult_22/SUMB[4][45] ), .CO(
        \mult_22/CARRYB[5][44] ), .S(\mult_22/SUMB[5][44] ) );
  FA_X1 \mult_22/S2_5_43  ( .A(\mult_22/ab[5][43] ), .B(
        \mult_22/CARRYB[4][43] ), .CI(\mult_22/SUMB[4][44] ), .CO(
        \mult_22/CARRYB[5][43] ), .S(\mult_22/SUMB[5][43] ) );
  FA_X1 \mult_22/S2_5_42  ( .A(\mult_22/ab[5][42] ), .B(
        \mult_22/CARRYB[4][42] ), .CI(\mult_22/SUMB[4][43] ), .CO(
        \mult_22/CARRYB[5][42] ), .S(\mult_22/SUMB[5][42] ) );
  FA_X1 \mult_22/S2_5_41  ( .A(\mult_22/ab[5][41] ), .B(
        \mult_22/CARRYB[4][41] ), .CI(\mult_22/SUMB[4][42] ), .CO(
        \mult_22/CARRYB[5][41] ), .S(\mult_22/SUMB[5][41] ) );
  FA_X1 \mult_22/S2_5_40  ( .A(\mult_22/ab[5][40] ), .B(
        \mult_22/CARRYB[4][40] ), .CI(\mult_22/SUMB[4][41] ), .CO(
        \mult_22/CARRYB[5][40] ), .S(\mult_22/SUMB[5][40] ) );
  FA_X1 \mult_22/S2_5_39  ( .A(\mult_22/ab[5][39] ), .B(
        \mult_22/CARRYB[4][39] ), .CI(\mult_22/SUMB[4][40] ), .CO(
        \mult_22/CARRYB[5][39] ), .S(\mult_22/SUMB[5][39] ) );
  FA_X1 \mult_22/S2_5_38  ( .A(\mult_22/ab[5][38] ), .B(
        \mult_22/CARRYB[4][38] ), .CI(\mult_22/SUMB[4][39] ), .CO(
        \mult_22/CARRYB[5][38] ), .S(\mult_22/SUMB[5][38] ) );
  FA_X1 \mult_22/S2_5_37  ( .A(\mult_22/ab[5][37] ), .B(
        \mult_22/CARRYB[4][37] ), .CI(\mult_22/SUMB[4][38] ), .CO(
        \mult_22/CARRYB[5][37] ), .S(\mult_22/SUMB[5][37] ) );
  FA_X1 \mult_22/S2_5_36  ( .A(\mult_22/ab[5][36] ), .B(
        \mult_22/CARRYB[4][36] ), .CI(\mult_22/SUMB[4][37] ), .CO(
        \mult_22/CARRYB[5][36] ), .S(\mult_22/SUMB[5][36] ) );
  FA_X1 \mult_22/S2_5_35  ( .A(\mult_22/ab[5][35] ), .B(
        \mult_22/CARRYB[4][35] ), .CI(\mult_22/SUMB[4][36] ), .CO(
        \mult_22/CARRYB[5][35] ), .S(\mult_22/SUMB[5][35] ) );
  FA_X1 \mult_22/S2_5_34  ( .A(\mult_22/ab[5][34] ), .B(
        \mult_22/CARRYB[4][34] ), .CI(\mult_22/SUMB[4][35] ), .CO(
        \mult_22/CARRYB[5][34] ), .S(\mult_22/SUMB[5][34] ) );
  FA_X1 \mult_22/S2_5_33  ( .A(\mult_22/ab[5][33] ), .B(
        \mult_22/CARRYB[4][33] ), .CI(\mult_22/SUMB[4][34] ), .CO(
        \mult_22/CARRYB[5][33] ), .S(\mult_22/SUMB[5][33] ) );
  FA_X1 \mult_22/S2_5_32  ( .A(\mult_22/ab[5][32] ), .B(
        \mult_22/CARRYB[4][32] ), .CI(\mult_22/SUMB[4][33] ), .CO(
        \mult_22/CARRYB[5][32] ), .S(\mult_22/SUMB[5][32] ) );
  FA_X1 \mult_22/S2_5_31  ( .A(\mult_22/ab[5][31] ), .B(
        \mult_22/CARRYB[4][31] ), .CI(\mult_22/SUMB[4][32] ), .CO(
        \mult_22/CARRYB[5][31] ), .S(\mult_22/SUMB[5][31] ) );
  FA_X1 \mult_22/S2_5_30  ( .A(\mult_22/ab[5][30] ), .B(
        \mult_22/CARRYB[4][30] ), .CI(\mult_22/SUMB[4][31] ), .CO(
        \mult_22/CARRYB[5][30] ), .S(\mult_22/SUMB[5][30] ) );
  FA_X1 \mult_22/S2_5_29  ( .A(\mult_22/ab[5][29] ), .B(
        \mult_22/CARRYB[4][29] ), .CI(\mult_22/SUMB[4][30] ), .CO(
        \mult_22/CARRYB[5][29] ), .S(\mult_22/SUMB[5][29] ) );
  FA_X1 \mult_22/S2_5_28  ( .A(\mult_22/ab[5][28] ), .B(
        \mult_22/CARRYB[4][28] ), .CI(\mult_22/SUMB[4][29] ), .CO(
        \mult_22/CARRYB[5][28] ), .S(\mult_22/SUMB[5][28] ) );
  FA_X1 \mult_22/S2_5_27  ( .A(\mult_22/ab[5][27] ), .B(
        \mult_22/CARRYB[4][27] ), .CI(\mult_22/SUMB[4][28] ), .CO(
        \mult_22/CARRYB[5][27] ), .S(\mult_22/SUMB[5][27] ) );
  FA_X1 \mult_22/S2_5_26  ( .A(\mult_22/ab[5][26] ), .B(
        \mult_22/CARRYB[4][26] ), .CI(\mult_22/SUMB[4][27] ), .CO(
        \mult_22/CARRYB[5][26] ), .S(\mult_22/SUMB[5][26] ) );
  FA_X1 \mult_22/S2_5_25  ( .A(\mult_22/ab[5][25] ), .B(
        \mult_22/CARRYB[4][25] ), .CI(\mult_22/SUMB[4][26] ), .CO(
        \mult_22/CARRYB[5][25] ), .S(\mult_22/SUMB[5][25] ) );
  FA_X1 \mult_22/S2_5_24  ( .A(\mult_22/ab[5][24] ), .B(
        \mult_22/CARRYB[4][24] ), .CI(\mult_22/SUMB[4][25] ), .CO(
        \mult_22/CARRYB[5][24] ), .S(\mult_22/SUMB[5][24] ) );
  FA_X1 \mult_22/S2_5_23  ( .A(\mult_22/ab[5][23] ), .B(
        \mult_22/CARRYB[4][23] ), .CI(\mult_22/SUMB[4][24] ), .CO(
        \mult_22/CARRYB[5][23] ), .S(\mult_22/SUMB[5][23] ) );
  FA_X1 \mult_22/S2_5_22  ( .A(\mult_22/ab[5][22] ), .B(
        \mult_22/CARRYB[4][22] ), .CI(\mult_22/SUMB[4][23] ), .CO(
        \mult_22/CARRYB[5][22] ), .S(\mult_22/SUMB[5][22] ) );
  FA_X1 \mult_22/S2_5_21  ( .A(\mult_22/ab[5][21] ), .B(
        \mult_22/CARRYB[4][21] ), .CI(\mult_22/SUMB[4][22] ), .CO(
        \mult_22/CARRYB[5][21] ), .S(\mult_22/SUMB[5][21] ) );
  FA_X1 \mult_22/S2_5_20  ( .A(\mult_22/ab[5][20] ), .B(
        \mult_22/CARRYB[4][20] ), .CI(\mult_22/SUMB[4][21] ), .CO(
        \mult_22/CARRYB[5][20] ), .S(\mult_22/SUMB[5][20] ) );
  FA_X1 \mult_22/S2_5_19  ( .A(\mult_22/ab[5][19] ), .B(
        \mult_22/CARRYB[4][19] ), .CI(\mult_22/SUMB[4][20] ), .CO(
        \mult_22/CARRYB[5][19] ), .S(\mult_22/SUMB[5][19] ) );
  FA_X1 \mult_22/S2_5_18  ( .A(\mult_22/ab[5][18] ), .B(
        \mult_22/CARRYB[4][18] ), .CI(\mult_22/SUMB[4][19] ), .CO(
        \mult_22/CARRYB[5][18] ), .S(\mult_22/SUMB[5][18] ) );
  FA_X1 \mult_22/S2_5_17  ( .A(\mult_22/ab[5][17] ), .B(
        \mult_22/CARRYB[4][17] ), .CI(\mult_22/SUMB[4][18] ), .CO(
        \mult_22/CARRYB[5][17] ), .S(\mult_22/SUMB[5][17] ) );
  FA_X1 \mult_22/S2_5_16  ( .A(\mult_22/ab[5][16] ), .B(
        \mult_22/CARRYB[4][16] ), .CI(\mult_22/SUMB[4][17] ), .CO(
        \mult_22/CARRYB[5][16] ), .S(\mult_22/SUMB[5][16] ) );
  FA_X1 \mult_22/S2_5_15  ( .A(\mult_22/ab[5][15] ), .B(
        \mult_22/CARRYB[4][15] ), .CI(\mult_22/SUMB[4][16] ), .CO(
        \mult_22/CARRYB[5][15] ), .S(\mult_22/SUMB[5][15] ) );
  FA_X1 \mult_22/S2_5_14  ( .A(\mult_22/ab[5][14] ), .B(
        \mult_22/CARRYB[4][14] ), .CI(\mult_22/SUMB[4][15] ), .CO(
        \mult_22/CARRYB[5][14] ), .S(\mult_22/SUMB[5][14] ) );
  FA_X1 \mult_22/S2_5_13  ( .A(\mult_22/ab[5][13] ), .B(
        \mult_22/CARRYB[4][13] ), .CI(\mult_22/SUMB[4][14] ), .CO(
        \mult_22/CARRYB[5][13] ), .S(\mult_22/SUMB[5][13] ) );
  FA_X1 \mult_22/S2_5_12  ( .A(\mult_22/ab[5][12] ), .B(
        \mult_22/CARRYB[4][12] ), .CI(\mult_22/SUMB[4][13] ), .CO(
        \mult_22/CARRYB[5][12] ), .S(\mult_22/SUMB[5][12] ) );
  FA_X1 \mult_22/S2_5_11  ( .A(\mult_22/ab[5][11] ), .B(
        \mult_22/CARRYB[4][11] ), .CI(\mult_22/SUMB[4][12] ), .CO(
        \mult_22/CARRYB[5][11] ), .S(\mult_22/SUMB[5][11] ) );
  FA_X1 \mult_22/S2_5_10  ( .A(\mult_22/ab[5][10] ), .B(
        \mult_22/CARRYB[4][10] ), .CI(\mult_22/SUMB[4][11] ), .CO(
        \mult_22/CARRYB[5][10] ), .S(\mult_22/SUMB[5][10] ) );
  FA_X1 \mult_22/S2_5_9  ( .A(\mult_22/ab[5][9] ), .B(\mult_22/CARRYB[4][9] ), 
        .CI(\mult_22/SUMB[4][10] ), .CO(\mult_22/CARRYB[5][9] ), .S(
        \mult_22/SUMB[5][9] ) );
  FA_X1 \mult_22/S2_5_8  ( .A(\mult_22/ab[5][8] ), .B(\mult_22/CARRYB[4][8] ), 
        .CI(\mult_22/SUMB[4][9] ), .CO(\mult_22/CARRYB[5][8] ), .S(
        \mult_22/SUMB[5][8] ) );
  FA_X1 \mult_22/S2_5_7  ( .A(\mult_22/ab[5][7] ), .B(\mult_22/CARRYB[4][7] ), 
        .CI(\mult_22/SUMB[4][8] ), .CO(\mult_22/CARRYB[5][7] ), .S(
        \mult_22/SUMB[5][7] ) );
  FA_X1 \mult_22/S2_5_6  ( .A(\mult_22/ab[5][6] ), .B(\mult_22/CARRYB[4][6] ), 
        .CI(\mult_22/SUMB[4][7] ), .CO(\mult_22/CARRYB[5][6] ), .S(
        \mult_22/SUMB[5][6] ) );
  FA_X1 \mult_22/S2_5_5  ( .A(\mult_22/ab[5][5] ), .B(\mult_22/CARRYB[4][5] ), 
        .CI(\mult_22/SUMB[4][6] ), .CO(\mult_22/CARRYB[5][5] ), .S(
        \mult_22/SUMB[5][5] ) );
  FA_X1 \mult_22/S2_5_4  ( .A(\mult_22/ab[5][4] ), .B(\mult_22/CARRYB[4][4] ), 
        .CI(\mult_22/SUMB[4][5] ), .CO(\mult_22/CARRYB[5][4] ), .S(
        \mult_22/SUMB[5][4] ) );
  FA_X1 \mult_22/S2_5_3  ( .A(\mult_22/ab[5][3] ), .B(\mult_22/CARRYB[4][3] ), 
        .CI(\mult_22/SUMB[4][4] ), .CO(\mult_22/CARRYB[5][3] ), .S(
        \mult_22/SUMB[5][3] ) );
  FA_X1 \mult_22/S2_5_2  ( .A(\mult_22/ab[5][2] ), .B(\mult_22/CARRYB[4][2] ), 
        .CI(\mult_22/SUMB[4][3] ), .CO(\mult_22/CARRYB[5][2] ), .S(
        \mult_22/SUMB[5][2] ) );
  FA_X1 \mult_22/S2_5_1  ( .A(\mult_22/ab[5][1] ), .B(\mult_22/CARRYB[4][1] ), 
        .CI(\mult_22/SUMB[4][2] ), .CO(\mult_22/CARRYB[5][1] ), .S(
        \mult_22/SUMB[5][1] ) );
  FA_X1 \mult_22/S1_5_0  ( .A(\mult_22/ab[5][0] ), .B(\mult_22/CARRYB[4][0] ), 
        .CI(\mult_22/SUMB[4][1] ), .CO(\mult_22/CARRYB[5][0] ), .S(N133) );
  FA_X1 \mult_22/S3_6_62  ( .A(\mult_22/ab[6][62] ), .B(
        \mult_22/CARRYB[5][62] ), .CI(\mult_22/ab[5][63] ), .CO(
        \mult_22/CARRYB[6][62] ), .S(\mult_22/SUMB[6][62] ) );
  FA_X1 \mult_22/S2_6_61  ( .A(\mult_22/ab[6][61] ), .B(
        \mult_22/CARRYB[5][61] ), .CI(\mult_22/SUMB[5][62] ), .CO(
        \mult_22/CARRYB[6][61] ), .S(\mult_22/SUMB[6][61] ) );
  FA_X1 \mult_22/S2_6_60  ( .A(\mult_22/ab[6][60] ), .B(
        \mult_22/CARRYB[5][60] ), .CI(\mult_22/SUMB[5][61] ), .CO(
        \mult_22/CARRYB[6][60] ), .S(\mult_22/SUMB[6][60] ) );
  FA_X1 \mult_22/S2_6_59  ( .A(\mult_22/CARRYB[5][59] ), .B(
        \mult_22/ab[6][59] ), .CI(\mult_22/SUMB[5][60] ), .CO(
        \mult_22/CARRYB[6][59] ), .S(\mult_22/SUMB[6][59] ) );
  FA_X1 \mult_22/S2_6_58  ( .A(\mult_22/CARRYB[5][58] ), .B(
        \mult_22/ab[6][58] ), .CI(\mult_22/SUMB[5][59] ), .CO(
        \mult_22/CARRYB[6][58] ), .S(\mult_22/SUMB[6][58] ) );
  FA_X1 \mult_22/S2_6_57  ( .A(\mult_22/ab[6][57] ), .B(
        \mult_22/CARRYB[5][57] ), .CI(\mult_22/SUMB[5][58] ), .CO(
        \mult_22/CARRYB[6][57] ), .S(\mult_22/SUMB[6][57] ) );
  FA_X1 \mult_22/S2_6_56  ( .A(\mult_22/ab[6][56] ), .B(
        \mult_22/CARRYB[5][56] ), .CI(\mult_22/SUMB[5][57] ), .CO(
        \mult_22/CARRYB[6][56] ), .S(\mult_22/SUMB[6][56] ) );
  FA_X1 \mult_22/S2_6_55  ( .A(\mult_22/CARRYB[5][55] ), .B(
        \mult_22/ab[6][55] ), .CI(\mult_22/SUMB[5][56] ), .CO(
        \mult_22/CARRYB[6][55] ), .S(\mult_22/SUMB[6][55] ) );
  FA_X1 \mult_22/S2_6_54  ( .A(\mult_22/ab[6][54] ), .B(
        \mult_22/CARRYB[5][54] ), .CI(\mult_22/SUMB[5][55] ), .CO(
        \mult_22/CARRYB[6][54] ), .S(\mult_22/SUMB[6][54] ) );
  FA_X1 \mult_22/S2_6_53  ( .A(\mult_22/ab[6][53] ), .B(
        \mult_22/CARRYB[5][53] ), .CI(\mult_22/SUMB[5][54] ), .CO(
        \mult_22/CARRYB[6][53] ), .S(\mult_22/SUMB[6][53] ) );
  FA_X1 \mult_22/S2_6_52  ( .A(\mult_22/ab[6][52] ), .B(
        \mult_22/CARRYB[5][52] ), .CI(\mult_22/SUMB[5][53] ), .CO(
        \mult_22/CARRYB[6][52] ), .S(\mult_22/SUMB[6][52] ) );
  FA_X1 \mult_22/S2_6_51  ( .A(\mult_22/ab[6][51] ), .B(
        \mult_22/CARRYB[5][51] ), .CI(\mult_22/SUMB[5][52] ), .CO(
        \mult_22/CARRYB[6][51] ), .S(\mult_22/SUMB[6][51] ) );
  FA_X1 \mult_22/S2_6_50  ( .A(\mult_22/ab[6][50] ), .B(
        \mult_22/CARRYB[5][50] ), .CI(\mult_22/SUMB[5][51] ), .CO(
        \mult_22/CARRYB[6][50] ), .S(\mult_22/SUMB[6][50] ) );
  FA_X1 \mult_22/S2_6_49  ( .A(\mult_22/ab[6][49] ), .B(
        \mult_22/CARRYB[5][49] ), .CI(\mult_22/SUMB[5][50] ), .CO(
        \mult_22/CARRYB[6][49] ), .S(\mult_22/SUMB[6][49] ) );
  FA_X1 \mult_22/S2_6_48  ( .A(\mult_22/ab[6][48] ), .B(
        \mult_22/CARRYB[5][48] ), .CI(\mult_22/SUMB[5][49] ), .CO(
        \mult_22/CARRYB[6][48] ), .S(\mult_22/SUMB[6][48] ) );
  FA_X1 \mult_22/S2_6_47  ( .A(\mult_22/ab[6][47] ), .B(
        \mult_22/CARRYB[5][47] ), .CI(\mult_22/SUMB[5][48] ), .CO(
        \mult_22/CARRYB[6][47] ), .S(\mult_22/SUMB[6][47] ) );
  FA_X1 \mult_22/S2_6_46  ( .A(\mult_22/ab[6][46] ), .B(
        \mult_22/CARRYB[5][46] ), .CI(\mult_22/SUMB[5][47] ), .CO(
        \mult_22/CARRYB[6][46] ), .S(\mult_22/SUMB[6][46] ) );
  FA_X1 \mult_22/S2_6_45  ( .A(\mult_22/ab[6][45] ), .B(
        \mult_22/CARRYB[5][45] ), .CI(\mult_22/SUMB[5][46] ), .CO(
        \mult_22/CARRYB[6][45] ), .S(\mult_22/SUMB[6][45] ) );
  FA_X1 \mult_22/S2_6_44  ( .A(\mult_22/ab[6][44] ), .B(
        \mult_22/CARRYB[5][44] ), .CI(\mult_22/SUMB[5][45] ), .CO(
        \mult_22/CARRYB[6][44] ), .S(\mult_22/SUMB[6][44] ) );
  FA_X1 \mult_22/S2_6_43  ( .A(\mult_22/ab[6][43] ), .B(
        \mult_22/CARRYB[5][43] ), .CI(\mult_22/SUMB[5][44] ), .CO(
        \mult_22/CARRYB[6][43] ), .S(\mult_22/SUMB[6][43] ) );
  FA_X1 \mult_22/S2_6_42  ( .A(\mult_22/ab[6][42] ), .B(
        \mult_22/CARRYB[5][42] ), .CI(\mult_22/SUMB[5][43] ), .CO(
        \mult_22/CARRYB[6][42] ), .S(\mult_22/SUMB[6][42] ) );
  FA_X1 \mult_22/S2_6_41  ( .A(\mult_22/ab[6][41] ), .B(
        \mult_22/CARRYB[5][41] ), .CI(\mult_22/SUMB[5][42] ), .CO(
        \mult_22/CARRYB[6][41] ), .S(\mult_22/SUMB[6][41] ) );
  FA_X1 \mult_22/S2_6_40  ( .A(\mult_22/ab[6][40] ), .B(
        \mult_22/CARRYB[5][40] ), .CI(\mult_22/SUMB[5][41] ), .CO(
        \mult_22/CARRYB[6][40] ), .S(\mult_22/SUMB[6][40] ) );
  FA_X1 \mult_22/S2_6_39  ( .A(\mult_22/ab[6][39] ), .B(
        \mult_22/CARRYB[5][39] ), .CI(\mult_22/SUMB[5][40] ), .CO(
        \mult_22/CARRYB[6][39] ), .S(\mult_22/SUMB[6][39] ) );
  FA_X1 \mult_22/S2_6_38  ( .A(\mult_22/ab[6][38] ), .B(
        \mult_22/CARRYB[5][38] ), .CI(\mult_22/SUMB[5][39] ), .CO(
        \mult_22/CARRYB[6][38] ), .S(\mult_22/SUMB[6][38] ) );
  FA_X1 \mult_22/S2_6_37  ( .A(\mult_22/ab[6][37] ), .B(
        \mult_22/CARRYB[5][37] ), .CI(\mult_22/SUMB[5][38] ), .CO(
        \mult_22/CARRYB[6][37] ), .S(\mult_22/SUMB[6][37] ) );
  FA_X1 \mult_22/S2_6_36  ( .A(\mult_22/ab[6][36] ), .B(
        \mult_22/CARRYB[5][36] ), .CI(\mult_22/SUMB[5][37] ), .CO(
        \mult_22/CARRYB[6][36] ), .S(\mult_22/SUMB[6][36] ) );
  FA_X1 \mult_22/S2_6_35  ( .A(\mult_22/ab[6][35] ), .B(
        \mult_22/CARRYB[5][35] ), .CI(\mult_22/SUMB[5][36] ), .CO(
        \mult_22/CARRYB[6][35] ), .S(\mult_22/SUMB[6][35] ) );
  FA_X1 \mult_22/S2_6_34  ( .A(\mult_22/ab[6][34] ), .B(
        \mult_22/CARRYB[5][34] ), .CI(\mult_22/SUMB[5][35] ), .CO(
        \mult_22/CARRYB[6][34] ), .S(\mult_22/SUMB[6][34] ) );
  FA_X1 \mult_22/S2_6_33  ( .A(\mult_22/ab[6][33] ), .B(
        \mult_22/CARRYB[5][33] ), .CI(\mult_22/SUMB[5][34] ), .CO(
        \mult_22/CARRYB[6][33] ), .S(\mult_22/SUMB[6][33] ) );
  FA_X1 \mult_22/S2_6_32  ( .A(\mult_22/ab[6][32] ), .B(
        \mult_22/CARRYB[5][32] ), .CI(\mult_22/SUMB[5][33] ), .CO(
        \mult_22/CARRYB[6][32] ), .S(\mult_22/SUMB[6][32] ) );
  FA_X1 \mult_22/S2_6_31  ( .A(\mult_22/ab[6][31] ), .B(
        \mult_22/CARRYB[5][31] ), .CI(\mult_22/SUMB[5][32] ), .CO(
        \mult_22/CARRYB[6][31] ), .S(\mult_22/SUMB[6][31] ) );
  FA_X1 \mult_22/S2_6_30  ( .A(\mult_22/ab[6][30] ), .B(
        \mult_22/CARRYB[5][30] ), .CI(\mult_22/SUMB[5][31] ), .CO(
        \mult_22/CARRYB[6][30] ), .S(\mult_22/SUMB[6][30] ) );
  FA_X1 \mult_22/S2_6_29  ( .A(\mult_22/ab[6][29] ), .B(
        \mult_22/CARRYB[5][29] ), .CI(\mult_22/SUMB[5][30] ), .CO(
        \mult_22/CARRYB[6][29] ), .S(\mult_22/SUMB[6][29] ) );
  FA_X1 \mult_22/S2_6_28  ( .A(\mult_22/ab[6][28] ), .B(
        \mult_22/CARRYB[5][28] ), .CI(\mult_22/SUMB[5][29] ), .CO(
        \mult_22/CARRYB[6][28] ), .S(\mult_22/SUMB[6][28] ) );
  FA_X1 \mult_22/S2_6_27  ( .A(\mult_22/ab[6][27] ), .B(
        \mult_22/CARRYB[5][27] ), .CI(\mult_22/SUMB[5][28] ), .CO(
        \mult_22/CARRYB[6][27] ), .S(\mult_22/SUMB[6][27] ) );
  FA_X1 \mult_22/S2_6_26  ( .A(\mult_22/ab[6][26] ), .B(
        \mult_22/CARRYB[5][26] ), .CI(\mult_22/SUMB[5][27] ), .CO(
        \mult_22/CARRYB[6][26] ), .S(\mult_22/SUMB[6][26] ) );
  FA_X1 \mult_22/S2_6_25  ( .A(\mult_22/ab[6][25] ), .B(
        \mult_22/CARRYB[5][25] ), .CI(\mult_22/SUMB[5][26] ), .CO(
        \mult_22/CARRYB[6][25] ), .S(\mult_22/SUMB[6][25] ) );
  FA_X1 \mult_22/S2_6_24  ( .A(\mult_22/ab[6][24] ), .B(
        \mult_22/CARRYB[5][24] ), .CI(\mult_22/SUMB[5][25] ), .CO(
        \mult_22/CARRYB[6][24] ), .S(\mult_22/SUMB[6][24] ) );
  FA_X1 \mult_22/S2_6_23  ( .A(\mult_22/ab[6][23] ), .B(
        \mult_22/CARRYB[5][23] ), .CI(\mult_22/SUMB[5][24] ), .CO(
        \mult_22/CARRYB[6][23] ), .S(\mult_22/SUMB[6][23] ) );
  FA_X1 \mult_22/S2_6_22  ( .A(\mult_22/ab[6][22] ), .B(
        \mult_22/CARRYB[5][22] ), .CI(\mult_22/SUMB[5][23] ), .CO(
        \mult_22/CARRYB[6][22] ), .S(\mult_22/SUMB[6][22] ) );
  FA_X1 \mult_22/S2_6_21  ( .A(\mult_22/ab[6][21] ), .B(
        \mult_22/CARRYB[5][21] ), .CI(\mult_22/SUMB[5][22] ), .CO(
        \mult_22/CARRYB[6][21] ), .S(\mult_22/SUMB[6][21] ) );
  FA_X1 \mult_22/S2_6_20  ( .A(\mult_22/ab[6][20] ), .B(
        \mult_22/CARRYB[5][20] ), .CI(\mult_22/SUMB[5][21] ), .CO(
        \mult_22/CARRYB[6][20] ), .S(\mult_22/SUMB[6][20] ) );
  FA_X1 \mult_22/S2_6_19  ( .A(\mult_22/ab[6][19] ), .B(
        \mult_22/CARRYB[5][19] ), .CI(\mult_22/SUMB[5][20] ), .CO(
        \mult_22/CARRYB[6][19] ), .S(\mult_22/SUMB[6][19] ) );
  FA_X1 \mult_22/S2_6_18  ( .A(\mult_22/ab[6][18] ), .B(
        \mult_22/CARRYB[5][18] ), .CI(\mult_22/SUMB[5][19] ), .CO(
        \mult_22/CARRYB[6][18] ), .S(\mult_22/SUMB[6][18] ) );
  FA_X1 \mult_22/S2_6_17  ( .A(\mult_22/ab[6][17] ), .B(
        \mult_22/CARRYB[5][17] ), .CI(\mult_22/SUMB[5][18] ), .CO(
        \mult_22/CARRYB[6][17] ), .S(\mult_22/SUMB[6][17] ) );
  FA_X1 \mult_22/S2_6_16  ( .A(\mult_22/ab[6][16] ), .B(
        \mult_22/CARRYB[5][16] ), .CI(\mult_22/SUMB[5][17] ), .CO(
        \mult_22/CARRYB[6][16] ), .S(\mult_22/SUMB[6][16] ) );
  FA_X1 \mult_22/S2_6_15  ( .A(\mult_22/ab[6][15] ), .B(
        \mult_22/CARRYB[5][15] ), .CI(\mult_22/SUMB[5][16] ), .CO(
        \mult_22/CARRYB[6][15] ), .S(\mult_22/SUMB[6][15] ) );
  FA_X1 \mult_22/S2_6_14  ( .A(\mult_22/ab[6][14] ), .B(
        \mult_22/CARRYB[5][14] ), .CI(\mult_22/SUMB[5][15] ), .CO(
        \mult_22/CARRYB[6][14] ), .S(\mult_22/SUMB[6][14] ) );
  FA_X1 \mult_22/S2_6_13  ( .A(\mult_22/ab[6][13] ), .B(
        \mult_22/CARRYB[5][13] ), .CI(\mult_22/SUMB[5][14] ), .CO(
        \mult_22/CARRYB[6][13] ), .S(\mult_22/SUMB[6][13] ) );
  FA_X1 \mult_22/S2_6_12  ( .A(\mult_22/ab[6][12] ), .B(
        \mult_22/CARRYB[5][12] ), .CI(\mult_22/SUMB[5][13] ), .CO(
        \mult_22/CARRYB[6][12] ), .S(\mult_22/SUMB[6][12] ) );
  FA_X1 \mult_22/S2_6_11  ( .A(\mult_22/ab[6][11] ), .B(
        \mult_22/CARRYB[5][11] ), .CI(\mult_22/SUMB[5][12] ), .CO(
        \mult_22/CARRYB[6][11] ), .S(\mult_22/SUMB[6][11] ) );
  FA_X1 \mult_22/S2_6_10  ( .A(\mult_22/ab[6][10] ), .B(
        \mult_22/CARRYB[5][10] ), .CI(\mult_22/SUMB[5][11] ), .CO(
        \mult_22/CARRYB[6][10] ), .S(\mult_22/SUMB[6][10] ) );
  FA_X1 \mult_22/S2_6_9  ( .A(\mult_22/ab[6][9] ), .B(\mult_22/CARRYB[5][9] ), 
        .CI(\mult_22/SUMB[5][10] ), .CO(\mult_22/CARRYB[6][9] ), .S(
        \mult_22/SUMB[6][9] ) );
  FA_X1 \mult_22/S2_6_8  ( .A(\mult_22/ab[6][8] ), .B(\mult_22/CARRYB[5][8] ), 
        .CI(\mult_22/SUMB[5][9] ), .CO(\mult_22/CARRYB[6][8] ), .S(
        \mult_22/SUMB[6][8] ) );
  FA_X1 \mult_22/S2_6_7  ( .A(\mult_22/ab[6][7] ), .B(\mult_22/CARRYB[5][7] ), 
        .CI(\mult_22/SUMB[5][8] ), .CO(\mult_22/CARRYB[6][7] ), .S(
        \mult_22/SUMB[6][7] ) );
  FA_X1 \mult_22/S2_6_6  ( .A(\mult_22/ab[6][6] ), .B(\mult_22/CARRYB[5][6] ), 
        .CI(\mult_22/SUMB[5][7] ), .CO(\mult_22/CARRYB[6][6] ), .S(
        \mult_22/SUMB[6][6] ) );
  FA_X1 \mult_22/S2_6_5  ( .A(\mult_22/ab[6][5] ), .B(\mult_22/CARRYB[5][5] ), 
        .CI(\mult_22/SUMB[5][6] ), .CO(\mult_22/CARRYB[6][5] ), .S(
        \mult_22/SUMB[6][5] ) );
  FA_X1 \mult_22/S2_6_4  ( .A(\mult_22/ab[6][4] ), .B(\mult_22/CARRYB[5][4] ), 
        .CI(\mult_22/SUMB[5][5] ), .CO(\mult_22/CARRYB[6][4] ), .S(
        \mult_22/SUMB[6][4] ) );
  FA_X1 \mult_22/S2_6_3  ( .A(\mult_22/ab[6][3] ), .B(\mult_22/CARRYB[5][3] ), 
        .CI(\mult_22/SUMB[5][4] ), .CO(\mult_22/CARRYB[6][3] ), .S(
        \mult_22/SUMB[6][3] ) );
  FA_X1 \mult_22/S2_6_2  ( .A(\mult_22/ab[6][2] ), .B(\mult_22/CARRYB[5][2] ), 
        .CI(\mult_22/SUMB[5][3] ), .CO(\mult_22/CARRYB[6][2] ), .S(
        \mult_22/SUMB[6][2] ) );
  FA_X1 \mult_22/S2_6_1  ( .A(\mult_22/ab[6][1] ), .B(\mult_22/CARRYB[5][1] ), 
        .CI(\mult_22/SUMB[5][2] ), .CO(\mult_22/CARRYB[6][1] ), .S(
        \mult_22/SUMB[6][1] ) );
  FA_X1 \mult_22/S1_6_0  ( .A(\mult_22/ab[6][0] ), .B(\mult_22/CARRYB[5][0] ), 
        .CI(\mult_22/SUMB[5][1] ), .CO(\mult_22/CARRYB[6][0] ), .S(N134) );
  FA_X1 \mult_22/S3_7_62  ( .A(\mult_22/ab[7][62] ), .B(
        \mult_22/CARRYB[6][62] ), .CI(\mult_22/ab[6][63] ), .CO(
        \mult_22/CARRYB[7][62] ), .S(\mult_22/SUMB[7][62] ) );
  FA_X1 \mult_22/S2_7_61  ( .A(\mult_22/ab[7][61] ), .B(
        \mult_22/CARRYB[6][61] ), .CI(\mult_22/SUMB[6][62] ), .CO(
        \mult_22/CARRYB[7][61] ), .S(\mult_22/SUMB[7][61] ) );
  FA_X1 \mult_22/S2_7_60  ( .A(\mult_22/ab[7][60] ), .B(
        \mult_22/CARRYB[6][60] ), .CI(\mult_22/SUMB[6][61] ), .CO(
        \mult_22/CARRYB[7][60] ), .S(\mult_22/SUMB[7][60] ) );
  FA_X1 \mult_22/S2_7_59  ( .A(\mult_22/ab[7][59] ), .B(
        \mult_22/CARRYB[6][59] ), .CI(\mult_22/SUMB[6][60] ), .CO(
        \mult_22/CARRYB[7][59] ), .S(\mult_22/SUMB[7][59] ) );
  FA_X1 \mult_22/S2_7_58  ( .A(\mult_22/CARRYB[6][58] ), .B(
        \mult_22/ab[7][58] ), .CI(\mult_22/SUMB[6][59] ), .CO(
        \mult_22/CARRYB[7][58] ), .S(\mult_22/SUMB[7][58] ) );
  FA_X1 \mult_22/S2_7_57  ( .A(\mult_22/CARRYB[6][57] ), .B(
        \mult_22/ab[7][57] ), .CI(\mult_22/SUMB[6][58] ), .CO(
        \mult_22/CARRYB[7][57] ), .S(\mult_22/SUMB[7][57] ) );
  FA_X1 \mult_22/S2_7_56  ( .A(\mult_22/ab[7][56] ), .B(
        \mult_22/CARRYB[6][56] ), .CI(\mult_22/SUMB[6][57] ), .CO(
        \mult_22/CARRYB[7][56] ), .S(\mult_22/SUMB[7][56] ) );
  FA_X1 \mult_22/S2_7_55  ( .A(\mult_22/ab[7][55] ), .B(
        \mult_22/CARRYB[6][55] ), .CI(\mult_22/SUMB[6][56] ), .CO(
        \mult_22/CARRYB[7][55] ), .S(\mult_22/SUMB[7][55] ) );
  FA_X1 \mult_22/S2_7_54  ( .A(\mult_22/ab[7][54] ), .B(
        \mult_22/CARRYB[6][54] ), .CI(\mult_22/SUMB[6][55] ), .CO(
        \mult_22/CARRYB[7][54] ), .S(\mult_22/SUMB[7][54] ) );
  FA_X1 \mult_22/S2_7_53  ( .A(\mult_22/ab[7][53] ), .B(
        \mult_22/CARRYB[6][53] ), .CI(\mult_22/SUMB[6][54] ), .CO(
        \mult_22/CARRYB[7][53] ), .S(\mult_22/SUMB[7][53] ) );
  FA_X1 \mult_22/S2_7_52  ( .A(\mult_22/ab[7][52] ), .B(
        \mult_22/CARRYB[6][52] ), .CI(\mult_22/SUMB[6][53] ), .CO(
        \mult_22/CARRYB[7][52] ), .S(\mult_22/SUMB[7][52] ) );
  FA_X1 \mult_22/S2_7_51  ( .A(\mult_22/ab[7][51] ), .B(
        \mult_22/CARRYB[6][51] ), .CI(\mult_22/SUMB[6][52] ), .CO(
        \mult_22/CARRYB[7][51] ), .S(\mult_22/SUMB[7][51] ) );
  FA_X1 \mult_22/S2_7_50  ( .A(\mult_22/ab[7][50] ), .B(
        \mult_22/CARRYB[6][50] ), .CI(\mult_22/SUMB[6][51] ), .CO(
        \mult_22/CARRYB[7][50] ), .S(\mult_22/SUMB[7][50] ) );
  FA_X1 \mult_22/S2_7_49  ( .A(\mult_22/ab[7][49] ), .B(
        \mult_22/CARRYB[6][49] ), .CI(\mult_22/SUMB[6][50] ), .CO(
        \mult_22/CARRYB[7][49] ), .S(\mult_22/SUMB[7][49] ) );
  FA_X1 \mult_22/S2_7_48  ( .A(\mult_22/ab[7][48] ), .B(
        \mult_22/CARRYB[6][48] ), .CI(\mult_22/SUMB[6][49] ), .CO(
        \mult_22/CARRYB[7][48] ), .S(\mult_22/SUMB[7][48] ) );
  FA_X1 \mult_22/S2_7_47  ( .A(\mult_22/ab[7][47] ), .B(
        \mult_22/CARRYB[6][47] ), .CI(\mult_22/SUMB[6][48] ), .CO(
        \mult_22/CARRYB[7][47] ), .S(\mult_22/SUMB[7][47] ) );
  FA_X1 \mult_22/S2_7_46  ( .A(\mult_22/ab[7][46] ), .B(
        \mult_22/CARRYB[6][46] ), .CI(\mult_22/SUMB[6][47] ), .CO(
        \mult_22/CARRYB[7][46] ), .S(\mult_22/SUMB[7][46] ) );
  FA_X1 \mult_22/S2_7_45  ( .A(\mult_22/ab[7][45] ), .B(
        \mult_22/CARRYB[6][45] ), .CI(\mult_22/SUMB[6][46] ), .CO(
        \mult_22/CARRYB[7][45] ), .S(\mult_22/SUMB[7][45] ) );
  FA_X1 \mult_22/S2_7_44  ( .A(\mult_22/ab[7][44] ), .B(
        \mult_22/CARRYB[6][44] ), .CI(\mult_22/SUMB[6][45] ), .CO(
        \mult_22/CARRYB[7][44] ), .S(\mult_22/SUMB[7][44] ) );
  FA_X1 \mult_22/S2_7_43  ( .A(\mult_22/ab[7][43] ), .B(
        \mult_22/CARRYB[6][43] ), .CI(\mult_22/SUMB[6][44] ), .CO(
        \mult_22/CARRYB[7][43] ), .S(\mult_22/SUMB[7][43] ) );
  FA_X1 \mult_22/S2_7_42  ( .A(\mult_22/ab[7][42] ), .B(
        \mult_22/CARRYB[6][42] ), .CI(\mult_22/SUMB[6][43] ), .CO(
        \mult_22/CARRYB[7][42] ), .S(\mult_22/SUMB[7][42] ) );
  FA_X1 \mult_22/S2_7_41  ( .A(\mult_22/ab[7][41] ), .B(
        \mult_22/CARRYB[6][41] ), .CI(\mult_22/SUMB[6][42] ), .CO(
        \mult_22/CARRYB[7][41] ), .S(\mult_22/SUMB[7][41] ) );
  FA_X1 \mult_22/S2_7_40  ( .A(\mult_22/ab[7][40] ), .B(
        \mult_22/CARRYB[6][40] ), .CI(\mult_22/SUMB[6][41] ), .CO(
        \mult_22/CARRYB[7][40] ), .S(\mult_22/SUMB[7][40] ) );
  FA_X1 \mult_22/S2_7_39  ( .A(\mult_22/ab[7][39] ), .B(
        \mult_22/CARRYB[6][39] ), .CI(\mult_22/SUMB[6][40] ), .CO(
        \mult_22/CARRYB[7][39] ), .S(\mult_22/SUMB[7][39] ) );
  FA_X1 \mult_22/S2_7_38  ( .A(\mult_22/ab[7][38] ), .B(
        \mult_22/CARRYB[6][38] ), .CI(\mult_22/SUMB[6][39] ), .CO(
        \mult_22/CARRYB[7][38] ), .S(\mult_22/SUMB[7][38] ) );
  FA_X1 \mult_22/S2_7_37  ( .A(\mult_22/ab[7][37] ), .B(
        \mult_22/CARRYB[6][37] ), .CI(\mult_22/SUMB[6][38] ), .CO(
        \mult_22/CARRYB[7][37] ), .S(\mult_22/SUMB[7][37] ) );
  FA_X1 \mult_22/S2_7_36  ( .A(\mult_22/ab[7][36] ), .B(
        \mult_22/CARRYB[6][36] ), .CI(\mult_22/SUMB[6][37] ), .CO(
        \mult_22/CARRYB[7][36] ), .S(\mult_22/SUMB[7][36] ) );
  FA_X1 \mult_22/S2_7_35  ( .A(\mult_22/ab[7][35] ), .B(
        \mult_22/CARRYB[6][35] ), .CI(\mult_22/SUMB[6][36] ), .CO(
        \mult_22/CARRYB[7][35] ), .S(\mult_22/SUMB[7][35] ) );
  FA_X1 \mult_22/S2_7_34  ( .A(\mult_22/ab[7][34] ), .B(
        \mult_22/CARRYB[6][34] ), .CI(\mult_22/SUMB[6][35] ), .CO(
        \mult_22/CARRYB[7][34] ), .S(\mult_22/SUMB[7][34] ) );
  FA_X1 \mult_22/S2_7_33  ( .A(\mult_22/ab[7][33] ), .B(
        \mult_22/CARRYB[6][33] ), .CI(\mult_22/SUMB[6][34] ), .CO(
        \mult_22/CARRYB[7][33] ), .S(\mult_22/SUMB[7][33] ) );
  FA_X1 \mult_22/S2_7_32  ( .A(\mult_22/ab[7][32] ), .B(
        \mult_22/CARRYB[6][32] ), .CI(\mult_22/SUMB[6][33] ), .CO(
        \mult_22/CARRYB[7][32] ), .S(\mult_22/SUMB[7][32] ) );
  FA_X1 \mult_22/S2_7_31  ( .A(\mult_22/ab[7][31] ), .B(
        \mult_22/CARRYB[6][31] ), .CI(\mult_22/SUMB[6][32] ), .CO(
        \mult_22/CARRYB[7][31] ), .S(\mult_22/SUMB[7][31] ) );
  FA_X1 \mult_22/S2_7_30  ( .A(\mult_22/ab[7][30] ), .B(
        \mult_22/CARRYB[6][30] ), .CI(\mult_22/SUMB[6][31] ), .CO(
        \mult_22/CARRYB[7][30] ), .S(\mult_22/SUMB[7][30] ) );
  FA_X1 \mult_22/S2_7_29  ( .A(\mult_22/ab[7][29] ), .B(
        \mult_22/CARRYB[6][29] ), .CI(\mult_22/SUMB[6][30] ), .CO(
        \mult_22/CARRYB[7][29] ), .S(\mult_22/SUMB[7][29] ) );
  FA_X1 \mult_22/S2_7_28  ( .A(\mult_22/ab[7][28] ), .B(
        \mult_22/CARRYB[6][28] ), .CI(\mult_22/SUMB[6][29] ), .CO(
        \mult_22/CARRYB[7][28] ), .S(\mult_22/SUMB[7][28] ) );
  FA_X1 \mult_22/S2_7_27  ( .A(\mult_22/ab[7][27] ), .B(
        \mult_22/CARRYB[6][27] ), .CI(\mult_22/SUMB[6][28] ), .CO(
        \mult_22/CARRYB[7][27] ), .S(\mult_22/SUMB[7][27] ) );
  FA_X1 \mult_22/S2_7_26  ( .A(\mult_22/ab[7][26] ), .B(
        \mult_22/CARRYB[6][26] ), .CI(\mult_22/SUMB[6][27] ), .CO(
        \mult_22/CARRYB[7][26] ), .S(\mult_22/SUMB[7][26] ) );
  FA_X1 \mult_22/S2_7_25  ( .A(\mult_22/ab[7][25] ), .B(
        \mult_22/CARRYB[6][25] ), .CI(\mult_22/SUMB[6][26] ), .CO(
        \mult_22/CARRYB[7][25] ), .S(\mult_22/SUMB[7][25] ) );
  FA_X1 \mult_22/S2_7_24  ( .A(\mult_22/ab[7][24] ), .B(
        \mult_22/CARRYB[6][24] ), .CI(\mult_22/SUMB[6][25] ), .CO(
        \mult_22/CARRYB[7][24] ), .S(\mult_22/SUMB[7][24] ) );
  FA_X1 \mult_22/S2_7_23  ( .A(\mult_22/ab[7][23] ), .B(
        \mult_22/CARRYB[6][23] ), .CI(\mult_22/SUMB[6][24] ), .CO(
        \mult_22/CARRYB[7][23] ), .S(\mult_22/SUMB[7][23] ) );
  FA_X1 \mult_22/S2_7_22  ( .A(\mult_22/ab[7][22] ), .B(
        \mult_22/CARRYB[6][22] ), .CI(\mult_22/SUMB[6][23] ), .CO(
        \mult_22/CARRYB[7][22] ), .S(\mult_22/SUMB[7][22] ) );
  FA_X1 \mult_22/S2_7_21  ( .A(\mult_22/ab[7][21] ), .B(
        \mult_22/CARRYB[6][21] ), .CI(\mult_22/SUMB[6][22] ), .CO(
        \mult_22/CARRYB[7][21] ), .S(\mult_22/SUMB[7][21] ) );
  FA_X1 \mult_22/S2_7_20  ( .A(\mult_22/ab[7][20] ), .B(
        \mult_22/CARRYB[6][20] ), .CI(\mult_22/SUMB[6][21] ), .CO(
        \mult_22/CARRYB[7][20] ), .S(\mult_22/SUMB[7][20] ) );
  FA_X1 \mult_22/S2_7_19  ( .A(\mult_22/ab[7][19] ), .B(
        \mult_22/CARRYB[6][19] ), .CI(\mult_22/SUMB[6][20] ), .CO(
        \mult_22/CARRYB[7][19] ), .S(\mult_22/SUMB[7][19] ) );
  FA_X1 \mult_22/S2_7_18  ( .A(\mult_22/ab[7][18] ), .B(
        \mult_22/CARRYB[6][18] ), .CI(\mult_22/SUMB[6][19] ), .CO(
        \mult_22/CARRYB[7][18] ), .S(\mult_22/SUMB[7][18] ) );
  FA_X1 \mult_22/S2_7_17  ( .A(\mult_22/ab[7][17] ), .B(
        \mult_22/CARRYB[6][17] ), .CI(\mult_22/SUMB[6][18] ), .CO(
        \mult_22/CARRYB[7][17] ), .S(\mult_22/SUMB[7][17] ) );
  FA_X1 \mult_22/S2_7_16  ( .A(\mult_22/ab[7][16] ), .B(
        \mult_22/CARRYB[6][16] ), .CI(\mult_22/SUMB[6][17] ), .CO(
        \mult_22/CARRYB[7][16] ), .S(\mult_22/SUMB[7][16] ) );
  FA_X1 \mult_22/S2_7_15  ( .A(\mult_22/ab[7][15] ), .B(
        \mult_22/CARRYB[6][15] ), .CI(\mult_22/SUMB[6][16] ), .CO(
        \mult_22/CARRYB[7][15] ), .S(\mult_22/SUMB[7][15] ) );
  FA_X1 \mult_22/S2_7_14  ( .A(\mult_22/ab[7][14] ), .B(
        \mult_22/CARRYB[6][14] ), .CI(\mult_22/SUMB[6][15] ), .CO(
        \mult_22/CARRYB[7][14] ), .S(\mult_22/SUMB[7][14] ) );
  FA_X1 \mult_22/S2_7_13  ( .A(\mult_22/ab[7][13] ), .B(
        \mult_22/CARRYB[6][13] ), .CI(\mult_22/SUMB[6][14] ), .CO(
        \mult_22/CARRYB[7][13] ), .S(\mult_22/SUMB[7][13] ) );
  FA_X1 \mult_22/S2_7_12  ( .A(\mult_22/ab[7][12] ), .B(
        \mult_22/CARRYB[6][12] ), .CI(\mult_22/SUMB[6][13] ), .CO(
        \mult_22/CARRYB[7][12] ), .S(\mult_22/SUMB[7][12] ) );
  FA_X1 \mult_22/S2_7_11  ( .A(\mult_22/ab[7][11] ), .B(
        \mult_22/CARRYB[6][11] ), .CI(\mult_22/SUMB[6][12] ), .CO(
        \mult_22/CARRYB[7][11] ), .S(\mult_22/SUMB[7][11] ) );
  FA_X1 \mult_22/S2_7_10  ( .A(\mult_22/ab[7][10] ), .B(
        \mult_22/CARRYB[6][10] ), .CI(\mult_22/SUMB[6][11] ), .CO(
        \mult_22/CARRYB[7][10] ), .S(\mult_22/SUMB[7][10] ) );
  FA_X1 \mult_22/S2_7_9  ( .A(\mult_22/ab[7][9] ), .B(\mult_22/CARRYB[6][9] ), 
        .CI(\mult_22/SUMB[6][10] ), .CO(\mult_22/CARRYB[7][9] ), .S(
        \mult_22/SUMB[7][9] ) );
  FA_X1 \mult_22/S2_7_8  ( .A(\mult_22/ab[7][8] ), .B(\mult_22/CARRYB[6][8] ), 
        .CI(\mult_22/SUMB[6][9] ), .CO(\mult_22/CARRYB[7][8] ), .S(
        \mult_22/SUMB[7][8] ) );
  FA_X1 \mult_22/S2_7_7  ( .A(\mult_22/ab[7][7] ), .B(\mult_22/CARRYB[6][7] ), 
        .CI(\mult_22/SUMB[6][8] ), .CO(\mult_22/CARRYB[7][7] ), .S(
        \mult_22/SUMB[7][7] ) );
  FA_X1 \mult_22/S2_7_6  ( .A(\mult_22/ab[7][6] ), .B(\mult_22/CARRYB[6][6] ), 
        .CI(\mult_22/SUMB[6][7] ), .CO(\mult_22/CARRYB[7][6] ), .S(
        \mult_22/SUMB[7][6] ) );
  FA_X1 \mult_22/S2_7_5  ( .A(\mult_22/ab[7][5] ), .B(\mult_22/CARRYB[6][5] ), 
        .CI(\mult_22/SUMB[6][6] ), .CO(\mult_22/CARRYB[7][5] ), .S(
        \mult_22/SUMB[7][5] ) );
  FA_X1 \mult_22/S2_7_4  ( .A(\mult_22/ab[7][4] ), .B(\mult_22/CARRYB[6][4] ), 
        .CI(\mult_22/SUMB[6][5] ), .CO(\mult_22/CARRYB[7][4] ), .S(
        \mult_22/SUMB[7][4] ) );
  FA_X1 \mult_22/S2_7_3  ( .A(\mult_22/ab[7][3] ), .B(\mult_22/CARRYB[6][3] ), 
        .CI(\mult_22/SUMB[6][4] ), .CO(\mult_22/CARRYB[7][3] ), .S(
        \mult_22/SUMB[7][3] ) );
  FA_X1 \mult_22/S2_7_2  ( .A(\mult_22/ab[7][2] ), .B(\mult_22/CARRYB[6][2] ), 
        .CI(\mult_22/SUMB[6][3] ), .CO(\mult_22/CARRYB[7][2] ), .S(
        \mult_22/SUMB[7][2] ) );
  FA_X1 \mult_22/S2_7_1  ( .A(\mult_22/ab[7][1] ), .B(\mult_22/CARRYB[6][1] ), 
        .CI(\mult_22/SUMB[6][2] ), .CO(\mult_22/CARRYB[7][1] ), .S(
        \mult_22/SUMB[7][1] ) );
  FA_X1 \mult_22/S1_7_0  ( .A(\mult_22/ab[7][0] ), .B(\mult_22/CARRYB[6][0] ), 
        .CI(\mult_22/SUMB[6][1] ), .CO(\mult_22/CARRYB[7][0] ), .S(N135) );
  FA_X1 \mult_22/S3_8_62  ( .A(\mult_22/ab[8][62] ), .B(
        \mult_22/CARRYB[7][62] ), .CI(\mult_22/ab[7][63] ), .CO(
        \mult_22/CARRYB[8][62] ), .S(\mult_22/SUMB[8][62] ) );
  FA_X1 \mult_22/S2_8_61  ( .A(\mult_22/ab[8][61] ), .B(
        \mult_22/CARRYB[7][61] ), .CI(\mult_22/SUMB[7][62] ), .CO(
        \mult_22/CARRYB[8][61] ), .S(\mult_22/SUMB[8][61] ) );
  FA_X1 \mult_22/S2_8_60  ( .A(\mult_22/ab[8][60] ), .B(
        \mult_22/CARRYB[7][60] ), .CI(\mult_22/SUMB[7][61] ), .CO(
        \mult_22/CARRYB[8][60] ), .S(\mult_22/SUMB[8][60] ) );
  FA_X1 \mult_22/S2_8_59  ( .A(\mult_22/ab[8][59] ), .B(
        \mult_22/CARRYB[7][59] ), .CI(\mult_22/SUMB[7][60] ), .CO(
        \mult_22/CARRYB[8][59] ), .S(\mult_22/SUMB[8][59] ) );
  FA_X1 \mult_22/S2_8_58  ( .A(\mult_22/CARRYB[7][58] ), .B(
        \mult_22/ab[8][58] ), .CI(\mult_22/SUMB[7][59] ), .CO(
        \mult_22/CARRYB[8][58] ), .S(\mult_22/SUMB[8][58] ) );
  FA_X1 \mult_22/S2_8_57  ( .A(\mult_22/CARRYB[7][57] ), .B(
        \mult_22/ab[8][57] ), .CI(\mult_22/SUMB[7][58] ), .CO(
        \mult_22/CARRYB[8][57] ), .S(\mult_22/SUMB[8][57] ) );
  FA_X1 \mult_22/S2_8_56  ( .A(\mult_22/CARRYB[7][56] ), .B(
        \mult_22/ab[8][56] ), .CI(\mult_22/SUMB[7][57] ), .CO(
        \mult_22/CARRYB[8][56] ), .S(\mult_22/SUMB[8][56] ) );
  FA_X1 \mult_22/S2_8_55  ( .A(\mult_22/ab[8][55] ), .B(
        \mult_22/CARRYB[7][55] ), .CI(\mult_22/SUMB[7][56] ), .CO(
        \mult_22/CARRYB[8][55] ), .S(\mult_22/SUMB[8][55] ) );
  FA_X1 \mult_22/S2_8_54  ( .A(\mult_22/ab[8][54] ), .B(
        \mult_22/CARRYB[7][54] ), .CI(\mult_22/SUMB[7][55] ), .CO(
        \mult_22/CARRYB[8][54] ), .S(\mult_22/SUMB[8][54] ) );
  FA_X1 \mult_22/S2_8_53  ( .A(\mult_22/CARRYB[7][53] ), .B(
        \mult_22/ab[8][53] ), .CI(\mult_22/SUMB[7][54] ), .CO(
        \mult_22/CARRYB[8][53] ), .S(\mult_22/SUMB[8][53] ) );
  FA_X1 \mult_22/S2_8_52  ( .A(\mult_22/ab[8][52] ), .B(
        \mult_22/CARRYB[7][52] ), .CI(\mult_22/SUMB[7][53] ), .CO(
        \mult_22/CARRYB[8][52] ), .S(\mult_22/SUMB[8][52] ) );
  FA_X1 \mult_22/S2_8_51  ( .A(\mult_22/ab[8][51] ), .B(
        \mult_22/CARRYB[7][51] ), .CI(\mult_22/SUMB[7][52] ), .CO(
        \mult_22/CARRYB[8][51] ), .S(\mult_22/SUMB[8][51] ) );
  FA_X1 \mult_22/S2_8_49  ( .A(\mult_22/ab[8][49] ), .B(
        \mult_22/CARRYB[7][49] ), .CI(\mult_22/SUMB[7][50] ), .CO(
        \mult_22/CARRYB[8][49] ), .S(\mult_22/SUMB[8][49] ) );
  FA_X1 \mult_22/S2_8_48  ( .A(\mult_22/ab[8][48] ), .B(
        \mult_22/CARRYB[7][48] ), .CI(\mult_22/SUMB[7][49] ), .CO(
        \mult_22/CARRYB[8][48] ), .S(\mult_22/SUMB[8][48] ) );
  FA_X1 \mult_22/S2_8_47  ( .A(\mult_22/ab[8][47] ), .B(
        \mult_22/CARRYB[7][47] ), .CI(\mult_22/SUMB[7][48] ), .CO(
        \mult_22/CARRYB[8][47] ), .S(\mult_22/SUMB[8][47] ) );
  FA_X1 \mult_22/S2_8_46  ( .A(\mult_22/ab[8][46] ), .B(
        \mult_22/CARRYB[7][46] ), .CI(\mult_22/SUMB[7][47] ), .CO(
        \mult_22/CARRYB[8][46] ), .S(\mult_22/SUMB[8][46] ) );
  FA_X1 \mult_22/S2_8_45  ( .A(\mult_22/ab[8][45] ), .B(
        \mult_22/CARRYB[7][45] ), .CI(\mult_22/SUMB[7][46] ), .CO(
        \mult_22/CARRYB[8][45] ), .S(\mult_22/SUMB[8][45] ) );
  FA_X1 \mult_22/S2_8_44  ( .A(\mult_22/ab[8][44] ), .B(
        \mult_22/CARRYB[7][44] ), .CI(\mult_22/SUMB[7][45] ), .CO(
        \mult_22/CARRYB[8][44] ), .S(\mult_22/SUMB[8][44] ) );
  FA_X1 \mult_22/S2_8_43  ( .A(\mult_22/ab[8][43] ), .B(
        \mult_22/CARRYB[7][43] ), .CI(\mult_22/SUMB[7][44] ), .CO(
        \mult_22/CARRYB[8][43] ), .S(\mult_22/SUMB[8][43] ) );
  FA_X1 \mult_22/S2_8_42  ( .A(\mult_22/ab[8][42] ), .B(
        \mult_22/CARRYB[7][42] ), .CI(\mult_22/SUMB[7][43] ), .CO(
        \mult_22/CARRYB[8][42] ), .S(\mult_22/SUMB[8][42] ) );
  FA_X1 \mult_22/S2_8_41  ( .A(\mult_22/ab[8][41] ), .B(
        \mult_22/CARRYB[7][41] ), .CI(\mult_22/SUMB[7][42] ), .CO(
        \mult_22/CARRYB[8][41] ), .S(\mult_22/SUMB[8][41] ) );
  FA_X1 \mult_22/S2_8_40  ( .A(\mult_22/ab[8][40] ), .B(
        \mult_22/CARRYB[7][40] ), .CI(\mult_22/SUMB[7][41] ), .CO(
        \mult_22/CARRYB[8][40] ), .S(\mult_22/SUMB[8][40] ) );
  FA_X1 \mult_22/S2_8_39  ( .A(\mult_22/ab[8][39] ), .B(
        \mult_22/CARRYB[7][39] ), .CI(\mult_22/SUMB[7][40] ), .CO(
        \mult_22/CARRYB[8][39] ), .S(\mult_22/SUMB[8][39] ) );
  FA_X1 \mult_22/S2_8_38  ( .A(\mult_22/ab[8][38] ), .B(
        \mult_22/CARRYB[7][38] ), .CI(\mult_22/SUMB[7][39] ), .CO(
        \mult_22/CARRYB[8][38] ), .S(\mult_22/SUMB[8][38] ) );
  FA_X1 \mult_22/S2_8_37  ( .A(\mult_22/ab[8][37] ), .B(
        \mult_22/CARRYB[7][37] ), .CI(\mult_22/SUMB[7][38] ), .CO(
        \mult_22/CARRYB[8][37] ), .S(\mult_22/SUMB[8][37] ) );
  FA_X1 \mult_22/S2_8_36  ( .A(\mult_22/ab[8][36] ), .B(
        \mult_22/CARRYB[7][36] ), .CI(\mult_22/SUMB[7][37] ), .CO(
        \mult_22/CARRYB[8][36] ), .S(\mult_22/SUMB[8][36] ) );
  FA_X1 \mult_22/S2_8_35  ( .A(\mult_22/ab[8][35] ), .B(
        \mult_22/CARRYB[7][35] ), .CI(\mult_22/SUMB[7][36] ), .CO(
        \mult_22/CARRYB[8][35] ), .S(\mult_22/SUMB[8][35] ) );
  FA_X1 \mult_22/S2_8_34  ( .A(\mult_22/ab[8][34] ), .B(
        \mult_22/CARRYB[7][34] ), .CI(\mult_22/SUMB[7][35] ), .CO(
        \mult_22/CARRYB[8][34] ), .S(\mult_22/SUMB[8][34] ) );
  FA_X1 \mult_22/S2_8_33  ( .A(\mult_22/ab[8][33] ), .B(
        \mult_22/CARRYB[7][33] ), .CI(\mult_22/SUMB[7][34] ), .CO(
        \mult_22/CARRYB[8][33] ), .S(\mult_22/SUMB[8][33] ) );
  FA_X1 \mult_22/S2_8_32  ( .A(\mult_22/ab[8][32] ), .B(
        \mult_22/CARRYB[7][32] ), .CI(\mult_22/SUMB[7][33] ), .CO(
        \mult_22/CARRYB[8][32] ), .S(\mult_22/SUMB[8][32] ) );
  FA_X1 \mult_22/S2_8_31  ( .A(\mult_22/ab[8][31] ), .B(
        \mult_22/CARRYB[7][31] ), .CI(\mult_22/SUMB[7][32] ), .CO(
        \mult_22/CARRYB[8][31] ), .S(\mult_22/SUMB[8][31] ) );
  FA_X1 \mult_22/S2_8_30  ( .A(\mult_22/ab[8][30] ), .B(
        \mult_22/CARRYB[7][30] ), .CI(\mult_22/SUMB[7][31] ), .CO(
        \mult_22/CARRYB[8][30] ), .S(\mult_22/SUMB[8][30] ) );
  FA_X1 \mult_22/S2_8_29  ( .A(\mult_22/ab[8][29] ), .B(
        \mult_22/CARRYB[7][29] ), .CI(\mult_22/SUMB[7][30] ), .CO(
        \mult_22/CARRYB[8][29] ), .S(\mult_22/SUMB[8][29] ) );
  FA_X1 \mult_22/S2_8_28  ( .A(\mult_22/ab[8][28] ), .B(
        \mult_22/CARRYB[7][28] ), .CI(\mult_22/SUMB[7][29] ), .CO(
        \mult_22/CARRYB[8][28] ), .S(\mult_22/SUMB[8][28] ) );
  FA_X1 \mult_22/S2_8_27  ( .A(\mult_22/ab[8][27] ), .B(
        \mult_22/CARRYB[7][27] ), .CI(\mult_22/SUMB[7][28] ), .CO(
        \mult_22/CARRYB[8][27] ), .S(\mult_22/SUMB[8][27] ) );
  FA_X1 \mult_22/S2_8_26  ( .A(\mult_22/ab[8][26] ), .B(
        \mult_22/CARRYB[7][26] ), .CI(\mult_22/SUMB[7][27] ), .CO(
        \mult_22/CARRYB[8][26] ), .S(\mult_22/SUMB[8][26] ) );
  FA_X1 \mult_22/S2_8_25  ( .A(\mult_22/ab[8][25] ), .B(
        \mult_22/CARRYB[7][25] ), .CI(\mult_22/SUMB[7][26] ), .CO(
        \mult_22/CARRYB[8][25] ), .S(\mult_22/SUMB[8][25] ) );
  FA_X1 \mult_22/S2_8_24  ( .A(\mult_22/ab[8][24] ), .B(
        \mult_22/CARRYB[7][24] ), .CI(\mult_22/SUMB[7][25] ), .CO(
        \mult_22/CARRYB[8][24] ), .S(\mult_22/SUMB[8][24] ) );
  FA_X1 \mult_22/S2_8_23  ( .A(\mult_22/ab[8][23] ), .B(
        \mult_22/CARRYB[7][23] ), .CI(\mult_22/SUMB[7][24] ), .CO(
        \mult_22/CARRYB[8][23] ), .S(\mult_22/SUMB[8][23] ) );
  FA_X1 \mult_22/S2_8_22  ( .A(\mult_22/ab[8][22] ), .B(
        \mult_22/CARRYB[7][22] ), .CI(\mult_22/SUMB[7][23] ), .CO(
        \mult_22/CARRYB[8][22] ), .S(\mult_22/SUMB[8][22] ) );
  FA_X1 \mult_22/S2_8_21  ( .A(\mult_22/ab[8][21] ), .B(
        \mult_22/CARRYB[7][21] ), .CI(\mult_22/SUMB[7][22] ), .CO(
        \mult_22/CARRYB[8][21] ), .S(\mult_22/SUMB[8][21] ) );
  FA_X1 \mult_22/S2_8_20  ( .A(\mult_22/ab[8][20] ), .B(
        \mult_22/CARRYB[7][20] ), .CI(\mult_22/SUMB[7][21] ), .CO(
        \mult_22/CARRYB[8][20] ), .S(\mult_22/SUMB[8][20] ) );
  FA_X1 \mult_22/S2_8_19  ( .A(\mult_22/ab[8][19] ), .B(
        \mult_22/CARRYB[7][19] ), .CI(\mult_22/SUMB[7][20] ), .CO(
        \mult_22/CARRYB[8][19] ), .S(\mult_22/SUMB[8][19] ) );
  FA_X1 \mult_22/S2_8_18  ( .A(\mult_22/ab[8][18] ), .B(
        \mult_22/CARRYB[7][18] ), .CI(\mult_22/SUMB[7][19] ), .CO(
        \mult_22/CARRYB[8][18] ), .S(\mult_22/SUMB[8][18] ) );
  FA_X1 \mult_22/S2_8_17  ( .A(\mult_22/ab[8][17] ), .B(
        \mult_22/CARRYB[7][17] ), .CI(\mult_22/SUMB[7][18] ), .CO(
        \mult_22/CARRYB[8][17] ), .S(\mult_22/SUMB[8][17] ) );
  FA_X1 \mult_22/S2_8_16  ( .A(\mult_22/ab[8][16] ), .B(
        \mult_22/CARRYB[7][16] ), .CI(\mult_22/SUMB[7][17] ), .CO(
        \mult_22/CARRYB[8][16] ), .S(\mult_22/SUMB[8][16] ) );
  FA_X1 \mult_22/S2_8_15  ( .A(\mult_22/ab[8][15] ), .B(
        \mult_22/CARRYB[7][15] ), .CI(\mult_22/SUMB[7][16] ), .CO(
        \mult_22/CARRYB[8][15] ), .S(\mult_22/SUMB[8][15] ) );
  FA_X1 \mult_22/S2_8_14  ( .A(\mult_22/ab[8][14] ), .B(
        \mult_22/CARRYB[7][14] ), .CI(\mult_22/SUMB[7][15] ), .CO(
        \mult_22/CARRYB[8][14] ), .S(\mult_22/SUMB[8][14] ) );
  FA_X1 \mult_22/S2_8_13  ( .A(\mult_22/ab[8][13] ), .B(
        \mult_22/CARRYB[7][13] ), .CI(\mult_22/SUMB[7][14] ), .CO(
        \mult_22/CARRYB[8][13] ), .S(\mult_22/SUMB[8][13] ) );
  FA_X1 \mult_22/S2_8_12  ( .A(\mult_22/ab[8][12] ), .B(
        \mult_22/CARRYB[7][12] ), .CI(\mult_22/SUMB[7][13] ), .CO(
        \mult_22/CARRYB[8][12] ), .S(\mult_22/SUMB[8][12] ) );
  FA_X1 \mult_22/S2_8_11  ( .A(\mult_22/ab[8][11] ), .B(
        \mult_22/CARRYB[7][11] ), .CI(\mult_22/SUMB[7][12] ), .CO(
        \mult_22/CARRYB[8][11] ), .S(\mult_22/SUMB[8][11] ) );
  FA_X1 \mult_22/S2_8_10  ( .A(\mult_22/ab[8][10] ), .B(
        \mult_22/CARRYB[7][10] ), .CI(\mult_22/SUMB[7][11] ), .CO(
        \mult_22/CARRYB[8][10] ), .S(\mult_22/SUMB[8][10] ) );
  FA_X1 \mult_22/S2_8_9  ( .A(\mult_22/ab[8][9] ), .B(\mult_22/CARRYB[7][9] ), 
        .CI(\mult_22/SUMB[7][10] ), .CO(\mult_22/CARRYB[8][9] ), .S(
        \mult_22/SUMB[8][9] ) );
  FA_X1 \mult_22/S2_8_8  ( .A(\mult_22/ab[8][8] ), .B(\mult_22/CARRYB[7][8] ), 
        .CI(\mult_22/SUMB[7][9] ), .CO(\mult_22/CARRYB[8][8] ), .S(
        \mult_22/SUMB[8][8] ) );
  FA_X1 \mult_22/S2_8_7  ( .A(\mult_22/ab[8][7] ), .B(\mult_22/CARRYB[7][7] ), 
        .CI(\mult_22/SUMB[7][8] ), .CO(\mult_22/CARRYB[8][7] ), .S(
        \mult_22/SUMB[8][7] ) );
  FA_X1 \mult_22/S2_8_6  ( .A(\mult_22/ab[8][6] ), .B(\mult_22/CARRYB[7][6] ), 
        .CI(\mult_22/SUMB[7][7] ), .CO(\mult_22/CARRYB[8][6] ), .S(
        \mult_22/SUMB[8][6] ) );
  FA_X1 \mult_22/S2_8_5  ( .A(\mult_22/ab[8][5] ), .B(\mult_22/CARRYB[7][5] ), 
        .CI(\mult_22/SUMB[7][6] ), .CO(\mult_22/CARRYB[8][5] ), .S(
        \mult_22/SUMB[8][5] ) );
  FA_X1 \mult_22/S2_8_4  ( .A(\mult_22/ab[8][4] ), .B(\mult_22/CARRYB[7][4] ), 
        .CI(\mult_22/SUMB[7][5] ), .CO(\mult_22/CARRYB[8][4] ), .S(
        \mult_22/SUMB[8][4] ) );
  FA_X1 \mult_22/S2_8_3  ( .A(\mult_22/ab[8][3] ), .B(\mult_22/CARRYB[7][3] ), 
        .CI(\mult_22/SUMB[7][4] ), .CO(\mult_22/CARRYB[8][3] ), .S(
        \mult_22/SUMB[8][3] ) );
  FA_X1 \mult_22/S2_8_2  ( .A(\mult_22/ab[8][2] ), .B(\mult_22/CARRYB[7][2] ), 
        .CI(\mult_22/SUMB[7][3] ), .CO(\mult_22/CARRYB[8][2] ), .S(
        \mult_22/SUMB[8][2] ) );
  FA_X1 \mult_22/S2_8_1  ( .A(\mult_22/ab[8][1] ), .B(\mult_22/CARRYB[7][1] ), 
        .CI(\mult_22/SUMB[7][2] ), .CO(\mult_22/CARRYB[8][1] ), .S(
        \mult_22/SUMB[8][1] ) );
  FA_X1 \mult_22/S1_8_0  ( .A(\mult_22/ab[8][0] ), .B(\mult_22/CARRYB[7][0] ), 
        .CI(\mult_22/SUMB[7][1] ), .CO(\mult_22/CARRYB[8][0] ), .S(N136) );
  FA_X1 \mult_22/S3_9_62  ( .A(\mult_22/ab[9][62] ), .B(
        \mult_22/CARRYB[8][62] ), .CI(\mult_22/ab[8][63] ), .CO(
        \mult_22/CARRYB[9][62] ), .S(\mult_22/SUMB[9][62] ) );
  FA_X1 \mult_22/S2_9_61  ( .A(\mult_22/ab[9][61] ), .B(
        \mult_22/CARRYB[8][61] ), .CI(\mult_22/SUMB[8][62] ), .CO(
        \mult_22/CARRYB[9][61] ), .S(\mult_22/SUMB[9][61] ) );
  FA_X1 \mult_22/S2_9_60  ( .A(\mult_22/ab[9][60] ), .B(
        \mult_22/CARRYB[8][60] ), .CI(\mult_22/SUMB[8][61] ), .CO(
        \mult_22/CARRYB[9][60] ), .S(\mult_22/SUMB[9][60] ) );
  FA_X1 \mult_22/S2_9_59  ( .A(\mult_22/ab[9][59] ), .B(
        \mult_22/CARRYB[8][59] ), .CI(\mult_22/SUMB[8][60] ), .CO(
        \mult_22/CARRYB[9][59] ), .S(\mult_22/SUMB[9][59] ) );
  FA_X1 \mult_22/S2_9_58  ( .A(\mult_22/CARRYB[8][58] ), .B(
        \mult_22/ab[9][58] ), .CI(\mult_22/SUMB[8][59] ), .CO(
        \mult_22/CARRYB[9][58] ), .S(\mult_22/SUMB[9][58] ) );
  FA_X1 \mult_22/S2_9_57  ( .A(\mult_22/ab[9][57] ), .B(
        \mult_22/CARRYB[8][57] ), .CI(\mult_22/SUMB[8][58] ), .CO(
        \mult_22/CARRYB[9][57] ), .S(\mult_22/SUMB[9][57] ) );
  FA_X1 \mult_22/S2_9_56  ( .A(\mult_22/CARRYB[8][56] ), .B(
        \mult_22/ab[9][56] ), .CI(\mult_22/SUMB[8][57] ), .CO(
        \mult_22/CARRYB[9][56] ), .S(\mult_22/SUMB[9][56] ) );
  FA_X1 \mult_22/S2_9_55  ( .A(\mult_22/CARRYB[8][55] ), .B(
        \mult_22/ab[9][55] ), .CI(\mult_22/SUMB[8][56] ), .CO(
        \mult_22/CARRYB[9][55] ), .S(\mult_22/SUMB[9][55] ) );
  FA_X1 \mult_22/S2_9_54  ( .A(\mult_22/ab[9][54] ), .B(
        \mult_22/CARRYB[8][54] ), .CI(\mult_22/SUMB[8][55] ), .CO(
        \mult_22/CARRYB[9][54] ), .S(\mult_22/SUMB[9][54] ) );
  FA_X1 \mult_22/S2_9_53  ( .A(\mult_22/ab[9][53] ), .B(
        \mult_22/CARRYB[8][53] ), .CI(\mult_22/SUMB[8][54] ), .CO(
        \mult_22/CARRYB[9][53] ), .S(\mult_22/SUMB[9][53] ) );
  FA_X1 \mult_22/S2_9_52  ( .A(\mult_22/ab[9][52] ), .B(
        \mult_22/CARRYB[8][52] ), .CI(\mult_22/SUMB[8][53] ), .CO(
        \mult_22/CARRYB[9][52] ), .S(\mult_22/SUMB[9][52] ) );
  FA_X1 \mult_22/S2_9_49  ( .A(\mult_22/ab[9][49] ), .B(
        \mult_22/CARRYB[8][49] ), .CI(\mult_22/SUMB[8][50] ), .CO(
        \mult_22/CARRYB[9][49] ), .S(\mult_22/SUMB[9][49] ) );
  FA_X1 \mult_22/S2_9_48  ( .A(\mult_22/ab[9][48] ), .B(
        \mult_22/CARRYB[8][48] ), .CI(\mult_22/SUMB[8][49] ), .CO(
        \mult_22/CARRYB[9][48] ), .S(\mult_22/SUMB[9][48] ) );
  FA_X1 \mult_22/S2_9_47  ( .A(\mult_22/ab[9][47] ), .B(
        \mult_22/CARRYB[8][47] ), .CI(\mult_22/SUMB[8][48] ), .CO(
        \mult_22/CARRYB[9][47] ), .S(\mult_22/SUMB[9][47] ) );
  FA_X1 \mult_22/S2_9_46  ( .A(\mult_22/ab[9][46] ), .B(
        \mult_22/CARRYB[8][46] ), .CI(\mult_22/SUMB[8][47] ), .CO(
        \mult_22/CARRYB[9][46] ), .S(\mult_22/SUMB[9][46] ) );
  FA_X1 \mult_22/S2_9_45  ( .A(\mult_22/ab[9][45] ), .B(
        \mult_22/CARRYB[8][45] ), .CI(\mult_22/SUMB[8][46] ), .CO(
        \mult_22/CARRYB[9][45] ), .S(\mult_22/SUMB[9][45] ) );
  FA_X1 \mult_22/S2_9_44  ( .A(\mult_22/ab[9][44] ), .B(
        \mult_22/CARRYB[8][44] ), .CI(\mult_22/SUMB[8][45] ), .CO(
        \mult_22/CARRYB[9][44] ), .S(\mult_22/SUMB[9][44] ) );
  FA_X1 \mult_22/S2_9_43  ( .A(\mult_22/ab[9][43] ), .B(
        \mult_22/CARRYB[8][43] ), .CI(\mult_22/SUMB[8][44] ), .CO(
        \mult_22/CARRYB[9][43] ), .S(\mult_22/SUMB[9][43] ) );
  FA_X1 \mult_22/S2_9_42  ( .A(\mult_22/ab[9][42] ), .B(
        \mult_22/CARRYB[8][42] ), .CI(\mult_22/SUMB[8][43] ), .CO(
        \mult_22/CARRYB[9][42] ), .S(\mult_22/SUMB[9][42] ) );
  FA_X1 \mult_22/S2_9_41  ( .A(\mult_22/ab[9][41] ), .B(
        \mult_22/CARRYB[8][41] ), .CI(\mult_22/SUMB[8][42] ), .CO(
        \mult_22/CARRYB[9][41] ), .S(\mult_22/SUMB[9][41] ) );
  FA_X1 \mult_22/S2_9_40  ( .A(\mult_22/ab[9][40] ), .B(
        \mult_22/CARRYB[8][40] ), .CI(\mult_22/SUMB[8][41] ), .CO(
        \mult_22/CARRYB[9][40] ), .S(\mult_22/SUMB[9][40] ) );
  FA_X1 \mult_22/S2_9_39  ( .A(\mult_22/ab[9][39] ), .B(
        \mult_22/CARRYB[8][39] ), .CI(\mult_22/SUMB[8][40] ), .CO(
        \mult_22/CARRYB[9][39] ), .S(\mult_22/SUMB[9][39] ) );
  FA_X1 \mult_22/S2_9_38  ( .A(\mult_22/ab[9][38] ), .B(
        \mult_22/CARRYB[8][38] ), .CI(\mult_22/SUMB[8][39] ), .CO(
        \mult_22/CARRYB[9][38] ), .S(\mult_22/SUMB[9][38] ) );
  FA_X1 \mult_22/S2_9_37  ( .A(\mult_22/ab[9][37] ), .B(
        \mult_22/CARRYB[8][37] ), .CI(\mult_22/SUMB[8][38] ), .CO(
        \mult_22/CARRYB[9][37] ), .S(\mult_22/SUMB[9][37] ) );
  FA_X1 \mult_22/S2_9_36  ( .A(\mult_22/ab[9][36] ), .B(
        \mult_22/CARRYB[8][36] ), .CI(\mult_22/SUMB[8][37] ), .CO(
        \mult_22/CARRYB[9][36] ), .S(\mult_22/SUMB[9][36] ) );
  FA_X1 \mult_22/S2_9_35  ( .A(\mult_22/ab[9][35] ), .B(
        \mult_22/CARRYB[8][35] ), .CI(\mult_22/SUMB[8][36] ), .CO(
        \mult_22/CARRYB[9][35] ), .S(\mult_22/SUMB[9][35] ) );
  FA_X1 \mult_22/S2_9_34  ( .A(\mult_22/ab[9][34] ), .B(
        \mult_22/CARRYB[8][34] ), .CI(\mult_22/SUMB[8][35] ), .CO(
        \mult_22/CARRYB[9][34] ), .S(\mult_22/SUMB[9][34] ) );
  FA_X1 \mult_22/S2_9_33  ( .A(\mult_22/ab[9][33] ), .B(
        \mult_22/CARRYB[8][33] ), .CI(\mult_22/SUMB[8][34] ), .CO(
        \mult_22/CARRYB[9][33] ), .S(\mult_22/SUMB[9][33] ) );
  FA_X1 \mult_22/S2_9_32  ( .A(\mult_22/ab[9][32] ), .B(
        \mult_22/CARRYB[8][32] ), .CI(\mult_22/SUMB[8][33] ), .CO(
        \mult_22/CARRYB[9][32] ), .S(\mult_22/SUMB[9][32] ) );
  FA_X1 \mult_22/S2_9_31  ( .A(\mult_22/ab[9][31] ), .B(
        \mult_22/CARRYB[8][31] ), .CI(\mult_22/SUMB[8][32] ), .CO(
        \mult_22/CARRYB[9][31] ), .S(\mult_22/SUMB[9][31] ) );
  FA_X1 \mult_22/S2_9_30  ( .A(\mult_22/ab[9][30] ), .B(
        \mult_22/CARRYB[8][30] ), .CI(\mult_22/SUMB[8][31] ), .CO(
        \mult_22/CARRYB[9][30] ), .S(\mult_22/SUMB[9][30] ) );
  FA_X1 \mult_22/S2_9_29  ( .A(\mult_22/ab[9][29] ), .B(
        \mult_22/CARRYB[8][29] ), .CI(\mult_22/SUMB[8][30] ), .CO(
        \mult_22/CARRYB[9][29] ), .S(\mult_22/SUMB[9][29] ) );
  FA_X1 \mult_22/S2_9_28  ( .A(\mult_22/ab[9][28] ), .B(
        \mult_22/CARRYB[8][28] ), .CI(\mult_22/SUMB[8][29] ), .CO(
        \mult_22/CARRYB[9][28] ), .S(\mult_22/SUMB[9][28] ) );
  FA_X1 \mult_22/S2_9_27  ( .A(\mult_22/ab[9][27] ), .B(
        \mult_22/CARRYB[8][27] ), .CI(\mult_22/SUMB[8][28] ), .CO(
        \mult_22/CARRYB[9][27] ), .S(\mult_22/SUMB[9][27] ) );
  FA_X1 \mult_22/S2_9_26  ( .A(\mult_22/ab[9][26] ), .B(
        \mult_22/CARRYB[8][26] ), .CI(\mult_22/SUMB[8][27] ), .CO(
        \mult_22/CARRYB[9][26] ), .S(\mult_22/SUMB[9][26] ) );
  FA_X1 \mult_22/S2_9_25  ( .A(\mult_22/ab[9][25] ), .B(
        \mult_22/CARRYB[8][25] ), .CI(\mult_22/SUMB[8][26] ), .CO(
        \mult_22/CARRYB[9][25] ), .S(\mult_22/SUMB[9][25] ) );
  FA_X1 \mult_22/S2_9_24  ( .A(\mult_22/ab[9][24] ), .B(
        \mult_22/CARRYB[8][24] ), .CI(\mult_22/SUMB[8][25] ), .CO(
        \mult_22/CARRYB[9][24] ), .S(\mult_22/SUMB[9][24] ) );
  FA_X1 \mult_22/S2_9_23  ( .A(\mult_22/ab[9][23] ), .B(
        \mult_22/CARRYB[8][23] ), .CI(\mult_22/SUMB[8][24] ), .CO(
        \mult_22/CARRYB[9][23] ), .S(\mult_22/SUMB[9][23] ) );
  FA_X1 \mult_22/S2_9_22  ( .A(\mult_22/ab[9][22] ), .B(
        \mult_22/CARRYB[8][22] ), .CI(\mult_22/SUMB[8][23] ), .CO(
        \mult_22/CARRYB[9][22] ), .S(\mult_22/SUMB[9][22] ) );
  FA_X1 \mult_22/S2_9_21  ( .A(\mult_22/ab[9][21] ), .B(
        \mult_22/CARRYB[8][21] ), .CI(\mult_22/SUMB[8][22] ), .CO(
        \mult_22/CARRYB[9][21] ), .S(\mult_22/SUMB[9][21] ) );
  FA_X1 \mult_22/S2_9_20  ( .A(\mult_22/ab[9][20] ), .B(
        \mult_22/CARRYB[8][20] ), .CI(\mult_22/SUMB[8][21] ), .CO(
        \mult_22/CARRYB[9][20] ), .S(\mult_22/SUMB[9][20] ) );
  FA_X1 \mult_22/S2_9_19  ( .A(\mult_22/ab[9][19] ), .B(
        \mult_22/CARRYB[8][19] ), .CI(\mult_22/SUMB[8][20] ), .CO(
        \mult_22/CARRYB[9][19] ), .S(\mult_22/SUMB[9][19] ) );
  FA_X1 \mult_22/S2_9_18  ( .A(\mult_22/ab[9][18] ), .B(
        \mult_22/CARRYB[8][18] ), .CI(\mult_22/SUMB[8][19] ), .CO(
        \mult_22/CARRYB[9][18] ), .S(\mult_22/SUMB[9][18] ) );
  FA_X1 \mult_22/S2_9_17  ( .A(\mult_22/ab[9][17] ), .B(
        \mult_22/CARRYB[8][17] ), .CI(\mult_22/SUMB[8][18] ), .CO(
        \mult_22/CARRYB[9][17] ), .S(\mult_22/SUMB[9][17] ) );
  FA_X1 \mult_22/S2_9_16  ( .A(\mult_22/ab[9][16] ), .B(
        \mult_22/CARRYB[8][16] ), .CI(\mult_22/SUMB[8][17] ), .CO(
        \mult_22/CARRYB[9][16] ), .S(\mult_22/SUMB[9][16] ) );
  FA_X1 \mult_22/S2_9_15  ( .A(\mult_22/ab[9][15] ), .B(
        \mult_22/CARRYB[8][15] ), .CI(\mult_22/SUMB[8][16] ), .CO(
        \mult_22/CARRYB[9][15] ), .S(\mult_22/SUMB[9][15] ) );
  FA_X1 \mult_22/S2_9_14  ( .A(\mult_22/ab[9][14] ), .B(
        \mult_22/CARRYB[8][14] ), .CI(\mult_22/SUMB[8][15] ), .CO(
        \mult_22/CARRYB[9][14] ), .S(\mult_22/SUMB[9][14] ) );
  FA_X1 \mult_22/S2_9_13  ( .A(\mult_22/ab[9][13] ), .B(
        \mult_22/CARRYB[8][13] ), .CI(\mult_22/SUMB[8][14] ), .CO(
        \mult_22/CARRYB[9][13] ), .S(\mult_22/SUMB[9][13] ) );
  FA_X1 \mult_22/S2_9_12  ( .A(\mult_22/ab[9][12] ), .B(
        \mult_22/CARRYB[8][12] ), .CI(\mult_22/SUMB[8][13] ), .CO(
        \mult_22/CARRYB[9][12] ), .S(\mult_22/SUMB[9][12] ) );
  FA_X1 \mult_22/S2_9_11  ( .A(\mult_22/ab[9][11] ), .B(
        \mult_22/CARRYB[8][11] ), .CI(\mult_22/SUMB[8][12] ), .CO(
        \mult_22/CARRYB[9][11] ), .S(\mult_22/SUMB[9][11] ) );
  FA_X1 \mult_22/S2_9_10  ( .A(\mult_22/ab[9][10] ), .B(
        \mult_22/CARRYB[8][10] ), .CI(\mult_22/SUMB[8][11] ), .CO(
        \mult_22/CARRYB[9][10] ), .S(\mult_22/SUMB[9][10] ) );
  FA_X1 \mult_22/S2_9_9  ( .A(\mult_22/ab[9][9] ), .B(\mult_22/CARRYB[8][9] ), 
        .CI(\mult_22/SUMB[8][10] ), .CO(\mult_22/CARRYB[9][9] ), .S(
        \mult_22/SUMB[9][9] ) );
  FA_X1 \mult_22/S2_9_8  ( .A(\mult_22/ab[9][8] ), .B(\mult_22/CARRYB[8][8] ), 
        .CI(\mult_22/SUMB[8][9] ), .CO(\mult_22/CARRYB[9][8] ), .S(
        \mult_22/SUMB[9][8] ) );
  FA_X1 \mult_22/S2_9_7  ( .A(\mult_22/ab[9][7] ), .B(\mult_22/CARRYB[8][7] ), 
        .CI(\mult_22/SUMB[8][8] ), .CO(\mult_22/CARRYB[9][7] ), .S(
        \mult_22/SUMB[9][7] ) );
  FA_X1 \mult_22/S2_9_6  ( .A(\mult_22/ab[9][6] ), .B(\mult_22/CARRYB[8][6] ), 
        .CI(\mult_22/SUMB[8][7] ), .CO(\mult_22/CARRYB[9][6] ), .S(
        \mult_22/SUMB[9][6] ) );
  FA_X1 \mult_22/S2_9_5  ( .A(\mult_22/ab[9][5] ), .B(\mult_22/CARRYB[8][5] ), 
        .CI(\mult_22/SUMB[8][6] ), .CO(\mult_22/CARRYB[9][5] ), .S(
        \mult_22/SUMB[9][5] ) );
  FA_X1 \mult_22/S2_9_4  ( .A(\mult_22/ab[9][4] ), .B(\mult_22/CARRYB[8][4] ), 
        .CI(\mult_22/SUMB[8][5] ), .CO(\mult_22/CARRYB[9][4] ), .S(
        \mult_22/SUMB[9][4] ) );
  FA_X1 \mult_22/S2_9_3  ( .A(\mult_22/ab[9][3] ), .B(\mult_22/CARRYB[8][3] ), 
        .CI(\mult_22/SUMB[8][4] ), .CO(\mult_22/CARRYB[9][3] ), .S(
        \mult_22/SUMB[9][3] ) );
  FA_X1 \mult_22/S2_9_2  ( .A(\mult_22/ab[9][2] ), .B(\mult_22/CARRYB[8][2] ), 
        .CI(\mult_22/SUMB[8][3] ), .CO(\mult_22/CARRYB[9][2] ), .S(
        \mult_22/SUMB[9][2] ) );
  FA_X1 \mult_22/S2_9_1  ( .A(\mult_22/ab[9][1] ), .B(\mult_22/CARRYB[8][1] ), 
        .CI(\mult_22/SUMB[8][2] ), .CO(\mult_22/CARRYB[9][1] ), .S(
        \mult_22/SUMB[9][1] ) );
  FA_X1 \mult_22/S1_9_0  ( .A(\mult_22/ab[9][0] ), .B(\mult_22/CARRYB[8][0] ), 
        .CI(\mult_22/SUMB[8][1] ), .CO(\mult_22/CARRYB[9][0] ), .S(N137) );
  FA_X1 \mult_22/S3_10_62  ( .A(\mult_22/ab[10][62] ), .B(
        \mult_22/CARRYB[9][62] ), .CI(\mult_22/ab[9][63] ), .CO(
        \mult_22/CARRYB[10][62] ), .S(\mult_22/SUMB[10][62] ) );
  FA_X1 \mult_22/S2_10_61  ( .A(\mult_22/ab[10][61] ), .B(
        \mult_22/CARRYB[9][61] ), .CI(\mult_22/SUMB[9][62] ), .CO(
        \mult_22/CARRYB[10][61] ), .S(\mult_22/SUMB[10][61] ) );
  FA_X1 \mult_22/S2_10_60  ( .A(\mult_22/ab[10][60] ), .B(
        \mult_22/CARRYB[9][60] ), .CI(\mult_22/SUMB[9][61] ), .CO(
        \mult_22/CARRYB[10][60] ), .S(\mult_22/SUMB[10][60] ) );
  FA_X1 \mult_22/S2_10_59  ( .A(\mult_22/ab[10][59] ), .B(
        \mult_22/CARRYB[9][59] ), .CI(\mult_22/SUMB[9][60] ), .CO(
        \mult_22/CARRYB[10][59] ), .S(\mult_22/SUMB[10][59] ) );
  FA_X1 \mult_22/S2_10_58  ( .A(\mult_22/ab[10][58] ), .B(
        \mult_22/CARRYB[9][58] ), .CI(\mult_22/SUMB[9][59] ), .CO(
        \mult_22/CARRYB[10][58] ), .S(\mult_22/SUMB[10][58] ) );
  FA_X1 \mult_22/S2_10_57  ( .A(\mult_22/ab[10][57] ), .B(
        \mult_22/CARRYB[9][57] ), .CI(\mult_22/SUMB[9][58] ), .CO(
        \mult_22/CARRYB[10][57] ), .S(\mult_22/SUMB[10][57] ) );
  FA_X1 \mult_22/S2_10_56  ( .A(\mult_22/CARRYB[9][56] ), .B(
        \mult_22/ab[10][56] ), .CI(\mult_22/SUMB[9][57] ), .CO(
        \mult_22/CARRYB[10][56] ), .S(\mult_22/SUMB[10][56] ) );
  FA_X1 \mult_22/S2_10_55  ( .A(\mult_22/CARRYB[9][55] ), .B(
        \mult_22/ab[10][55] ), .CI(\mult_22/SUMB[9][56] ), .CO(
        \mult_22/CARRYB[10][55] ), .S(\mult_22/SUMB[10][55] ) );
  FA_X1 \mult_22/S2_10_54  ( .A(\mult_22/CARRYB[9][54] ), .B(
        \mult_22/ab[10][54] ), .CI(\mult_22/SUMB[9][55] ), .CO(
        \mult_22/CARRYB[10][54] ), .S(\mult_22/SUMB[10][54] ) );
  FA_X1 \mult_22/S2_10_53  ( .A(\mult_22/ab[10][53] ), .B(
        \mult_22/CARRYB[9][53] ), .CI(\mult_22/SUMB[9][54] ), .CO(
        \mult_22/CARRYB[10][53] ), .S(\mult_22/SUMB[10][53] ) );
  FA_X1 \mult_22/S2_10_52  ( .A(\mult_22/ab[10][52] ), .B(
        \mult_22/CARRYB[9][52] ), .CI(\mult_22/SUMB[9][53] ), .CO(
        \mult_22/CARRYB[10][52] ), .S(\mult_22/SUMB[10][52] ) );
  FA_X1 \mult_22/S2_10_51  ( .A(\mult_22/ab[10][51] ), .B(
        \mult_22/CARRYB[9][51] ), .CI(\mult_22/SUMB[9][52] ), .CO(
        \mult_22/CARRYB[10][51] ), .S(\mult_22/SUMB[10][51] ) );
  FA_X1 \mult_22/S2_10_50  ( .A(\mult_22/ab[10][50] ), .B(
        \mult_22/CARRYB[9][50] ), .CI(\mult_22/SUMB[9][51] ), .CO(
        \mult_22/CARRYB[10][50] ), .S(\mult_22/SUMB[10][50] ) );
  FA_X1 \mult_22/S2_10_49  ( .A(\mult_22/ab[10][49] ), .B(
        \mult_22/CARRYB[9][49] ), .CI(\mult_22/SUMB[9][50] ), .CO(
        \mult_22/CARRYB[10][49] ), .S(\mult_22/SUMB[10][49] ) );
  FA_X1 \mult_22/S2_10_48  ( .A(\mult_22/ab[10][48] ), .B(
        \mult_22/CARRYB[9][48] ), .CI(\mult_22/SUMB[9][49] ), .CO(
        \mult_22/CARRYB[10][48] ), .S(\mult_22/SUMB[10][48] ) );
  FA_X1 \mult_22/S2_10_47  ( .A(\mult_22/ab[10][47] ), .B(
        \mult_22/CARRYB[9][47] ), .CI(\mult_22/SUMB[9][48] ), .CO(
        \mult_22/CARRYB[10][47] ), .S(\mult_22/SUMB[10][47] ) );
  FA_X1 \mult_22/S2_10_46  ( .A(\mult_22/ab[10][46] ), .B(
        \mult_22/CARRYB[9][46] ), .CI(\mult_22/SUMB[9][47] ), .CO(
        \mult_22/CARRYB[10][46] ), .S(\mult_22/SUMB[10][46] ) );
  FA_X1 \mult_22/S2_10_45  ( .A(\mult_22/ab[10][45] ), .B(
        \mult_22/CARRYB[9][45] ), .CI(\mult_22/SUMB[9][46] ), .CO(
        \mult_22/CARRYB[10][45] ), .S(\mult_22/SUMB[10][45] ) );
  FA_X1 \mult_22/S2_10_44  ( .A(\mult_22/ab[10][44] ), .B(
        \mult_22/CARRYB[9][44] ), .CI(\mult_22/SUMB[9][45] ), .CO(
        \mult_22/CARRYB[10][44] ), .S(\mult_22/SUMB[10][44] ) );
  FA_X1 \mult_22/S2_10_43  ( .A(\mult_22/ab[10][43] ), .B(
        \mult_22/CARRYB[9][43] ), .CI(\mult_22/SUMB[9][44] ), .CO(
        \mult_22/CARRYB[10][43] ), .S(\mult_22/SUMB[10][43] ) );
  FA_X1 \mult_22/S2_10_42  ( .A(\mult_22/ab[10][42] ), .B(
        \mult_22/CARRYB[9][42] ), .CI(\mult_22/SUMB[9][43] ), .CO(
        \mult_22/CARRYB[10][42] ), .S(\mult_22/SUMB[10][42] ) );
  FA_X1 \mult_22/S2_10_41  ( .A(\mult_22/ab[10][41] ), .B(
        \mult_22/CARRYB[9][41] ), .CI(\mult_22/SUMB[9][42] ), .CO(
        \mult_22/CARRYB[10][41] ), .S(\mult_22/SUMB[10][41] ) );
  FA_X1 \mult_22/S2_10_40  ( .A(\mult_22/ab[10][40] ), .B(
        \mult_22/CARRYB[9][40] ), .CI(\mult_22/SUMB[9][41] ), .CO(
        \mult_22/CARRYB[10][40] ), .S(\mult_22/SUMB[10][40] ) );
  FA_X1 \mult_22/S2_10_39  ( .A(\mult_22/ab[10][39] ), .B(
        \mult_22/CARRYB[9][39] ), .CI(\mult_22/SUMB[9][40] ), .CO(
        \mult_22/CARRYB[10][39] ), .S(\mult_22/SUMB[10][39] ) );
  FA_X1 \mult_22/S2_10_38  ( .A(\mult_22/ab[10][38] ), .B(
        \mult_22/CARRYB[9][38] ), .CI(\mult_22/SUMB[9][39] ), .CO(
        \mult_22/CARRYB[10][38] ), .S(\mult_22/SUMB[10][38] ) );
  FA_X1 \mult_22/S2_10_37  ( .A(\mult_22/ab[10][37] ), .B(
        \mult_22/CARRYB[9][37] ), .CI(\mult_22/SUMB[9][38] ), .CO(
        \mult_22/CARRYB[10][37] ), .S(\mult_22/SUMB[10][37] ) );
  FA_X1 \mult_22/S2_10_36  ( .A(\mult_22/ab[10][36] ), .B(
        \mult_22/CARRYB[9][36] ), .CI(\mult_22/SUMB[9][37] ), .CO(
        \mult_22/CARRYB[10][36] ), .S(\mult_22/SUMB[10][36] ) );
  FA_X1 \mult_22/S2_10_35  ( .A(\mult_22/ab[10][35] ), .B(
        \mult_22/CARRYB[9][35] ), .CI(\mult_22/SUMB[9][36] ), .CO(
        \mult_22/CARRYB[10][35] ), .S(\mult_22/SUMB[10][35] ) );
  FA_X1 \mult_22/S2_10_34  ( .A(\mult_22/ab[10][34] ), .B(
        \mult_22/CARRYB[9][34] ), .CI(\mult_22/SUMB[9][35] ), .CO(
        \mult_22/CARRYB[10][34] ), .S(\mult_22/SUMB[10][34] ) );
  FA_X1 \mult_22/S2_10_33  ( .A(\mult_22/ab[10][33] ), .B(
        \mult_22/CARRYB[9][33] ), .CI(\mult_22/SUMB[9][34] ), .CO(
        \mult_22/CARRYB[10][33] ), .S(\mult_22/SUMB[10][33] ) );
  FA_X1 \mult_22/S2_10_32  ( .A(\mult_22/ab[10][32] ), .B(
        \mult_22/CARRYB[9][32] ), .CI(\mult_22/SUMB[9][33] ), .CO(
        \mult_22/CARRYB[10][32] ), .S(\mult_22/SUMB[10][32] ) );
  FA_X1 \mult_22/S2_10_31  ( .A(\mult_22/ab[10][31] ), .B(
        \mult_22/CARRYB[9][31] ), .CI(\mult_22/SUMB[9][32] ), .CO(
        \mult_22/CARRYB[10][31] ), .S(\mult_22/SUMB[10][31] ) );
  FA_X1 \mult_22/S2_10_30  ( .A(\mult_22/ab[10][30] ), .B(
        \mult_22/CARRYB[9][30] ), .CI(\mult_22/SUMB[9][31] ), .CO(
        \mult_22/CARRYB[10][30] ), .S(\mult_22/SUMB[10][30] ) );
  FA_X1 \mult_22/S2_10_29  ( .A(\mult_22/ab[10][29] ), .B(
        \mult_22/CARRYB[9][29] ), .CI(\mult_22/SUMB[9][30] ), .CO(
        \mult_22/CARRYB[10][29] ), .S(\mult_22/SUMB[10][29] ) );
  FA_X1 \mult_22/S2_10_28  ( .A(\mult_22/ab[10][28] ), .B(
        \mult_22/CARRYB[9][28] ), .CI(\mult_22/SUMB[9][29] ), .CO(
        \mult_22/CARRYB[10][28] ), .S(\mult_22/SUMB[10][28] ) );
  FA_X1 \mult_22/S2_10_27  ( .A(\mult_22/ab[10][27] ), .B(
        \mult_22/CARRYB[9][27] ), .CI(\mult_22/SUMB[9][28] ), .CO(
        \mult_22/CARRYB[10][27] ), .S(\mult_22/SUMB[10][27] ) );
  FA_X1 \mult_22/S2_10_26  ( .A(\mult_22/ab[10][26] ), .B(
        \mult_22/CARRYB[9][26] ), .CI(\mult_22/SUMB[9][27] ), .CO(
        \mult_22/CARRYB[10][26] ), .S(\mult_22/SUMB[10][26] ) );
  FA_X1 \mult_22/S2_10_25  ( .A(\mult_22/ab[10][25] ), .B(
        \mult_22/CARRYB[9][25] ), .CI(\mult_22/SUMB[9][26] ), .CO(
        \mult_22/CARRYB[10][25] ), .S(\mult_22/SUMB[10][25] ) );
  FA_X1 \mult_22/S2_10_24  ( .A(\mult_22/ab[10][24] ), .B(
        \mult_22/CARRYB[9][24] ), .CI(\mult_22/SUMB[9][25] ), .CO(
        \mult_22/CARRYB[10][24] ), .S(\mult_22/SUMB[10][24] ) );
  FA_X1 \mult_22/S2_10_23  ( .A(\mult_22/ab[10][23] ), .B(
        \mult_22/CARRYB[9][23] ), .CI(\mult_22/SUMB[9][24] ), .CO(
        \mult_22/CARRYB[10][23] ), .S(\mult_22/SUMB[10][23] ) );
  FA_X1 \mult_22/S2_10_22  ( .A(\mult_22/ab[10][22] ), .B(
        \mult_22/CARRYB[9][22] ), .CI(\mult_22/SUMB[9][23] ), .CO(
        \mult_22/CARRYB[10][22] ), .S(\mult_22/SUMB[10][22] ) );
  FA_X1 \mult_22/S2_10_21  ( .A(\mult_22/ab[10][21] ), .B(
        \mult_22/CARRYB[9][21] ), .CI(\mult_22/SUMB[9][22] ), .CO(
        \mult_22/CARRYB[10][21] ), .S(\mult_22/SUMB[10][21] ) );
  FA_X1 \mult_22/S2_10_20  ( .A(\mult_22/ab[10][20] ), .B(
        \mult_22/CARRYB[9][20] ), .CI(\mult_22/SUMB[9][21] ), .CO(
        \mult_22/CARRYB[10][20] ), .S(\mult_22/SUMB[10][20] ) );
  FA_X1 \mult_22/S2_10_19  ( .A(\mult_22/ab[10][19] ), .B(
        \mult_22/CARRYB[9][19] ), .CI(\mult_22/SUMB[9][20] ), .CO(
        \mult_22/CARRYB[10][19] ), .S(\mult_22/SUMB[10][19] ) );
  FA_X1 \mult_22/S2_10_18  ( .A(\mult_22/ab[10][18] ), .B(
        \mult_22/CARRYB[9][18] ), .CI(\mult_22/SUMB[9][19] ), .CO(
        \mult_22/CARRYB[10][18] ), .S(\mult_22/SUMB[10][18] ) );
  FA_X1 \mult_22/S2_10_17  ( .A(\mult_22/ab[10][17] ), .B(
        \mult_22/CARRYB[9][17] ), .CI(\mult_22/SUMB[9][18] ), .CO(
        \mult_22/CARRYB[10][17] ), .S(\mult_22/SUMB[10][17] ) );
  FA_X1 \mult_22/S2_10_16  ( .A(\mult_22/ab[10][16] ), .B(
        \mult_22/CARRYB[9][16] ), .CI(\mult_22/SUMB[9][17] ), .CO(
        \mult_22/CARRYB[10][16] ), .S(\mult_22/SUMB[10][16] ) );
  FA_X1 \mult_22/S2_10_15  ( .A(\mult_22/ab[10][15] ), .B(
        \mult_22/CARRYB[9][15] ), .CI(\mult_22/SUMB[9][16] ), .CO(
        \mult_22/CARRYB[10][15] ), .S(\mult_22/SUMB[10][15] ) );
  FA_X1 \mult_22/S2_10_14  ( .A(\mult_22/ab[10][14] ), .B(
        \mult_22/CARRYB[9][14] ), .CI(\mult_22/SUMB[9][15] ), .CO(
        \mult_22/CARRYB[10][14] ), .S(\mult_22/SUMB[10][14] ) );
  FA_X1 \mult_22/S2_10_13  ( .A(\mult_22/ab[10][13] ), .B(
        \mult_22/CARRYB[9][13] ), .CI(\mult_22/SUMB[9][14] ), .CO(
        \mult_22/CARRYB[10][13] ), .S(\mult_22/SUMB[10][13] ) );
  FA_X1 \mult_22/S2_10_12  ( .A(\mult_22/ab[10][12] ), .B(
        \mult_22/CARRYB[9][12] ), .CI(\mult_22/SUMB[9][13] ), .CO(
        \mult_22/CARRYB[10][12] ), .S(\mult_22/SUMB[10][12] ) );
  FA_X1 \mult_22/S2_10_11  ( .A(\mult_22/ab[10][11] ), .B(
        \mult_22/CARRYB[9][11] ), .CI(\mult_22/SUMB[9][12] ), .CO(
        \mult_22/CARRYB[10][11] ), .S(\mult_22/SUMB[10][11] ) );
  FA_X1 \mult_22/S2_10_10  ( .A(\mult_22/ab[10][10] ), .B(
        \mult_22/CARRYB[9][10] ), .CI(\mult_22/SUMB[9][11] ), .CO(
        \mult_22/CARRYB[10][10] ), .S(\mult_22/SUMB[10][10] ) );
  FA_X1 \mult_22/S2_10_9  ( .A(\mult_22/ab[10][9] ), .B(\mult_22/CARRYB[9][9] ), .CI(\mult_22/SUMB[9][10] ), .CO(\mult_22/CARRYB[10][9] ), .S(
        \mult_22/SUMB[10][9] ) );
  FA_X1 \mult_22/S2_10_8  ( .A(\mult_22/ab[10][8] ), .B(\mult_22/CARRYB[9][8] ), .CI(\mult_22/SUMB[9][9] ), .CO(\mult_22/CARRYB[10][8] ), .S(
        \mult_22/SUMB[10][8] ) );
  FA_X1 \mult_22/S2_10_7  ( .A(\mult_22/ab[10][7] ), .B(\mult_22/CARRYB[9][7] ), .CI(\mult_22/SUMB[9][8] ), .CO(\mult_22/CARRYB[10][7] ), .S(
        \mult_22/SUMB[10][7] ) );
  FA_X1 \mult_22/S2_10_6  ( .A(\mult_22/ab[10][6] ), .B(\mult_22/CARRYB[9][6] ), .CI(\mult_22/SUMB[9][7] ), .CO(\mult_22/CARRYB[10][6] ), .S(
        \mult_22/SUMB[10][6] ) );
  FA_X1 \mult_22/S2_10_5  ( .A(\mult_22/ab[10][5] ), .B(\mult_22/CARRYB[9][5] ), .CI(\mult_22/SUMB[9][6] ), .CO(\mult_22/CARRYB[10][5] ), .S(
        \mult_22/SUMB[10][5] ) );
  FA_X1 \mult_22/S2_10_4  ( .A(\mult_22/ab[10][4] ), .B(\mult_22/CARRYB[9][4] ), .CI(\mult_22/SUMB[9][5] ), .CO(\mult_22/CARRYB[10][4] ), .S(
        \mult_22/SUMB[10][4] ) );
  FA_X1 \mult_22/S2_10_3  ( .A(\mult_22/ab[10][3] ), .B(\mult_22/CARRYB[9][3] ), .CI(\mult_22/SUMB[9][4] ), .CO(\mult_22/CARRYB[10][3] ), .S(
        \mult_22/SUMB[10][3] ) );
  FA_X1 \mult_22/S2_10_2  ( .A(\mult_22/ab[10][2] ), .B(\mult_22/CARRYB[9][2] ), .CI(\mult_22/SUMB[9][3] ), .CO(\mult_22/CARRYB[10][2] ), .S(
        \mult_22/SUMB[10][2] ) );
  FA_X1 \mult_22/S2_10_1  ( .A(\mult_22/ab[10][1] ), .B(\mult_22/CARRYB[9][1] ), .CI(\mult_22/SUMB[9][2] ), .CO(\mult_22/CARRYB[10][1] ), .S(
        \mult_22/SUMB[10][1] ) );
  FA_X1 \mult_22/S1_10_0  ( .A(\mult_22/ab[10][0] ), .B(\mult_22/CARRYB[9][0] ), .CI(\mult_22/SUMB[9][1] ), .CO(\mult_22/CARRYB[10][0] ), .S(N138) );
  FA_X1 \mult_22/S3_11_62  ( .A(\mult_22/ab[11][62] ), .B(
        \mult_22/CARRYB[10][62] ), .CI(\mult_22/ab[10][63] ), .CO(
        \mult_22/CARRYB[11][62] ), .S(\mult_22/SUMB[11][62] ) );
  FA_X1 \mult_22/S2_11_61  ( .A(\mult_22/ab[11][61] ), .B(
        \mult_22/CARRYB[10][61] ), .CI(\mult_22/SUMB[10][62] ), .CO(
        \mult_22/CARRYB[11][61] ), .S(\mult_22/SUMB[11][61] ) );
  FA_X1 \mult_22/S2_11_60  ( .A(\mult_22/ab[11][60] ), .B(
        \mult_22/CARRYB[10][60] ), .CI(\mult_22/SUMB[10][61] ), .CO(
        \mult_22/CARRYB[11][60] ), .S(\mult_22/SUMB[11][60] ) );
  FA_X1 \mult_22/S2_11_59  ( .A(\mult_22/ab[11][59] ), .B(
        \mult_22/CARRYB[10][59] ), .CI(\mult_22/SUMB[10][60] ), .CO(
        \mult_22/CARRYB[11][59] ), .S(\mult_22/SUMB[11][59] ) );
  FA_X1 \mult_22/S2_11_58  ( .A(\mult_22/ab[11][58] ), .B(
        \mult_22/CARRYB[10][58] ), .CI(\mult_22/SUMB[10][59] ), .CO(
        \mult_22/CARRYB[11][58] ), .S(\mult_22/SUMB[11][58] ) );
  FA_X1 \mult_22/S2_11_57  ( .A(\mult_22/ab[11][57] ), .B(
        \mult_22/CARRYB[10][57] ), .CI(\mult_22/SUMB[10][58] ), .CO(
        \mult_22/CARRYB[11][57] ), .S(\mult_22/SUMB[11][57] ) );
  FA_X1 \mult_22/S2_11_56  ( .A(\mult_22/CARRYB[10][56] ), .B(
        \mult_22/ab[11][56] ), .CI(\mult_22/SUMB[10][57] ), .CO(
        \mult_22/CARRYB[11][56] ), .S(\mult_22/SUMB[11][56] ) );
  FA_X1 \mult_22/S2_11_55  ( .A(\mult_22/ab[11][55] ), .B(
        \mult_22/CARRYB[10][55] ), .CI(\mult_22/SUMB[10][56] ), .CO(
        \mult_22/CARRYB[11][55] ), .S(\mult_22/SUMB[11][55] ) );
  FA_X1 \mult_22/S2_11_54  ( .A(\mult_22/CARRYB[10][54] ), .B(
        \mult_22/ab[11][54] ), .CI(\mult_22/SUMB[10][55] ), .CO(
        \mult_22/CARRYB[11][54] ), .S(\mult_22/SUMB[11][54] ) );
  FA_X1 \mult_22/S2_11_53  ( .A(\mult_22/CARRYB[10][53] ), .B(
        \mult_22/ab[11][53] ), .CI(\mult_22/SUMB[10][54] ), .CO(
        \mult_22/CARRYB[11][53] ), .S(\mult_22/SUMB[11][53] ) );
  FA_X1 \mult_22/S2_11_52  ( .A(\mult_22/ab[11][52] ), .B(
        \mult_22/CARRYB[10][52] ), .CI(\mult_22/SUMB[10][53] ), .CO(
        \mult_22/CARRYB[11][52] ), .S(\mult_22/SUMB[11][52] ) );
  FA_X1 \mult_22/S2_11_51  ( .A(\mult_22/ab[11][51] ), .B(
        \mult_22/CARRYB[10][51] ), .CI(\mult_22/SUMB[10][52] ), .CO(
        \mult_22/CARRYB[11][51] ), .S(\mult_22/SUMB[11][51] ) );
  FA_X1 \mult_22/S2_11_50  ( .A(\mult_22/ab[11][50] ), .B(
        \mult_22/CARRYB[10][50] ), .CI(\mult_22/SUMB[10][51] ), .CO(
        \mult_22/CARRYB[11][50] ), .S(\mult_22/SUMB[11][50] ) );
  FA_X1 \mult_22/S2_11_49  ( .A(\mult_22/ab[11][49] ), .B(
        \mult_22/CARRYB[10][49] ), .CI(\mult_22/SUMB[10][50] ), .CO(
        \mult_22/CARRYB[11][49] ), .S(\mult_22/SUMB[11][49] ) );
  FA_X1 \mult_22/S2_11_48  ( .A(\mult_22/ab[11][48] ), .B(
        \mult_22/CARRYB[10][48] ), .CI(\mult_22/SUMB[10][49] ), .CO(
        \mult_22/CARRYB[11][48] ), .S(\mult_22/SUMB[11][48] ) );
  FA_X1 \mult_22/S2_11_45  ( .A(\mult_22/ab[11][45] ), .B(
        \mult_22/CARRYB[10][45] ), .CI(\mult_22/SUMB[10][46] ), .CO(
        \mult_22/CARRYB[11][45] ), .S(\mult_22/SUMB[11][45] ) );
  FA_X1 \mult_22/S2_11_44  ( .A(\mult_22/ab[11][44] ), .B(
        \mult_22/CARRYB[10][44] ), .CI(\mult_22/SUMB[10][45] ), .CO(
        \mult_22/CARRYB[11][44] ), .S(\mult_22/SUMB[11][44] ) );
  FA_X1 \mult_22/S2_11_43  ( .A(\mult_22/ab[11][43] ), .B(
        \mult_22/CARRYB[10][43] ), .CI(\mult_22/SUMB[10][44] ), .CO(
        \mult_22/CARRYB[11][43] ), .S(\mult_22/SUMB[11][43] ) );
  FA_X1 \mult_22/S2_11_42  ( .A(\mult_22/ab[11][42] ), .B(
        \mult_22/CARRYB[10][42] ), .CI(\mult_22/SUMB[10][43] ), .CO(
        \mult_22/CARRYB[11][42] ), .S(\mult_22/SUMB[11][42] ) );
  FA_X1 \mult_22/S2_11_41  ( .A(\mult_22/ab[11][41] ), .B(
        \mult_22/CARRYB[10][41] ), .CI(\mult_22/SUMB[10][42] ), .CO(
        \mult_22/CARRYB[11][41] ), .S(\mult_22/SUMB[11][41] ) );
  FA_X1 \mult_22/S2_11_40  ( .A(\mult_22/ab[11][40] ), .B(
        \mult_22/CARRYB[10][40] ), .CI(\mult_22/SUMB[10][41] ), .CO(
        \mult_22/CARRYB[11][40] ), .S(\mult_22/SUMB[11][40] ) );
  FA_X1 \mult_22/S2_11_39  ( .A(\mult_22/ab[11][39] ), .B(
        \mult_22/CARRYB[10][39] ), .CI(\mult_22/SUMB[10][40] ), .CO(
        \mult_22/CARRYB[11][39] ), .S(\mult_22/SUMB[11][39] ) );
  FA_X1 \mult_22/S2_11_38  ( .A(\mult_22/ab[11][38] ), .B(
        \mult_22/CARRYB[10][38] ), .CI(\mult_22/SUMB[10][39] ), .CO(
        \mult_22/CARRYB[11][38] ), .S(\mult_22/SUMB[11][38] ) );
  FA_X1 \mult_22/S2_11_37  ( .A(\mult_22/ab[11][37] ), .B(
        \mult_22/CARRYB[10][37] ), .CI(\mult_22/SUMB[10][38] ), .CO(
        \mult_22/CARRYB[11][37] ), .S(\mult_22/SUMB[11][37] ) );
  FA_X1 \mult_22/S2_11_36  ( .A(\mult_22/ab[11][36] ), .B(
        \mult_22/CARRYB[10][36] ), .CI(\mult_22/SUMB[10][37] ), .CO(
        \mult_22/CARRYB[11][36] ), .S(\mult_22/SUMB[11][36] ) );
  FA_X1 \mult_22/S2_11_35  ( .A(\mult_22/ab[11][35] ), .B(
        \mult_22/CARRYB[10][35] ), .CI(\mult_22/SUMB[10][36] ), .CO(
        \mult_22/CARRYB[11][35] ), .S(\mult_22/SUMB[11][35] ) );
  FA_X1 \mult_22/S2_11_34  ( .A(\mult_22/ab[11][34] ), .B(
        \mult_22/CARRYB[10][34] ), .CI(\mult_22/SUMB[10][35] ), .CO(
        \mult_22/CARRYB[11][34] ), .S(\mult_22/SUMB[11][34] ) );
  FA_X1 \mult_22/S2_11_33  ( .A(\mult_22/ab[11][33] ), .B(
        \mult_22/CARRYB[10][33] ), .CI(\mult_22/SUMB[10][34] ), .CO(
        \mult_22/CARRYB[11][33] ), .S(\mult_22/SUMB[11][33] ) );
  FA_X1 \mult_22/S2_11_32  ( .A(\mult_22/ab[11][32] ), .B(
        \mult_22/CARRYB[10][32] ), .CI(\mult_22/SUMB[10][33] ), .CO(
        \mult_22/CARRYB[11][32] ), .S(\mult_22/SUMB[11][32] ) );
  FA_X1 \mult_22/S2_11_31  ( .A(\mult_22/ab[11][31] ), .B(
        \mult_22/CARRYB[10][31] ), .CI(\mult_22/SUMB[10][32] ), .CO(
        \mult_22/CARRYB[11][31] ), .S(\mult_22/SUMB[11][31] ) );
  FA_X1 \mult_22/S2_11_30  ( .A(\mult_22/ab[11][30] ), .B(
        \mult_22/CARRYB[10][30] ), .CI(\mult_22/SUMB[10][31] ), .CO(
        \mult_22/CARRYB[11][30] ), .S(\mult_22/SUMB[11][30] ) );
  FA_X1 \mult_22/S2_11_29  ( .A(\mult_22/ab[11][29] ), .B(
        \mult_22/CARRYB[10][29] ), .CI(\mult_22/SUMB[10][30] ), .CO(
        \mult_22/CARRYB[11][29] ), .S(\mult_22/SUMB[11][29] ) );
  FA_X1 \mult_22/S2_11_28  ( .A(\mult_22/ab[11][28] ), .B(
        \mult_22/CARRYB[10][28] ), .CI(\mult_22/SUMB[10][29] ), .CO(
        \mult_22/CARRYB[11][28] ), .S(\mult_22/SUMB[11][28] ) );
  FA_X1 \mult_22/S2_11_27  ( .A(\mult_22/ab[11][27] ), .B(
        \mult_22/CARRYB[10][27] ), .CI(\mult_22/SUMB[10][28] ), .CO(
        \mult_22/CARRYB[11][27] ), .S(\mult_22/SUMB[11][27] ) );
  FA_X1 \mult_22/S2_11_26  ( .A(\mult_22/ab[11][26] ), .B(
        \mult_22/CARRYB[10][26] ), .CI(\mult_22/SUMB[10][27] ), .CO(
        \mult_22/CARRYB[11][26] ), .S(\mult_22/SUMB[11][26] ) );
  FA_X1 \mult_22/S2_11_25  ( .A(\mult_22/ab[11][25] ), .B(
        \mult_22/CARRYB[10][25] ), .CI(\mult_22/SUMB[10][26] ), .CO(
        \mult_22/CARRYB[11][25] ), .S(\mult_22/SUMB[11][25] ) );
  FA_X1 \mult_22/S2_11_24  ( .A(\mult_22/ab[11][24] ), .B(
        \mult_22/CARRYB[10][24] ), .CI(\mult_22/SUMB[10][25] ), .CO(
        \mult_22/CARRYB[11][24] ), .S(\mult_22/SUMB[11][24] ) );
  FA_X1 \mult_22/S2_11_23  ( .A(\mult_22/ab[11][23] ), .B(
        \mult_22/CARRYB[10][23] ), .CI(\mult_22/SUMB[10][24] ), .CO(
        \mult_22/CARRYB[11][23] ), .S(\mult_22/SUMB[11][23] ) );
  FA_X1 \mult_22/S2_11_22  ( .A(\mult_22/ab[11][22] ), .B(
        \mult_22/CARRYB[10][22] ), .CI(\mult_22/SUMB[10][23] ), .CO(
        \mult_22/CARRYB[11][22] ), .S(\mult_22/SUMB[11][22] ) );
  FA_X1 \mult_22/S2_11_21  ( .A(\mult_22/ab[11][21] ), .B(
        \mult_22/CARRYB[10][21] ), .CI(\mult_22/SUMB[10][22] ), .CO(
        \mult_22/CARRYB[11][21] ), .S(\mult_22/SUMB[11][21] ) );
  FA_X1 \mult_22/S2_11_20  ( .A(\mult_22/ab[11][20] ), .B(
        \mult_22/CARRYB[10][20] ), .CI(\mult_22/SUMB[10][21] ), .CO(
        \mult_22/CARRYB[11][20] ), .S(\mult_22/SUMB[11][20] ) );
  FA_X1 \mult_22/S2_11_19  ( .A(\mult_22/ab[11][19] ), .B(
        \mult_22/CARRYB[10][19] ), .CI(\mult_22/SUMB[10][20] ), .CO(
        \mult_22/CARRYB[11][19] ), .S(\mult_22/SUMB[11][19] ) );
  FA_X1 \mult_22/S2_11_18  ( .A(\mult_22/ab[11][18] ), .B(
        \mult_22/CARRYB[10][18] ), .CI(\mult_22/SUMB[10][19] ), .CO(
        \mult_22/CARRYB[11][18] ), .S(\mult_22/SUMB[11][18] ) );
  FA_X1 \mult_22/S2_11_17  ( .A(\mult_22/ab[11][17] ), .B(
        \mult_22/CARRYB[10][17] ), .CI(\mult_22/SUMB[10][18] ), .CO(
        \mult_22/CARRYB[11][17] ), .S(\mult_22/SUMB[11][17] ) );
  FA_X1 \mult_22/S2_11_16  ( .A(\mult_22/ab[11][16] ), .B(
        \mult_22/CARRYB[10][16] ), .CI(\mult_22/SUMB[10][17] ), .CO(
        \mult_22/CARRYB[11][16] ), .S(\mult_22/SUMB[11][16] ) );
  FA_X1 \mult_22/S2_11_15  ( .A(\mult_22/ab[11][15] ), .B(
        \mult_22/CARRYB[10][15] ), .CI(\mult_22/SUMB[10][16] ), .CO(
        \mult_22/CARRYB[11][15] ), .S(\mult_22/SUMB[11][15] ) );
  FA_X1 \mult_22/S2_11_14  ( .A(\mult_22/ab[11][14] ), .B(
        \mult_22/CARRYB[10][14] ), .CI(\mult_22/SUMB[10][15] ), .CO(
        \mult_22/CARRYB[11][14] ), .S(\mult_22/SUMB[11][14] ) );
  FA_X1 \mult_22/S2_11_13  ( .A(\mult_22/ab[11][13] ), .B(
        \mult_22/CARRYB[10][13] ), .CI(\mult_22/SUMB[10][14] ), .CO(
        \mult_22/CARRYB[11][13] ), .S(\mult_22/SUMB[11][13] ) );
  FA_X1 \mult_22/S2_11_12  ( .A(\mult_22/ab[11][12] ), .B(
        \mult_22/CARRYB[10][12] ), .CI(\mult_22/SUMB[10][13] ), .CO(
        \mult_22/CARRYB[11][12] ), .S(\mult_22/SUMB[11][12] ) );
  FA_X1 \mult_22/S2_11_11  ( .A(\mult_22/ab[11][11] ), .B(
        \mult_22/CARRYB[10][11] ), .CI(\mult_22/SUMB[10][12] ), .CO(
        \mult_22/CARRYB[11][11] ), .S(\mult_22/SUMB[11][11] ) );
  FA_X1 \mult_22/S2_11_10  ( .A(\mult_22/ab[11][10] ), .B(
        \mult_22/CARRYB[10][10] ), .CI(\mult_22/SUMB[10][11] ), .CO(
        \mult_22/CARRYB[11][10] ), .S(\mult_22/SUMB[11][10] ) );
  FA_X1 \mult_22/S2_11_9  ( .A(\mult_22/ab[11][9] ), .B(
        \mult_22/CARRYB[10][9] ), .CI(\mult_22/SUMB[10][10] ), .CO(
        \mult_22/CARRYB[11][9] ), .S(\mult_22/SUMB[11][9] ) );
  FA_X1 \mult_22/S2_11_8  ( .A(\mult_22/ab[11][8] ), .B(
        \mult_22/CARRYB[10][8] ), .CI(\mult_22/SUMB[10][9] ), .CO(
        \mult_22/CARRYB[11][8] ), .S(\mult_22/SUMB[11][8] ) );
  FA_X1 \mult_22/S2_11_7  ( .A(\mult_22/ab[11][7] ), .B(
        \mult_22/CARRYB[10][7] ), .CI(\mult_22/SUMB[10][8] ), .CO(
        \mult_22/CARRYB[11][7] ), .S(\mult_22/SUMB[11][7] ) );
  FA_X1 \mult_22/S2_11_6  ( .A(\mult_22/ab[11][6] ), .B(
        \mult_22/CARRYB[10][6] ), .CI(\mult_22/SUMB[10][7] ), .CO(
        \mult_22/CARRYB[11][6] ), .S(\mult_22/SUMB[11][6] ) );
  FA_X1 \mult_22/S2_11_5  ( .A(\mult_22/ab[11][5] ), .B(
        \mult_22/CARRYB[10][5] ), .CI(\mult_22/SUMB[10][6] ), .CO(
        \mult_22/CARRYB[11][5] ), .S(\mult_22/SUMB[11][5] ) );
  FA_X1 \mult_22/S2_11_4  ( .A(\mult_22/ab[11][4] ), .B(
        \mult_22/CARRYB[10][4] ), .CI(\mult_22/SUMB[10][5] ), .CO(
        \mult_22/CARRYB[11][4] ), .S(\mult_22/SUMB[11][4] ) );
  FA_X1 \mult_22/S2_11_3  ( .A(\mult_22/ab[11][3] ), .B(
        \mult_22/CARRYB[10][3] ), .CI(\mult_22/SUMB[10][4] ), .CO(
        \mult_22/CARRYB[11][3] ), .S(\mult_22/SUMB[11][3] ) );
  FA_X1 \mult_22/S2_11_2  ( .A(\mult_22/ab[11][2] ), .B(
        \mult_22/CARRYB[10][2] ), .CI(\mult_22/SUMB[10][3] ), .CO(
        \mult_22/CARRYB[11][2] ), .S(\mult_22/SUMB[11][2] ) );
  FA_X1 \mult_22/S2_11_1  ( .A(\mult_22/ab[11][1] ), .B(
        \mult_22/CARRYB[10][1] ), .CI(\mult_22/SUMB[10][2] ), .CO(
        \mult_22/CARRYB[11][1] ), .S(\mult_22/SUMB[11][1] ) );
  FA_X1 \mult_22/S1_11_0  ( .A(\mult_22/ab[11][0] ), .B(
        \mult_22/CARRYB[10][0] ), .CI(\mult_22/SUMB[10][1] ), .CO(
        \mult_22/CARRYB[11][0] ), .S(N139) );
  FA_X1 \mult_22/S3_12_62  ( .A(\mult_22/ab[12][62] ), .B(
        \mult_22/CARRYB[11][62] ), .CI(\mult_22/ab[11][63] ), .CO(
        \mult_22/CARRYB[12][62] ), .S(\mult_22/SUMB[12][62] ) );
  FA_X1 \mult_22/S2_12_61  ( .A(\mult_22/ab[12][61] ), .B(
        \mult_22/CARRYB[11][61] ), .CI(\mult_22/SUMB[11][62] ), .CO(
        \mult_22/CARRYB[12][61] ), .S(\mult_22/SUMB[12][61] ) );
  FA_X1 \mult_22/S2_12_60  ( .A(\mult_22/ab[12][60] ), .B(
        \mult_22/CARRYB[11][60] ), .CI(\mult_22/SUMB[11][61] ), .CO(
        \mult_22/CARRYB[12][60] ), .S(\mult_22/SUMB[12][60] ) );
  FA_X1 \mult_22/S2_12_59  ( .A(\mult_22/ab[12][59] ), .B(
        \mult_22/CARRYB[11][59] ), .CI(\mult_22/SUMB[11][60] ), .CO(
        \mult_22/CARRYB[12][59] ), .S(\mult_22/SUMB[12][59] ) );
  FA_X1 \mult_22/S2_12_58  ( .A(\mult_22/ab[12][58] ), .B(
        \mult_22/CARRYB[11][58] ), .CI(\mult_22/SUMB[11][59] ), .CO(
        \mult_22/CARRYB[12][58] ), .S(\mult_22/SUMB[12][58] ) );
  FA_X1 \mult_22/S2_12_57  ( .A(\mult_22/ab[12][57] ), .B(
        \mult_22/CARRYB[11][57] ), .CI(\mult_22/SUMB[11][58] ), .CO(
        \mult_22/CARRYB[12][57] ), .S(\mult_22/SUMB[12][57] ) );
  FA_X1 \mult_22/S2_12_56  ( .A(\mult_22/ab[12][56] ), .B(
        \mult_22/CARRYB[11][56] ), .CI(\mult_22/SUMB[11][57] ), .CO(
        \mult_22/CARRYB[12][56] ), .S(\mult_22/SUMB[12][56] ) );
  FA_X1 \mult_22/S2_12_55  ( .A(\mult_22/ab[12][55] ), .B(
        \mult_22/CARRYB[11][55] ), .CI(\mult_22/SUMB[11][56] ), .CO(
        \mult_22/CARRYB[12][55] ), .S(\mult_22/SUMB[12][55] ) );
  FA_X1 \mult_22/S2_12_54  ( .A(\mult_22/CARRYB[11][54] ), .B(
        \mult_22/ab[12][54] ), .CI(\mult_22/SUMB[11][55] ), .CO(
        \mult_22/CARRYB[12][54] ), .S(\mult_22/SUMB[12][54] ) );
  FA_X1 \mult_22/S2_12_53  ( .A(\mult_22/ab[12][53] ), .B(
        \mult_22/CARRYB[11][53] ), .CI(\mult_22/SUMB[11][54] ), .CO(
        \mult_22/CARRYB[12][53] ), .S(\mult_22/SUMB[12][53] ) );
  FA_X1 \mult_22/S2_12_52  ( .A(\mult_22/CARRYB[11][52] ), .B(
        \mult_22/ab[12][52] ), .CI(\mult_22/SUMB[11][53] ), .CO(
        \mult_22/CARRYB[12][52] ), .S(\mult_22/SUMB[12][52] ) );
  FA_X1 \mult_22/S2_12_51  ( .A(\mult_22/ab[12][51] ), .B(
        \mult_22/CARRYB[11][51] ), .CI(\mult_22/SUMB[11][52] ), .CO(
        \mult_22/CARRYB[12][51] ), .S(\mult_22/SUMB[12][51] ) );
  FA_X1 \mult_22/S2_12_50  ( .A(\mult_22/ab[12][50] ), .B(
        \mult_22/CARRYB[11][50] ), .CI(\mult_22/SUMB[11][51] ), .CO(
        \mult_22/CARRYB[12][50] ), .S(\mult_22/SUMB[12][50] ) );
  FA_X1 \mult_22/S2_12_49  ( .A(\mult_22/ab[12][49] ), .B(
        \mult_22/CARRYB[11][49] ), .CI(\mult_22/SUMB[11][50] ), .CO(
        \mult_22/CARRYB[12][49] ), .S(\mult_22/SUMB[12][49] ) );
  FA_X1 \mult_22/S2_12_48  ( .A(\mult_22/ab[12][48] ), .B(
        \mult_22/CARRYB[11][48] ), .CI(\mult_22/SUMB[11][49] ), .CO(
        \mult_22/CARRYB[12][48] ), .S(\mult_22/SUMB[12][48] ) );
  FA_X1 \mult_22/S2_12_47  ( .A(\mult_22/ab[12][47] ), .B(
        \mult_22/CARRYB[11][47] ), .CI(\mult_22/SUMB[11][48] ), .CO(
        \mult_22/CARRYB[12][47] ), .S(\mult_22/SUMB[12][47] ) );
  FA_X1 \mult_22/S2_12_46  ( .A(\mult_22/CARRYB[11][46] ), .B(
        \mult_22/ab[12][46] ), .CI(\mult_22/SUMB[11][47] ), .CO(
        \mult_22/CARRYB[12][46] ), .S(\mult_22/SUMB[12][46] ) );
  FA_X1 \mult_22/S2_12_45  ( .A(\mult_22/ab[12][45] ), .B(
        \mult_22/CARRYB[11][45] ), .CI(\mult_22/SUMB[11][46] ), .CO(
        \mult_22/CARRYB[12][45] ), .S(\mult_22/SUMB[12][45] ) );
  FA_X1 \mult_22/S2_12_44  ( .A(\mult_22/ab[12][44] ), .B(
        \mult_22/CARRYB[11][44] ), .CI(\mult_22/SUMB[11][45] ), .CO(
        \mult_22/CARRYB[12][44] ), .S(\mult_22/SUMB[12][44] ) );
  FA_X1 \mult_22/S2_12_43  ( .A(\mult_22/ab[12][43] ), .B(
        \mult_22/CARRYB[11][43] ), .CI(\mult_22/SUMB[11][44] ), .CO(
        \mult_22/CARRYB[12][43] ), .S(\mult_22/SUMB[12][43] ) );
  FA_X1 \mult_22/S2_12_42  ( .A(\mult_22/ab[12][42] ), .B(
        \mult_22/CARRYB[11][42] ), .CI(\mult_22/SUMB[11][43] ), .CO(
        \mult_22/CARRYB[12][42] ), .S(\mult_22/SUMB[12][42] ) );
  FA_X1 \mult_22/S2_12_41  ( .A(\mult_22/ab[12][41] ), .B(
        \mult_22/CARRYB[11][41] ), .CI(\mult_22/SUMB[11][42] ), .CO(
        \mult_22/CARRYB[12][41] ), .S(\mult_22/SUMB[12][41] ) );
  FA_X1 \mult_22/S2_12_40  ( .A(\mult_22/ab[12][40] ), .B(
        \mult_22/CARRYB[11][40] ), .CI(\mult_22/SUMB[11][41] ), .CO(
        \mult_22/CARRYB[12][40] ), .S(\mult_22/SUMB[12][40] ) );
  FA_X1 \mult_22/S2_12_39  ( .A(\mult_22/ab[12][39] ), .B(
        \mult_22/CARRYB[11][39] ), .CI(\mult_22/SUMB[11][40] ), .CO(
        \mult_22/CARRYB[12][39] ), .S(\mult_22/SUMB[12][39] ) );
  FA_X1 \mult_22/S2_12_38  ( .A(\mult_22/ab[12][38] ), .B(
        \mult_22/CARRYB[11][38] ), .CI(\mult_22/SUMB[11][39] ), .CO(
        \mult_22/CARRYB[12][38] ), .S(\mult_22/SUMB[12][38] ) );
  FA_X1 \mult_22/S2_12_37  ( .A(\mult_22/ab[12][37] ), .B(
        \mult_22/CARRYB[11][37] ), .CI(\mult_22/SUMB[11][38] ), .CO(
        \mult_22/CARRYB[12][37] ), .S(\mult_22/SUMB[12][37] ) );
  FA_X1 \mult_22/S2_12_36  ( .A(\mult_22/ab[12][36] ), .B(
        \mult_22/CARRYB[11][36] ), .CI(\mult_22/SUMB[11][37] ), .CO(
        \mult_22/CARRYB[12][36] ), .S(\mult_22/SUMB[12][36] ) );
  FA_X1 \mult_22/S2_12_35  ( .A(\mult_22/ab[12][35] ), .B(
        \mult_22/CARRYB[11][35] ), .CI(\mult_22/SUMB[11][36] ), .CO(
        \mult_22/CARRYB[12][35] ), .S(\mult_22/SUMB[12][35] ) );
  FA_X1 \mult_22/S2_12_34  ( .A(\mult_22/ab[12][34] ), .B(
        \mult_22/CARRYB[11][34] ), .CI(\mult_22/SUMB[11][35] ), .CO(
        \mult_22/CARRYB[12][34] ), .S(\mult_22/SUMB[12][34] ) );
  FA_X1 \mult_22/S2_12_33  ( .A(\mult_22/ab[12][33] ), .B(
        \mult_22/CARRYB[11][33] ), .CI(\mult_22/SUMB[11][34] ), .CO(
        \mult_22/CARRYB[12][33] ), .S(\mult_22/SUMB[12][33] ) );
  FA_X1 \mult_22/S2_12_32  ( .A(\mult_22/ab[12][32] ), .B(
        \mult_22/CARRYB[11][32] ), .CI(\mult_22/SUMB[11][33] ), .CO(
        \mult_22/CARRYB[12][32] ), .S(\mult_22/SUMB[12][32] ) );
  FA_X1 \mult_22/S2_12_31  ( .A(\mult_22/ab[12][31] ), .B(
        \mult_22/CARRYB[11][31] ), .CI(\mult_22/SUMB[11][32] ), .CO(
        \mult_22/CARRYB[12][31] ), .S(\mult_22/SUMB[12][31] ) );
  FA_X1 \mult_22/S2_12_30  ( .A(\mult_22/ab[12][30] ), .B(
        \mult_22/CARRYB[11][30] ), .CI(\mult_22/SUMB[11][31] ), .CO(
        \mult_22/CARRYB[12][30] ), .S(\mult_22/SUMB[12][30] ) );
  FA_X1 \mult_22/S2_12_29  ( .A(\mult_22/ab[12][29] ), .B(
        \mult_22/CARRYB[11][29] ), .CI(\mult_22/SUMB[11][30] ), .CO(
        \mult_22/CARRYB[12][29] ), .S(\mult_22/SUMB[12][29] ) );
  FA_X1 \mult_22/S2_12_28  ( .A(\mult_22/ab[12][28] ), .B(
        \mult_22/CARRYB[11][28] ), .CI(\mult_22/SUMB[11][29] ), .CO(
        \mult_22/CARRYB[12][28] ), .S(\mult_22/SUMB[12][28] ) );
  FA_X1 \mult_22/S2_12_27  ( .A(\mult_22/ab[12][27] ), .B(
        \mult_22/CARRYB[11][27] ), .CI(\mult_22/SUMB[11][28] ), .CO(
        \mult_22/CARRYB[12][27] ), .S(\mult_22/SUMB[12][27] ) );
  FA_X1 \mult_22/S2_12_26  ( .A(\mult_22/ab[12][26] ), .B(
        \mult_22/CARRYB[11][26] ), .CI(\mult_22/SUMB[11][27] ), .CO(
        \mult_22/CARRYB[12][26] ), .S(\mult_22/SUMB[12][26] ) );
  FA_X1 \mult_22/S2_12_25  ( .A(\mult_22/ab[12][25] ), .B(
        \mult_22/CARRYB[11][25] ), .CI(\mult_22/SUMB[11][26] ), .CO(
        \mult_22/CARRYB[12][25] ), .S(\mult_22/SUMB[12][25] ) );
  FA_X1 \mult_22/S2_12_24  ( .A(\mult_22/ab[12][24] ), .B(
        \mult_22/CARRYB[11][24] ), .CI(\mult_22/SUMB[11][25] ), .CO(
        \mult_22/CARRYB[12][24] ), .S(\mult_22/SUMB[12][24] ) );
  FA_X1 \mult_22/S2_12_23  ( .A(\mult_22/ab[12][23] ), .B(
        \mult_22/CARRYB[11][23] ), .CI(\mult_22/SUMB[11][24] ), .CO(
        \mult_22/CARRYB[12][23] ), .S(\mult_22/SUMB[12][23] ) );
  FA_X1 \mult_22/S2_12_22  ( .A(\mult_22/ab[12][22] ), .B(
        \mult_22/CARRYB[11][22] ), .CI(\mult_22/SUMB[11][23] ), .CO(
        \mult_22/CARRYB[12][22] ), .S(\mult_22/SUMB[12][22] ) );
  FA_X1 \mult_22/S2_12_21  ( .A(\mult_22/ab[12][21] ), .B(
        \mult_22/CARRYB[11][21] ), .CI(\mult_22/SUMB[11][22] ), .CO(
        \mult_22/CARRYB[12][21] ), .S(\mult_22/SUMB[12][21] ) );
  FA_X1 \mult_22/S2_12_20  ( .A(\mult_22/ab[12][20] ), .B(
        \mult_22/CARRYB[11][20] ), .CI(\mult_22/SUMB[11][21] ), .CO(
        \mult_22/CARRYB[12][20] ), .S(\mult_22/SUMB[12][20] ) );
  FA_X1 \mult_22/S2_12_19  ( .A(\mult_22/ab[12][19] ), .B(
        \mult_22/CARRYB[11][19] ), .CI(\mult_22/SUMB[11][20] ), .CO(
        \mult_22/CARRYB[12][19] ), .S(\mult_22/SUMB[12][19] ) );
  FA_X1 \mult_22/S2_12_18  ( .A(\mult_22/ab[12][18] ), .B(
        \mult_22/CARRYB[11][18] ), .CI(\mult_22/SUMB[11][19] ), .CO(
        \mult_22/CARRYB[12][18] ), .S(\mult_22/SUMB[12][18] ) );
  FA_X1 \mult_22/S2_12_17  ( .A(\mult_22/ab[12][17] ), .B(
        \mult_22/CARRYB[11][17] ), .CI(\mult_22/SUMB[11][18] ), .CO(
        \mult_22/CARRYB[12][17] ), .S(\mult_22/SUMB[12][17] ) );
  FA_X1 \mult_22/S2_12_16  ( .A(\mult_22/ab[12][16] ), .B(
        \mult_22/CARRYB[11][16] ), .CI(\mult_22/SUMB[11][17] ), .CO(
        \mult_22/CARRYB[12][16] ), .S(\mult_22/SUMB[12][16] ) );
  FA_X1 \mult_22/S2_12_15  ( .A(\mult_22/ab[12][15] ), .B(
        \mult_22/CARRYB[11][15] ), .CI(\mult_22/SUMB[11][16] ), .CO(
        \mult_22/CARRYB[12][15] ), .S(\mult_22/SUMB[12][15] ) );
  FA_X1 \mult_22/S2_12_14  ( .A(\mult_22/ab[12][14] ), .B(
        \mult_22/CARRYB[11][14] ), .CI(\mult_22/SUMB[11][15] ), .CO(
        \mult_22/CARRYB[12][14] ), .S(\mult_22/SUMB[12][14] ) );
  FA_X1 \mult_22/S2_12_13  ( .A(\mult_22/ab[12][13] ), .B(
        \mult_22/CARRYB[11][13] ), .CI(\mult_22/SUMB[11][14] ), .CO(
        \mult_22/CARRYB[12][13] ), .S(\mult_22/SUMB[12][13] ) );
  FA_X1 \mult_22/S2_12_12  ( .A(\mult_22/ab[12][12] ), .B(
        \mult_22/CARRYB[11][12] ), .CI(\mult_22/SUMB[11][13] ), .CO(
        \mult_22/CARRYB[12][12] ), .S(\mult_22/SUMB[12][12] ) );
  FA_X1 \mult_22/S2_12_11  ( .A(\mult_22/ab[12][11] ), .B(
        \mult_22/CARRYB[11][11] ), .CI(\mult_22/SUMB[11][12] ), .CO(
        \mult_22/CARRYB[12][11] ), .S(\mult_22/SUMB[12][11] ) );
  FA_X1 \mult_22/S2_12_10  ( .A(\mult_22/ab[12][10] ), .B(
        \mult_22/CARRYB[11][10] ), .CI(\mult_22/SUMB[11][11] ), .CO(
        \mult_22/CARRYB[12][10] ), .S(\mult_22/SUMB[12][10] ) );
  FA_X1 \mult_22/S2_12_9  ( .A(\mult_22/ab[12][9] ), .B(
        \mult_22/CARRYB[11][9] ), .CI(\mult_22/SUMB[11][10] ), .CO(
        \mult_22/CARRYB[12][9] ), .S(\mult_22/SUMB[12][9] ) );
  FA_X1 \mult_22/S2_12_8  ( .A(\mult_22/ab[12][8] ), .B(
        \mult_22/CARRYB[11][8] ), .CI(\mult_22/SUMB[11][9] ), .CO(
        \mult_22/CARRYB[12][8] ), .S(\mult_22/SUMB[12][8] ) );
  FA_X1 \mult_22/S2_12_7  ( .A(\mult_22/ab[12][7] ), .B(
        \mult_22/CARRYB[11][7] ), .CI(\mult_22/SUMB[11][8] ), .CO(
        \mult_22/CARRYB[12][7] ), .S(\mult_22/SUMB[12][7] ) );
  FA_X1 \mult_22/S2_12_6  ( .A(\mult_22/ab[12][6] ), .B(
        \mult_22/CARRYB[11][6] ), .CI(\mult_22/SUMB[11][7] ), .CO(
        \mult_22/CARRYB[12][6] ), .S(\mult_22/SUMB[12][6] ) );
  FA_X1 \mult_22/S2_12_5  ( .A(\mult_22/ab[12][5] ), .B(
        \mult_22/CARRYB[11][5] ), .CI(\mult_22/SUMB[11][6] ), .CO(
        \mult_22/CARRYB[12][5] ), .S(\mult_22/SUMB[12][5] ) );
  FA_X1 \mult_22/S2_12_4  ( .A(\mult_22/ab[12][4] ), .B(
        \mult_22/CARRYB[11][4] ), .CI(\mult_22/SUMB[11][5] ), .CO(
        \mult_22/CARRYB[12][4] ), .S(\mult_22/SUMB[12][4] ) );
  FA_X1 \mult_22/S2_12_3  ( .A(\mult_22/ab[12][3] ), .B(
        \mult_22/CARRYB[11][3] ), .CI(\mult_22/SUMB[11][4] ), .CO(
        \mult_22/CARRYB[12][3] ), .S(\mult_22/SUMB[12][3] ) );
  FA_X1 \mult_22/S2_12_2  ( .A(\mult_22/ab[12][2] ), .B(
        \mult_22/CARRYB[11][2] ), .CI(\mult_22/SUMB[11][3] ), .CO(
        \mult_22/CARRYB[12][2] ), .S(\mult_22/SUMB[12][2] ) );
  FA_X1 \mult_22/S2_12_1  ( .A(\mult_22/ab[12][1] ), .B(
        \mult_22/CARRYB[11][1] ), .CI(\mult_22/SUMB[11][2] ), .CO(
        \mult_22/CARRYB[12][1] ), .S(\mult_22/SUMB[12][1] ) );
  FA_X1 \mult_22/S1_12_0  ( .A(\mult_22/ab[12][0] ), .B(
        \mult_22/CARRYB[11][0] ), .CI(\mult_22/SUMB[11][1] ), .CO(
        \mult_22/CARRYB[12][0] ), .S(N140) );
  FA_X1 \mult_22/S3_13_62  ( .A(\mult_22/ab[13][62] ), .B(
        \mult_22/CARRYB[12][62] ), .CI(\mult_22/ab[12][63] ), .CO(
        \mult_22/CARRYB[13][62] ), .S(\mult_22/SUMB[13][62] ) );
  FA_X1 \mult_22/S2_13_61  ( .A(\mult_22/ab[13][61] ), .B(
        \mult_22/CARRYB[12][61] ), .CI(\mult_22/SUMB[12][62] ), .CO(
        \mult_22/CARRYB[13][61] ), .S(\mult_22/SUMB[13][61] ) );
  FA_X1 \mult_22/S2_13_60  ( .A(\mult_22/ab[13][60] ), .B(
        \mult_22/CARRYB[12][60] ), .CI(\mult_22/SUMB[12][61] ), .CO(
        \mult_22/CARRYB[13][60] ), .S(\mult_22/SUMB[13][60] ) );
  FA_X1 \mult_22/S2_13_59  ( .A(\mult_22/ab[13][59] ), .B(
        \mult_22/CARRYB[12][59] ), .CI(\mult_22/SUMB[12][60] ), .CO(
        \mult_22/CARRYB[13][59] ), .S(\mult_22/SUMB[13][59] ) );
  FA_X1 \mult_22/S2_13_58  ( .A(\mult_22/ab[13][58] ), .B(
        \mult_22/CARRYB[12][58] ), .CI(\mult_22/SUMB[12][59] ), .CO(
        \mult_22/CARRYB[13][58] ), .S(\mult_22/SUMB[13][58] ) );
  FA_X1 \mult_22/S2_13_57  ( .A(\mult_22/ab[13][57] ), .B(
        \mult_22/CARRYB[12][57] ), .CI(\mult_22/SUMB[12][58] ), .CO(
        \mult_22/CARRYB[13][57] ), .S(\mult_22/SUMB[13][57] ) );
  FA_X1 \mult_22/S2_13_56  ( .A(\mult_22/ab[13][56] ), .B(
        \mult_22/CARRYB[12][56] ), .CI(\mult_22/SUMB[12][57] ), .CO(
        \mult_22/CARRYB[13][56] ), .S(\mult_22/SUMB[13][56] ) );
  FA_X1 \mult_22/S2_13_55  ( .A(\mult_22/ab[13][55] ), .B(
        \mult_22/CARRYB[12][55] ), .CI(\mult_22/SUMB[12][56] ), .CO(
        \mult_22/CARRYB[13][55] ), .S(\mult_22/SUMB[13][55] ) );
  FA_X1 \mult_22/S2_13_54  ( .A(\mult_22/CARRYB[12][54] ), .B(
        \mult_22/ab[13][54] ), .CI(\mult_22/SUMB[12][55] ), .CO(
        \mult_22/CARRYB[13][54] ), .S(\mult_22/SUMB[13][54] ) );
  FA_X1 \mult_22/S2_13_53  ( .A(\mult_22/ab[13][53] ), .B(
        \mult_22/CARRYB[12][53] ), .CI(\mult_22/SUMB[12][54] ), .CO(
        \mult_22/CARRYB[13][53] ), .S(\mult_22/SUMB[13][53] ) );
  FA_X1 \mult_22/S2_13_52  ( .A(\mult_22/CARRYB[12][52] ), .B(
        \mult_22/ab[13][52] ), .CI(\mult_22/SUMB[12][53] ), .CO(
        \mult_22/CARRYB[13][52] ), .S(\mult_22/SUMB[13][52] ) );
  FA_X1 \mult_22/S2_13_51  ( .A(\mult_22/CARRYB[12][51] ), .B(
        \mult_22/ab[13][51] ), .CI(\mult_22/SUMB[12][52] ), .CO(
        \mult_22/CARRYB[13][51] ), .S(\mult_22/SUMB[13][51] ) );
  FA_X1 \mult_22/S2_13_50  ( .A(\mult_22/ab[13][50] ), .B(
        \mult_22/CARRYB[12][50] ), .CI(\mult_22/SUMB[12][51] ), .CO(
        \mult_22/CARRYB[13][50] ), .S(\mult_22/SUMB[13][50] ) );
  FA_X1 \mult_22/S2_13_49  ( .A(\mult_22/ab[13][49] ), .B(
        \mult_22/CARRYB[12][49] ), .CI(\mult_22/SUMB[12][50] ), .CO(
        \mult_22/CARRYB[13][49] ), .S(\mult_22/SUMB[13][49] ) );
  FA_X1 \mult_22/S2_13_48  ( .A(\mult_22/ab[13][48] ), .B(
        \mult_22/CARRYB[12][48] ), .CI(\mult_22/SUMB[12][49] ), .CO(
        \mult_22/CARRYB[13][48] ), .S(\mult_22/SUMB[13][48] ) );
  FA_X1 \mult_22/S2_13_47  ( .A(\mult_22/ab[13][47] ), .B(
        \mult_22/CARRYB[12][47] ), .CI(\mult_22/SUMB[12][48] ), .CO(
        \mult_22/CARRYB[13][47] ), .S(\mult_22/SUMB[13][47] ) );
  FA_X1 \mult_22/S2_13_46  ( .A(\mult_22/ab[13][46] ), .B(
        \mult_22/CARRYB[12][46] ), .CI(\mult_22/SUMB[12][47] ), .CO(
        \mult_22/CARRYB[13][46] ), .S(\mult_22/SUMB[13][46] ) );
  FA_X1 \mult_22/S2_13_45  ( .A(\mult_22/ab[13][45] ), .B(
        \mult_22/CARRYB[12][45] ), .CI(\mult_22/SUMB[12][46] ), .CO(
        \mult_22/CARRYB[13][45] ), .S(\mult_22/SUMB[13][45] ) );
  FA_X1 \mult_22/S2_13_44  ( .A(\mult_22/ab[13][44] ), .B(
        \mult_22/CARRYB[12][44] ), .CI(\mult_22/SUMB[12][45] ), .CO(
        \mult_22/CARRYB[13][44] ), .S(\mult_22/SUMB[13][44] ) );
  FA_X1 \mult_22/S2_13_43  ( .A(\mult_22/ab[13][43] ), .B(
        \mult_22/CARRYB[12][43] ), .CI(\mult_22/SUMB[12][44] ), .CO(
        \mult_22/CARRYB[13][43] ), .S(\mult_22/SUMB[13][43] ) );
  FA_X1 \mult_22/S2_13_42  ( .A(\mult_22/ab[13][42] ), .B(
        \mult_22/CARRYB[12][42] ), .CI(\mult_22/SUMB[12][43] ), .CO(
        \mult_22/CARRYB[13][42] ), .S(\mult_22/SUMB[13][42] ) );
  FA_X1 \mult_22/S2_13_41  ( .A(\mult_22/ab[13][41] ), .B(
        \mult_22/CARRYB[12][41] ), .CI(\mult_22/SUMB[12][42] ), .CO(
        \mult_22/CARRYB[13][41] ), .S(\mult_22/SUMB[13][41] ) );
  FA_X1 \mult_22/S2_13_40  ( .A(\mult_22/ab[13][40] ), .B(
        \mult_22/CARRYB[12][40] ), .CI(\mult_22/SUMB[12][41] ), .CO(
        \mult_22/CARRYB[13][40] ), .S(\mult_22/SUMB[13][40] ) );
  FA_X1 \mult_22/S2_13_39  ( .A(\mult_22/ab[13][39] ), .B(
        \mult_22/CARRYB[12][39] ), .CI(\mult_22/SUMB[12][40] ), .CO(
        \mult_22/CARRYB[13][39] ), .S(\mult_22/SUMB[13][39] ) );
  FA_X1 \mult_22/S2_13_38  ( .A(\mult_22/ab[13][38] ), .B(
        \mult_22/CARRYB[12][38] ), .CI(\mult_22/SUMB[12][39] ), .CO(
        \mult_22/CARRYB[13][38] ), .S(\mult_22/SUMB[13][38] ) );
  FA_X1 \mult_22/S2_13_37  ( .A(\mult_22/ab[13][37] ), .B(
        \mult_22/CARRYB[12][37] ), .CI(\mult_22/SUMB[12][38] ), .CO(
        \mult_22/CARRYB[13][37] ), .S(\mult_22/SUMB[13][37] ) );
  FA_X1 \mult_22/S2_13_36  ( .A(\mult_22/ab[13][36] ), .B(
        \mult_22/CARRYB[12][36] ), .CI(\mult_22/SUMB[12][37] ), .CO(
        \mult_22/CARRYB[13][36] ), .S(\mult_22/SUMB[13][36] ) );
  FA_X1 \mult_22/S2_13_35  ( .A(\mult_22/ab[13][35] ), .B(
        \mult_22/CARRYB[12][35] ), .CI(\mult_22/SUMB[12][36] ), .CO(
        \mult_22/CARRYB[13][35] ), .S(\mult_22/SUMB[13][35] ) );
  FA_X1 \mult_22/S2_13_34  ( .A(\mult_22/ab[13][34] ), .B(
        \mult_22/CARRYB[12][34] ), .CI(\mult_22/SUMB[12][35] ), .CO(
        \mult_22/CARRYB[13][34] ), .S(\mult_22/SUMB[13][34] ) );
  FA_X1 \mult_22/S2_13_33  ( .A(\mult_22/ab[13][33] ), .B(
        \mult_22/CARRYB[12][33] ), .CI(\mult_22/SUMB[12][34] ), .CO(
        \mult_22/CARRYB[13][33] ), .S(\mult_22/SUMB[13][33] ) );
  FA_X1 \mult_22/S2_13_32  ( .A(\mult_22/ab[13][32] ), .B(
        \mult_22/CARRYB[12][32] ), .CI(\mult_22/SUMB[12][33] ), .CO(
        \mult_22/CARRYB[13][32] ), .S(\mult_22/SUMB[13][32] ) );
  FA_X1 \mult_22/S2_13_31  ( .A(\mult_22/ab[13][31] ), .B(
        \mult_22/CARRYB[12][31] ), .CI(\mult_22/SUMB[12][32] ), .CO(
        \mult_22/CARRYB[13][31] ), .S(\mult_22/SUMB[13][31] ) );
  FA_X1 \mult_22/S2_13_30  ( .A(\mult_22/ab[13][30] ), .B(
        \mult_22/CARRYB[12][30] ), .CI(\mult_22/SUMB[12][31] ), .CO(
        \mult_22/CARRYB[13][30] ), .S(\mult_22/SUMB[13][30] ) );
  FA_X1 \mult_22/S2_13_29  ( .A(\mult_22/ab[13][29] ), .B(
        \mult_22/CARRYB[12][29] ), .CI(\mult_22/SUMB[12][30] ), .CO(
        \mult_22/CARRYB[13][29] ), .S(\mult_22/SUMB[13][29] ) );
  FA_X1 \mult_22/S2_13_28  ( .A(\mult_22/ab[13][28] ), .B(
        \mult_22/CARRYB[12][28] ), .CI(\mult_22/SUMB[12][29] ), .CO(
        \mult_22/CARRYB[13][28] ), .S(\mult_22/SUMB[13][28] ) );
  FA_X1 \mult_22/S2_13_27  ( .A(\mult_22/ab[13][27] ), .B(
        \mult_22/CARRYB[12][27] ), .CI(\mult_22/SUMB[12][28] ), .CO(
        \mult_22/CARRYB[13][27] ), .S(\mult_22/SUMB[13][27] ) );
  FA_X1 \mult_22/S2_13_26  ( .A(\mult_22/ab[13][26] ), .B(
        \mult_22/CARRYB[12][26] ), .CI(\mult_22/SUMB[12][27] ), .CO(
        \mult_22/CARRYB[13][26] ), .S(\mult_22/SUMB[13][26] ) );
  FA_X1 \mult_22/S2_13_25  ( .A(\mult_22/ab[13][25] ), .B(
        \mult_22/CARRYB[12][25] ), .CI(\mult_22/SUMB[12][26] ), .CO(
        \mult_22/CARRYB[13][25] ), .S(\mult_22/SUMB[13][25] ) );
  FA_X1 \mult_22/S2_13_24  ( .A(\mult_22/ab[13][24] ), .B(
        \mult_22/CARRYB[12][24] ), .CI(\mult_22/SUMB[12][25] ), .CO(
        \mult_22/CARRYB[13][24] ), .S(\mult_22/SUMB[13][24] ) );
  FA_X1 \mult_22/S2_13_23  ( .A(\mult_22/ab[13][23] ), .B(
        \mult_22/CARRYB[12][23] ), .CI(\mult_22/SUMB[12][24] ), .CO(
        \mult_22/CARRYB[13][23] ), .S(\mult_22/SUMB[13][23] ) );
  FA_X1 \mult_22/S2_13_22  ( .A(\mult_22/ab[13][22] ), .B(
        \mult_22/CARRYB[12][22] ), .CI(\mult_22/SUMB[12][23] ), .CO(
        \mult_22/CARRYB[13][22] ), .S(\mult_22/SUMB[13][22] ) );
  FA_X1 \mult_22/S2_13_21  ( .A(\mult_22/ab[13][21] ), .B(
        \mult_22/CARRYB[12][21] ), .CI(\mult_22/SUMB[12][22] ), .CO(
        \mult_22/CARRYB[13][21] ), .S(\mult_22/SUMB[13][21] ) );
  FA_X1 \mult_22/S2_13_20  ( .A(\mult_22/ab[13][20] ), .B(
        \mult_22/CARRYB[12][20] ), .CI(\mult_22/SUMB[12][21] ), .CO(
        \mult_22/CARRYB[13][20] ), .S(\mult_22/SUMB[13][20] ) );
  FA_X1 \mult_22/S2_13_19  ( .A(\mult_22/ab[13][19] ), .B(
        \mult_22/CARRYB[12][19] ), .CI(\mult_22/SUMB[12][20] ), .CO(
        \mult_22/CARRYB[13][19] ), .S(\mult_22/SUMB[13][19] ) );
  FA_X1 \mult_22/S2_13_18  ( .A(\mult_22/ab[13][18] ), .B(
        \mult_22/CARRYB[12][18] ), .CI(\mult_22/SUMB[12][19] ), .CO(
        \mult_22/CARRYB[13][18] ), .S(\mult_22/SUMB[13][18] ) );
  FA_X1 \mult_22/S2_13_17  ( .A(\mult_22/ab[13][17] ), .B(
        \mult_22/CARRYB[12][17] ), .CI(\mult_22/SUMB[12][18] ), .CO(
        \mult_22/CARRYB[13][17] ), .S(\mult_22/SUMB[13][17] ) );
  FA_X1 \mult_22/S2_13_16  ( .A(\mult_22/ab[13][16] ), .B(
        \mult_22/CARRYB[12][16] ), .CI(\mult_22/SUMB[12][17] ), .CO(
        \mult_22/CARRYB[13][16] ), .S(\mult_22/SUMB[13][16] ) );
  FA_X1 \mult_22/S2_13_15  ( .A(\mult_22/ab[13][15] ), .B(
        \mult_22/CARRYB[12][15] ), .CI(\mult_22/SUMB[12][16] ), .CO(
        \mult_22/CARRYB[13][15] ), .S(\mult_22/SUMB[13][15] ) );
  FA_X1 \mult_22/S2_13_14  ( .A(\mult_22/ab[13][14] ), .B(
        \mult_22/CARRYB[12][14] ), .CI(\mult_22/SUMB[12][15] ), .CO(
        \mult_22/CARRYB[13][14] ), .S(\mult_22/SUMB[13][14] ) );
  FA_X1 \mult_22/S2_13_13  ( .A(\mult_22/ab[13][13] ), .B(
        \mult_22/CARRYB[12][13] ), .CI(\mult_22/SUMB[12][14] ), .CO(
        \mult_22/CARRYB[13][13] ), .S(\mult_22/SUMB[13][13] ) );
  FA_X1 \mult_22/S2_13_12  ( .A(\mult_22/ab[13][12] ), .B(
        \mult_22/CARRYB[12][12] ), .CI(\mult_22/SUMB[12][13] ), .CO(
        \mult_22/CARRYB[13][12] ), .S(\mult_22/SUMB[13][12] ) );
  FA_X1 \mult_22/S2_13_11  ( .A(\mult_22/ab[13][11] ), .B(
        \mult_22/CARRYB[12][11] ), .CI(\mult_22/SUMB[12][12] ), .CO(
        \mult_22/CARRYB[13][11] ), .S(\mult_22/SUMB[13][11] ) );
  FA_X1 \mult_22/S2_13_10  ( .A(\mult_22/ab[13][10] ), .B(
        \mult_22/CARRYB[12][10] ), .CI(\mult_22/SUMB[12][11] ), .CO(
        \mult_22/CARRYB[13][10] ), .S(\mult_22/SUMB[13][10] ) );
  FA_X1 \mult_22/S2_13_9  ( .A(\mult_22/ab[13][9] ), .B(
        \mult_22/CARRYB[12][9] ), .CI(\mult_22/SUMB[12][10] ), .CO(
        \mult_22/CARRYB[13][9] ), .S(\mult_22/SUMB[13][9] ) );
  FA_X1 \mult_22/S2_13_8  ( .A(\mult_22/ab[13][8] ), .B(
        \mult_22/CARRYB[12][8] ), .CI(\mult_22/SUMB[12][9] ), .CO(
        \mult_22/CARRYB[13][8] ), .S(\mult_22/SUMB[13][8] ) );
  FA_X1 \mult_22/S2_13_7  ( .A(\mult_22/ab[13][7] ), .B(
        \mult_22/CARRYB[12][7] ), .CI(\mult_22/SUMB[12][8] ), .CO(
        \mult_22/CARRYB[13][7] ), .S(\mult_22/SUMB[13][7] ) );
  FA_X1 \mult_22/S2_13_6  ( .A(\mult_22/ab[13][6] ), .B(
        \mult_22/CARRYB[12][6] ), .CI(\mult_22/SUMB[12][7] ), .CO(
        \mult_22/CARRYB[13][6] ), .S(\mult_22/SUMB[13][6] ) );
  FA_X1 \mult_22/S2_13_5  ( .A(\mult_22/ab[13][5] ), .B(
        \mult_22/CARRYB[12][5] ), .CI(\mult_22/SUMB[12][6] ), .CO(
        \mult_22/CARRYB[13][5] ), .S(\mult_22/SUMB[13][5] ) );
  FA_X1 \mult_22/S2_13_4  ( .A(\mult_22/ab[13][4] ), .B(
        \mult_22/CARRYB[12][4] ), .CI(\mult_22/SUMB[12][5] ), .CO(
        \mult_22/CARRYB[13][4] ), .S(\mult_22/SUMB[13][4] ) );
  FA_X1 \mult_22/S2_13_3  ( .A(\mult_22/ab[13][3] ), .B(
        \mult_22/CARRYB[12][3] ), .CI(\mult_22/SUMB[12][4] ), .CO(
        \mult_22/CARRYB[13][3] ), .S(\mult_22/SUMB[13][3] ) );
  FA_X1 \mult_22/S2_13_2  ( .A(\mult_22/ab[13][2] ), .B(
        \mult_22/CARRYB[12][2] ), .CI(\mult_22/SUMB[12][3] ), .CO(
        \mult_22/CARRYB[13][2] ), .S(\mult_22/SUMB[13][2] ) );
  FA_X1 \mult_22/S2_13_1  ( .A(\mult_22/ab[13][1] ), .B(
        \mult_22/CARRYB[12][1] ), .CI(\mult_22/SUMB[12][2] ), .CO(
        \mult_22/CARRYB[13][1] ), .S(\mult_22/SUMB[13][1] ) );
  FA_X1 \mult_22/S1_13_0  ( .A(\mult_22/ab[13][0] ), .B(
        \mult_22/CARRYB[12][0] ), .CI(\mult_22/SUMB[12][1] ), .CO(
        \mult_22/CARRYB[13][0] ), .S(N141) );
  FA_X1 \mult_22/S3_14_62  ( .A(\mult_22/ab[14][62] ), .B(
        \mult_22/CARRYB[13][62] ), .CI(\mult_22/ab[13][63] ), .CO(
        \mult_22/CARRYB[14][62] ), .S(\mult_22/SUMB[14][62] ) );
  FA_X1 \mult_22/S2_14_61  ( .A(\mult_22/ab[14][61] ), .B(
        \mult_22/CARRYB[13][61] ), .CI(\mult_22/SUMB[13][62] ), .CO(
        \mult_22/CARRYB[14][61] ), .S(\mult_22/SUMB[14][61] ) );
  FA_X1 \mult_22/S2_14_60  ( .A(\mult_22/ab[14][60] ), .B(
        \mult_22/CARRYB[13][60] ), .CI(\mult_22/SUMB[13][61] ), .CO(
        \mult_22/CARRYB[14][60] ), .S(\mult_22/SUMB[14][60] ) );
  FA_X1 \mult_22/S2_14_59  ( .A(\mult_22/ab[14][59] ), .B(
        \mult_22/CARRYB[13][59] ), .CI(\mult_22/SUMB[13][60] ), .CO(
        \mult_22/CARRYB[14][59] ), .S(\mult_22/SUMB[14][59] ) );
  FA_X1 \mult_22/S2_14_58  ( .A(\mult_22/ab[14][58] ), .B(
        \mult_22/CARRYB[13][58] ), .CI(\mult_22/SUMB[13][59] ), .CO(
        \mult_22/CARRYB[14][58] ), .S(\mult_22/SUMB[14][58] ) );
  FA_X1 \mult_22/S2_14_57  ( .A(\mult_22/ab[14][57] ), .B(
        \mult_22/CARRYB[13][57] ), .CI(\mult_22/SUMB[13][58] ), .CO(
        \mult_22/CARRYB[14][57] ), .S(\mult_22/SUMB[14][57] ) );
  FA_X1 \mult_22/S2_14_56  ( .A(\mult_22/ab[14][56] ), .B(
        \mult_22/CARRYB[13][56] ), .CI(\mult_22/SUMB[13][57] ), .CO(
        \mult_22/CARRYB[14][56] ), .S(\mult_22/SUMB[14][56] ) );
  FA_X1 \mult_22/S2_14_55  ( .A(\mult_22/ab[14][55] ), .B(
        \mult_22/CARRYB[13][55] ), .CI(\mult_22/SUMB[13][56] ), .CO(
        \mult_22/CARRYB[14][55] ), .S(\mult_22/SUMB[14][55] ) );
  FA_X1 \mult_22/S2_14_54  ( .A(\mult_22/ab[14][54] ), .B(
        \mult_22/CARRYB[13][54] ), .CI(\mult_22/SUMB[13][55] ), .CO(
        \mult_22/CARRYB[14][54] ), .S(\mult_22/SUMB[14][54] ) );
  FA_X1 \mult_22/S2_14_53  ( .A(\mult_22/ab[14][53] ), .B(
        \mult_22/CARRYB[13][53] ), .CI(\mult_22/SUMB[13][54] ), .CO(
        \mult_22/CARRYB[14][53] ), .S(\mult_22/SUMB[14][53] ) );
  FA_X1 \mult_22/S2_14_52  ( .A(\mult_22/CARRYB[13][52] ), .B(
        \mult_22/ab[14][52] ), .CI(\mult_22/SUMB[13][53] ), .CO(
        \mult_22/CARRYB[14][52] ), .S(\mult_22/SUMB[14][52] ) );
  FA_X1 \mult_22/S2_14_51  ( .A(\mult_22/ab[14][51] ), .B(
        \mult_22/CARRYB[13][51] ), .CI(\mult_22/SUMB[13][52] ), .CO(
        \mult_22/CARRYB[14][51] ), .S(\mult_22/SUMB[14][51] ) );
  FA_X1 \mult_22/S2_14_50  ( .A(\mult_22/CARRYB[13][50] ), .B(
        \mult_22/ab[14][50] ), .CI(\mult_22/SUMB[13][51] ), .CO(
        \mult_22/CARRYB[14][50] ), .S(\mult_22/SUMB[14][50] ) );
  FA_X1 \mult_22/S2_14_49  ( .A(\mult_22/ab[14][49] ), .B(
        \mult_22/CARRYB[13][49] ), .CI(\mult_22/SUMB[13][50] ), .CO(
        \mult_22/CARRYB[14][49] ), .S(\mult_22/SUMB[14][49] ) );
  FA_X1 \mult_22/S2_14_48  ( .A(\mult_22/ab[14][48] ), .B(
        \mult_22/CARRYB[13][48] ), .CI(\mult_22/SUMB[13][49] ), .CO(
        \mult_22/CARRYB[14][48] ), .S(\mult_22/SUMB[14][48] ) );
  FA_X1 \mult_22/S2_14_46  ( .A(\mult_22/ab[14][46] ), .B(
        \mult_22/CARRYB[13][46] ), .CI(\mult_22/SUMB[13][47] ), .CO(
        \mult_22/CARRYB[14][46] ), .S(\mult_22/SUMB[14][46] ) );
  FA_X1 \mult_22/S2_14_45  ( .A(\mult_22/ab[14][45] ), .B(
        \mult_22/CARRYB[13][45] ), .CI(\mult_22/SUMB[13][46] ), .CO(
        \mult_22/CARRYB[14][45] ), .S(\mult_22/SUMB[14][45] ) );
  FA_X1 \mult_22/S2_14_44  ( .A(\mult_22/ab[14][44] ), .B(
        \mult_22/CARRYB[13][44] ), .CI(\mult_22/SUMB[13][45] ), .CO(
        \mult_22/CARRYB[14][44] ), .S(\mult_22/SUMB[14][44] ) );
  FA_X1 \mult_22/S2_14_43  ( .A(\mult_22/ab[14][43] ), .B(
        \mult_22/CARRYB[13][43] ), .CI(\mult_22/SUMB[13][44] ), .CO(
        \mult_22/CARRYB[14][43] ), .S(\mult_22/SUMB[14][43] ) );
  FA_X1 \mult_22/S2_14_42  ( .A(\mult_22/ab[14][42] ), .B(
        \mult_22/CARRYB[13][42] ), .CI(\mult_22/SUMB[13][43] ), .CO(
        \mult_22/CARRYB[14][42] ), .S(\mult_22/SUMB[14][42] ) );
  FA_X1 \mult_22/S2_14_41  ( .A(\mult_22/ab[14][41] ), .B(
        \mult_22/CARRYB[13][41] ), .CI(\mult_22/SUMB[13][42] ), .CO(
        \mult_22/CARRYB[14][41] ), .S(\mult_22/SUMB[14][41] ) );
  FA_X1 \mult_22/S2_14_40  ( .A(\mult_22/ab[14][40] ), .B(
        \mult_22/CARRYB[13][40] ), .CI(\mult_22/SUMB[13][41] ), .CO(
        \mult_22/CARRYB[14][40] ), .S(\mult_22/SUMB[14][40] ) );
  FA_X1 \mult_22/S2_14_39  ( .A(\mult_22/ab[14][39] ), .B(
        \mult_22/CARRYB[13][39] ), .CI(\mult_22/SUMB[13][40] ), .CO(
        \mult_22/CARRYB[14][39] ), .S(\mult_22/SUMB[14][39] ) );
  FA_X1 \mult_22/S2_14_38  ( .A(\mult_22/ab[14][38] ), .B(
        \mult_22/CARRYB[13][38] ), .CI(\mult_22/SUMB[13][39] ), .CO(
        \mult_22/CARRYB[14][38] ), .S(\mult_22/SUMB[14][38] ) );
  FA_X1 \mult_22/S2_14_37  ( .A(\mult_22/ab[14][37] ), .B(
        \mult_22/CARRYB[13][37] ), .CI(\mult_22/SUMB[13][38] ), .CO(
        \mult_22/CARRYB[14][37] ), .S(\mult_22/SUMB[14][37] ) );
  FA_X1 \mult_22/S2_14_36  ( .A(\mult_22/ab[14][36] ), .B(
        \mult_22/CARRYB[13][36] ), .CI(\mult_22/SUMB[13][37] ), .CO(
        \mult_22/CARRYB[14][36] ), .S(\mult_22/SUMB[14][36] ) );
  FA_X1 \mult_22/S2_14_35  ( .A(\mult_22/ab[14][35] ), .B(
        \mult_22/CARRYB[13][35] ), .CI(\mult_22/SUMB[13][36] ), .CO(
        \mult_22/CARRYB[14][35] ), .S(\mult_22/SUMB[14][35] ) );
  FA_X1 \mult_22/S2_14_34  ( .A(\mult_22/ab[14][34] ), .B(
        \mult_22/CARRYB[13][34] ), .CI(\mult_22/SUMB[13][35] ), .CO(
        \mult_22/CARRYB[14][34] ), .S(\mult_22/SUMB[14][34] ) );
  FA_X1 \mult_22/S2_14_33  ( .A(\mult_22/ab[14][33] ), .B(
        \mult_22/CARRYB[13][33] ), .CI(\mult_22/SUMB[13][34] ), .CO(
        \mult_22/CARRYB[14][33] ), .S(\mult_22/SUMB[14][33] ) );
  FA_X1 \mult_22/S2_14_32  ( .A(\mult_22/ab[14][32] ), .B(
        \mult_22/CARRYB[13][32] ), .CI(\mult_22/SUMB[13][33] ), .CO(
        \mult_22/CARRYB[14][32] ), .S(\mult_22/SUMB[14][32] ) );
  FA_X1 \mult_22/S2_14_31  ( .A(\mult_22/ab[14][31] ), .B(
        \mult_22/CARRYB[13][31] ), .CI(\mult_22/SUMB[13][32] ), .CO(
        \mult_22/CARRYB[14][31] ), .S(\mult_22/SUMB[14][31] ) );
  FA_X1 \mult_22/S2_14_30  ( .A(\mult_22/ab[14][30] ), .B(
        \mult_22/CARRYB[13][30] ), .CI(\mult_22/SUMB[13][31] ), .CO(
        \mult_22/CARRYB[14][30] ), .S(\mult_22/SUMB[14][30] ) );
  FA_X1 \mult_22/S2_14_29  ( .A(\mult_22/ab[14][29] ), .B(
        \mult_22/CARRYB[13][29] ), .CI(\mult_22/SUMB[13][30] ), .CO(
        \mult_22/CARRYB[14][29] ), .S(\mult_22/SUMB[14][29] ) );
  FA_X1 \mult_22/S2_14_28  ( .A(\mult_22/ab[14][28] ), .B(
        \mult_22/CARRYB[13][28] ), .CI(\mult_22/SUMB[13][29] ), .CO(
        \mult_22/CARRYB[14][28] ), .S(\mult_22/SUMB[14][28] ) );
  FA_X1 \mult_22/S2_14_27  ( .A(\mult_22/ab[14][27] ), .B(
        \mult_22/CARRYB[13][27] ), .CI(\mult_22/SUMB[13][28] ), .CO(
        \mult_22/CARRYB[14][27] ), .S(\mult_22/SUMB[14][27] ) );
  FA_X1 \mult_22/S2_14_26  ( .A(\mult_22/ab[14][26] ), .B(
        \mult_22/CARRYB[13][26] ), .CI(\mult_22/SUMB[13][27] ), .CO(
        \mult_22/CARRYB[14][26] ), .S(\mult_22/SUMB[14][26] ) );
  FA_X1 \mult_22/S2_14_25  ( .A(\mult_22/ab[14][25] ), .B(
        \mult_22/CARRYB[13][25] ), .CI(\mult_22/SUMB[13][26] ), .CO(
        \mult_22/CARRYB[14][25] ), .S(\mult_22/SUMB[14][25] ) );
  FA_X1 \mult_22/S2_14_24  ( .A(\mult_22/ab[14][24] ), .B(
        \mult_22/CARRYB[13][24] ), .CI(\mult_22/SUMB[13][25] ), .CO(
        \mult_22/CARRYB[14][24] ), .S(\mult_22/SUMB[14][24] ) );
  FA_X1 \mult_22/S2_14_23  ( .A(\mult_22/ab[14][23] ), .B(
        \mult_22/CARRYB[13][23] ), .CI(\mult_22/SUMB[13][24] ), .CO(
        \mult_22/CARRYB[14][23] ), .S(\mult_22/SUMB[14][23] ) );
  FA_X1 \mult_22/S2_14_22  ( .A(\mult_22/ab[14][22] ), .B(
        \mult_22/CARRYB[13][22] ), .CI(\mult_22/SUMB[13][23] ), .CO(
        \mult_22/CARRYB[14][22] ), .S(\mult_22/SUMB[14][22] ) );
  FA_X1 \mult_22/S2_14_21  ( .A(\mult_22/ab[14][21] ), .B(
        \mult_22/CARRYB[13][21] ), .CI(\mult_22/SUMB[13][22] ), .CO(
        \mult_22/CARRYB[14][21] ), .S(\mult_22/SUMB[14][21] ) );
  FA_X1 \mult_22/S2_14_20  ( .A(\mult_22/ab[14][20] ), .B(
        \mult_22/CARRYB[13][20] ), .CI(\mult_22/SUMB[13][21] ), .CO(
        \mult_22/CARRYB[14][20] ), .S(\mult_22/SUMB[14][20] ) );
  FA_X1 \mult_22/S2_14_19  ( .A(\mult_22/ab[14][19] ), .B(
        \mult_22/CARRYB[13][19] ), .CI(\mult_22/SUMB[13][20] ), .CO(
        \mult_22/CARRYB[14][19] ), .S(\mult_22/SUMB[14][19] ) );
  FA_X1 \mult_22/S2_14_18  ( .A(\mult_22/ab[14][18] ), .B(
        \mult_22/CARRYB[13][18] ), .CI(\mult_22/SUMB[13][19] ), .CO(
        \mult_22/CARRYB[14][18] ), .S(\mult_22/SUMB[14][18] ) );
  FA_X1 \mult_22/S2_14_17  ( .A(\mult_22/ab[14][17] ), .B(
        \mult_22/CARRYB[13][17] ), .CI(\mult_22/SUMB[13][18] ), .CO(
        \mult_22/CARRYB[14][17] ), .S(\mult_22/SUMB[14][17] ) );
  FA_X1 \mult_22/S2_14_16  ( .A(\mult_22/ab[14][16] ), .B(
        \mult_22/CARRYB[13][16] ), .CI(\mult_22/SUMB[13][17] ), .CO(
        \mult_22/CARRYB[14][16] ), .S(\mult_22/SUMB[14][16] ) );
  FA_X1 \mult_22/S2_14_15  ( .A(\mult_22/ab[14][15] ), .B(
        \mult_22/CARRYB[13][15] ), .CI(\mult_22/SUMB[13][16] ), .CO(
        \mult_22/CARRYB[14][15] ), .S(\mult_22/SUMB[14][15] ) );
  FA_X1 \mult_22/S2_14_14  ( .A(\mult_22/ab[14][14] ), .B(
        \mult_22/CARRYB[13][14] ), .CI(\mult_22/SUMB[13][15] ), .CO(
        \mult_22/CARRYB[14][14] ), .S(\mult_22/SUMB[14][14] ) );
  FA_X1 \mult_22/S2_14_13  ( .A(\mult_22/ab[14][13] ), .B(
        \mult_22/CARRYB[13][13] ), .CI(\mult_22/SUMB[13][14] ), .CO(
        \mult_22/CARRYB[14][13] ), .S(\mult_22/SUMB[14][13] ) );
  FA_X1 \mult_22/S2_14_12  ( .A(\mult_22/ab[14][12] ), .B(
        \mult_22/CARRYB[13][12] ), .CI(\mult_22/SUMB[13][13] ), .CO(
        \mult_22/CARRYB[14][12] ), .S(\mult_22/SUMB[14][12] ) );
  FA_X1 \mult_22/S2_14_11  ( .A(\mult_22/ab[14][11] ), .B(
        \mult_22/CARRYB[13][11] ), .CI(\mult_22/SUMB[13][12] ), .CO(
        \mult_22/CARRYB[14][11] ), .S(\mult_22/SUMB[14][11] ) );
  FA_X1 \mult_22/S2_14_10  ( .A(\mult_22/ab[14][10] ), .B(
        \mult_22/CARRYB[13][10] ), .CI(\mult_22/SUMB[13][11] ), .CO(
        \mult_22/CARRYB[14][10] ), .S(\mult_22/SUMB[14][10] ) );
  FA_X1 \mult_22/S2_14_9  ( .A(\mult_22/ab[14][9] ), .B(
        \mult_22/CARRYB[13][9] ), .CI(\mult_22/SUMB[13][10] ), .CO(
        \mult_22/CARRYB[14][9] ), .S(\mult_22/SUMB[14][9] ) );
  FA_X1 \mult_22/S2_14_8  ( .A(\mult_22/ab[14][8] ), .B(
        \mult_22/CARRYB[13][8] ), .CI(\mult_22/SUMB[13][9] ), .CO(
        \mult_22/CARRYB[14][8] ), .S(\mult_22/SUMB[14][8] ) );
  FA_X1 \mult_22/S2_14_7  ( .A(\mult_22/ab[14][7] ), .B(
        \mult_22/CARRYB[13][7] ), .CI(\mult_22/SUMB[13][8] ), .CO(
        \mult_22/CARRYB[14][7] ), .S(\mult_22/SUMB[14][7] ) );
  FA_X1 \mult_22/S2_14_6  ( .A(\mult_22/ab[14][6] ), .B(
        \mult_22/CARRYB[13][6] ), .CI(\mult_22/SUMB[13][7] ), .CO(
        \mult_22/CARRYB[14][6] ), .S(\mult_22/SUMB[14][6] ) );
  FA_X1 \mult_22/S2_14_5  ( .A(\mult_22/ab[14][5] ), .B(
        \mult_22/CARRYB[13][5] ), .CI(\mult_22/SUMB[13][6] ), .CO(
        \mult_22/CARRYB[14][5] ), .S(\mult_22/SUMB[14][5] ) );
  FA_X1 \mult_22/S2_14_4  ( .A(\mult_22/ab[14][4] ), .B(
        \mult_22/CARRYB[13][4] ), .CI(\mult_22/SUMB[13][5] ), .CO(
        \mult_22/CARRYB[14][4] ), .S(\mult_22/SUMB[14][4] ) );
  FA_X1 \mult_22/S2_14_3  ( .A(\mult_22/ab[14][3] ), .B(
        \mult_22/CARRYB[13][3] ), .CI(\mult_22/SUMB[13][4] ), .CO(
        \mult_22/CARRYB[14][3] ), .S(\mult_22/SUMB[14][3] ) );
  FA_X1 \mult_22/S2_14_2  ( .A(\mult_22/ab[14][2] ), .B(
        \mult_22/CARRYB[13][2] ), .CI(\mult_22/SUMB[13][3] ), .CO(
        \mult_22/CARRYB[14][2] ), .S(\mult_22/SUMB[14][2] ) );
  FA_X1 \mult_22/S2_14_1  ( .A(\mult_22/ab[14][1] ), .B(
        \mult_22/CARRYB[13][1] ), .CI(\mult_22/SUMB[13][2] ), .CO(
        \mult_22/CARRYB[14][1] ), .S(\mult_22/SUMB[14][1] ) );
  FA_X1 \mult_22/S1_14_0  ( .A(\mult_22/ab[14][0] ), .B(
        \mult_22/CARRYB[13][0] ), .CI(\mult_22/SUMB[13][1] ), .CO(
        \mult_22/CARRYB[14][0] ), .S(N142) );
  FA_X1 \mult_22/S3_15_62  ( .A(\mult_22/ab[15][62] ), .B(
        \mult_22/CARRYB[14][62] ), .CI(\mult_22/ab[14][63] ), .CO(
        \mult_22/CARRYB[15][62] ), .S(\mult_22/SUMB[15][62] ) );
  FA_X1 \mult_22/S2_15_61  ( .A(\mult_22/ab[15][61] ), .B(
        \mult_22/CARRYB[14][61] ), .CI(\mult_22/SUMB[14][62] ), .CO(
        \mult_22/CARRYB[15][61] ), .S(\mult_22/SUMB[15][61] ) );
  FA_X1 \mult_22/S2_15_60  ( .A(\mult_22/ab[15][60] ), .B(
        \mult_22/CARRYB[14][60] ), .CI(\mult_22/SUMB[14][61] ), .CO(
        \mult_22/CARRYB[15][60] ), .S(\mult_22/SUMB[15][60] ) );
  FA_X1 \mult_22/S2_15_59  ( .A(\mult_22/ab[15][59] ), .B(
        \mult_22/CARRYB[14][59] ), .CI(\mult_22/SUMB[14][60] ), .CO(
        \mult_22/CARRYB[15][59] ), .S(\mult_22/SUMB[15][59] ) );
  FA_X1 \mult_22/S2_15_58  ( .A(\mult_22/ab[15][58] ), .B(
        \mult_22/CARRYB[14][58] ), .CI(\mult_22/SUMB[14][59] ), .CO(
        \mult_22/CARRYB[15][58] ), .S(\mult_22/SUMB[15][58] ) );
  FA_X1 \mult_22/S2_15_57  ( .A(\mult_22/ab[15][57] ), .B(
        \mult_22/CARRYB[14][57] ), .CI(\mult_22/SUMB[14][58] ), .CO(
        \mult_22/CARRYB[15][57] ), .S(\mult_22/SUMB[15][57] ) );
  FA_X1 \mult_22/S2_15_56  ( .A(\mult_22/ab[15][56] ), .B(
        \mult_22/CARRYB[14][56] ), .CI(\mult_22/SUMB[14][57] ), .CO(
        \mult_22/CARRYB[15][56] ), .S(\mult_22/SUMB[15][56] ) );
  FA_X1 \mult_22/S2_15_55  ( .A(\mult_22/ab[15][55] ), .B(
        \mult_22/CARRYB[14][55] ), .CI(\mult_22/SUMB[14][56] ), .CO(
        \mult_22/CARRYB[15][55] ), .S(\mult_22/SUMB[15][55] ) );
  FA_X1 \mult_22/S2_15_54  ( .A(\mult_22/ab[15][54] ), .B(
        \mult_22/CARRYB[14][54] ), .CI(\mult_22/SUMB[14][55] ), .CO(
        \mult_22/CARRYB[15][54] ), .S(\mult_22/SUMB[15][54] ) );
  FA_X1 \mult_22/S2_15_53  ( .A(\mult_22/ab[15][53] ), .B(
        \mult_22/CARRYB[14][53] ), .CI(\mult_22/SUMB[14][54] ), .CO(
        \mult_22/CARRYB[15][53] ), .S(\mult_22/SUMB[15][53] ) );
  FA_X1 \mult_22/S2_15_52  ( .A(\mult_22/CARRYB[14][52] ), .B(
        \mult_22/ab[15][52] ), .CI(\mult_22/SUMB[14][53] ), .CO(
        \mult_22/CARRYB[15][52] ), .S(\mult_22/SUMB[15][52] ) );
  FA_X1 \mult_22/S2_15_51  ( .A(\mult_22/ab[15][51] ), .B(
        \mult_22/CARRYB[14][51] ), .CI(\mult_22/SUMB[14][52] ), .CO(
        \mult_22/CARRYB[15][51] ), .S(\mult_22/SUMB[15][51] ) );
  FA_X1 \mult_22/S2_15_50  ( .A(\mult_22/CARRYB[14][50] ), .B(
        \mult_22/ab[15][50] ), .CI(\mult_22/SUMB[14][51] ), .CO(
        \mult_22/CARRYB[15][50] ), .S(\mult_22/SUMB[15][50] ) );
  FA_X1 \mult_22/S2_15_49  ( .A(\mult_22/CARRYB[14][49] ), .B(
        \mult_22/ab[15][49] ), .CI(\mult_22/SUMB[14][50] ), .CO(
        \mult_22/CARRYB[15][49] ), .S(\mult_22/SUMB[15][49] ) );
  FA_X1 \mult_22/S2_15_48  ( .A(\mult_22/ab[15][48] ), .B(
        \mult_22/CARRYB[14][48] ), .CI(\mult_22/SUMB[14][49] ), .CO(
        \mult_22/CARRYB[15][48] ), .S(\mult_22/SUMB[15][48] ) );
  FA_X1 \mult_22/S2_15_47  ( .A(\mult_22/ab[15][47] ), .B(
        \mult_22/CARRYB[14][47] ), .CI(\mult_22/SUMB[14][48] ), .CO(
        \mult_22/CARRYB[15][47] ), .S(\mult_22/SUMB[15][47] ) );
  FA_X1 \mult_22/S2_15_46  ( .A(\mult_22/ab[15][46] ), .B(
        \mult_22/CARRYB[14][46] ), .CI(\mult_22/SUMB[14][47] ), .CO(
        \mult_22/CARRYB[15][46] ), .S(\mult_22/SUMB[15][46] ) );
  FA_X1 \mult_22/S2_15_45  ( .A(\mult_22/ab[15][45] ), .B(
        \mult_22/CARRYB[14][45] ), .CI(\mult_22/SUMB[14][46] ), .CO(
        \mult_22/CARRYB[15][45] ), .S(\mult_22/SUMB[15][45] ) );
  FA_X1 \mult_22/S2_15_44  ( .A(\mult_22/ab[15][44] ), .B(
        \mult_22/CARRYB[14][44] ), .CI(\mult_22/SUMB[14][45] ), .CO(
        \mult_22/CARRYB[15][44] ), .S(\mult_22/SUMB[15][44] ) );
  FA_X1 \mult_22/S2_15_43  ( .A(\mult_22/ab[15][43] ), .B(
        \mult_22/CARRYB[14][43] ), .CI(\mult_22/SUMB[14][44] ), .CO(
        \mult_22/CARRYB[15][43] ), .S(\mult_22/SUMB[15][43] ) );
  FA_X1 \mult_22/S2_15_42  ( .A(\mult_22/ab[15][42] ), .B(
        \mult_22/CARRYB[14][42] ), .CI(\mult_22/SUMB[14][43] ), .CO(
        \mult_22/CARRYB[15][42] ), .S(\mult_22/SUMB[15][42] ) );
  FA_X1 \mult_22/S2_15_41  ( .A(\mult_22/ab[15][41] ), .B(
        \mult_22/CARRYB[14][41] ), .CI(\mult_22/SUMB[14][42] ), .CO(
        \mult_22/CARRYB[15][41] ), .S(\mult_22/SUMB[15][41] ) );
  FA_X1 \mult_22/S2_15_40  ( .A(\mult_22/ab[15][40] ), .B(
        \mult_22/CARRYB[14][40] ), .CI(\mult_22/SUMB[14][41] ), .CO(
        \mult_22/CARRYB[15][40] ), .S(\mult_22/SUMB[15][40] ) );
  FA_X1 \mult_22/S2_15_39  ( .A(\mult_22/ab[15][39] ), .B(
        \mult_22/CARRYB[14][39] ), .CI(\mult_22/SUMB[14][40] ), .CO(
        \mult_22/CARRYB[15][39] ), .S(\mult_22/SUMB[15][39] ) );
  FA_X1 \mult_22/S2_15_38  ( .A(\mult_22/ab[15][38] ), .B(
        \mult_22/CARRYB[14][38] ), .CI(\mult_22/SUMB[14][39] ), .CO(
        \mult_22/CARRYB[15][38] ), .S(\mult_22/SUMB[15][38] ) );
  FA_X1 \mult_22/S2_15_37  ( .A(\mult_22/ab[15][37] ), .B(
        \mult_22/CARRYB[14][37] ), .CI(\mult_22/SUMB[14][38] ), .CO(
        \mult_22/CARRYB[15][37] ), .S(\mult_22/SUMB[15][37] ) );
  FA_X1 \mult_22/S2_15_36  ( .A(\mult_22/ab[15][36] ), .B(
        \mult_22/CARRYB[14][36] ), .CI(\mult_22/SUMB[14][37] ), .CO(
        \mult_22/CARRYB[15][36] ), .S(\mult_22/SUMB[15][36] ) );
  FA_X1 \mult_22/S2_15_35  ( .A(\mult_22/ab[15][35] ), .B(
        \mult_22/CARRYB[14][35] ), .CI(\mult_22/SUMB[14][36] ), .CO(
        \mult_22/CARRYB[15][35] ), .S(\mult_22/SUMB[15][35] ) );
  FA_X1 \mult_22/S2_15_34  ( .A(\mult_22/ab[15][34] ), .B(
        \mult_22/CARRYB[14][34] ), .CI(\mult_22/SUMB[14][35] ), .CO(
        \mult_22/CARRYB[15][34] ), .S(\mult_22/SUMB[15][34] ) );
  FA_X1 \mult_22/S2_15_33  ( .A(\mult_22/ab[15][33] ), .B(
        \mult_22/CARRYB[14][33] ), .CI(\mult_22/SUMB[14][34] ), .CO(
        \mult_22/CARRYB[15][33] ), .S(\mult_22/SUMB[15][33] ) );
  FA_X1 \mult_22/S2_15_32  ( .A(\mult_22/ab[15][32] ), .B(
        \mult_22/CARRYB[14][32] ), .CI(\mult_22/SUMB[14][33] ), .CO(
        \mult_22/CARRYB[15][32] ), .S(\mult_22/SUMB[15][32] ) );
  FA_X1 \mult_22/S2_15_31  ( .A(\mult_22/ab[15][31] ), .B(
        \mult_22/CARRYB[14][31] ), .CI(\mult_22/SUMB[14][32] ), .CO(
        \mult_22/CARRYB[15][31] ), .S(\mult_22/SUMB[15][31] ) );
  FA_X1 \mult_22/S2_15_30  ( .A(\mult_22/ab[15][30] ), .B(
        \mult_22/CARRYB[14][30] ), .CI(\mult_22/SUMB[14][31] ), .CO(
        \mult_22/CARRYB[15][30] ), .S(\mult_22/SUMB[15][30] ) );
  FA_X1 \mult_22/S2_15_29  ( .A(\mult_22/ab[15][29] ), .B(
        \mult_22/CARRYB[14][29] ), .CI(\mult_22/SUMB[14][30] ), .CO(
        \mult_22/CARRYB[15][29] ), .S(\mult_22/SUMB[15][29] ) );
  FA_X1 \mult_22/S2_15_28  ( .A(\mult_22/ab[15][28] ), .B(
        \mult_22/CARRYB[14][28] ), .CI(\mult_22/SUMB[14][29] ), .CO(
        \mult_22/CARRYB[15][28] ), .S(\mult_22/SUMB[15][28] ) );
  FA_X1 \mult_22/S2_15_27  ( .A(\mult_22/ab[15][27] ), .B(
        \mult_22/CARRYB[14][27] ), .CI(\mult_22/SUMB[14][28] ), .CO(
        \mult_22/CARRYB[15][27] ), .S(\mult_22/SUMB[15][27] ) );
  FA_X1 \mult_22/S2_15_26  ( .A(\mult_22/ab[15][26] ), .B(
        \mult_22/CARRYB[14][26] ), .CI(\mult_22/SUMB[14][27] ), .CO(
        \mult_22/CARRYB[15][26] ), .S(\mult_22/SUMB[15][26] ) );
  FA_X1 \mult_22/S2_15_25  ( .A(\mult_22/ab[15][25] ), .B(
        \mult_22/CARRYB[14][25] ), .CI(\mult_22/SUMB[14][26] ), .CO(
        \mult_22/CARRYB[15][25] ), .S(\mult_22/SUMB[15][25] ) );
  FA_X1 \mult_22/S2_15_24  ( .A(\mult_22/ab[15][24] ), .B(
        \mult_22/CARRYB[14][24] ), .CI(\mult_22/SUMB[14][25] ), .CO(
        \mult_22/CARRYB[15][24] ), .S(\mult_22/SUMB[15][24] ) );
  FA_X1 \mult_22/S2_15_23  ( .A(\mult_22/ab[15][23] ), .B(
        \mult_22/CARRYB[14][23] ), .CI(\mult_22/SUMB[14][24] ), .CO(
        \mult_22/CARRYB[15][23] ), .S(\mult_22/SUMB[15][23] ) );
  FA_X1 \mult_22/S2_15_22  ( .A(\mult_22/ab[15][22] ), .B(
        \mult_22/CARRYB[14][22] ), .CI(\mult_22/SUMB[14][23] ), .CO(
        \mult_22/CARRYB[15][22] ), .S(\mult_22/SUMB[15][22] ) );
  FA_X1 \mult_22/S2_15_21  ( .A(\mult_22/ab[15][21] ), .B(
        \mult_22/CARRYB[14][21] ), .CI(\mult_22/SUMB[14][22] ), .CO(
        \mult_22/CARRYB[15][21] ), .S(\mult_22/SUMB[15][21] ) );
  FA_X1 \mult_22/S2_15_20  ( .A(\mult_22/ab[15][20] ), .B(
        \mult_22/CARRYB[14][20] ), .CI(\mult_22/SUMB[14][21] ), .CO(
        \mult_22/CARRYB[15][20] ), .S(\mult_22/SUMB[15][20] ) );
  FA_X1 \mult_22/S2_15_19  ( .A(\mult_22/ab[15][19] ), .B(
        \mult_22/CARRYB[14][19] ), .CI(\mult_22/SUMB[14][20] ), .CO(
        \mult_22/CARRYB[15][19] ), .S(\mult_22/SUMB[15][19] ) );
  FA_X1 \mult_22/S2_15_18  ( .A(\mult_22/ab[15][18] ), .B(
        \mult_22/CARRYB[14][18] ), .CI(\mult_22/SUMB[14][19] ), .CO(
        \mult_22/CARRYB[15][18] ), .S(\mult_22/SUMB[15][18] ) );
  FA_X1 \mult_22/S2_15_17  ( .A(\mult_22/ab[15][17] ), .B(
        \mult_22/CARRYB[14][17] ), .CI(\mult_22/SUMB[14][18] ), .CO(
        \mult_22/CARRYB[15][17] ), .S(\mult_22/SUMB[15][17] ) );
  FA_X1 \mult_22/S2_15_16  ( .A(\mult_22/ab[15][16] ), .B(
        \mult_22/CARRYB[14][16] ), .CI(\mult_22/SUMB[14][17] ), .CO(
        \mult_22/CARRYB[15][16] ), .S(\mult_22/SUMB[15][16] ) );
  FA_X1 \mult_22/S2_15_15  ( .A(\mult_22/ab[15][15] ), .B(
        \mult_22/CARRYB[14][15] ), .CI(\mult_22/SUMB[14][16] ), .CO(
        \mult_22/CARRYB[15][15] ), .S(\mult_22/SUMB[15][15] ) );
  FA_X1 \mult_22/S2_15_14  ( .A(\mult_22/ab[15][14] ), .B(
        \mult_22/CARRYB[14][14] ), .CI(\mult_22/SUMB[14][15] ), .CO(
        \mult_22/CARRYB[15][14] ), .S(\mult_22/SUMB[15][14] ) );
  FA_X1 \mult_22/S2_15_13  ( .A(\mult_22/ab[15][13] ), .B(
        \mult_22/CARRYB[14][13] ), .CI(\mult_22/SUMB[14][14] ), .CO(
        \mult_22/CARRYB[15][13] ), .S(\mult_22/SUMB[15][13] ) );
  FA_X1 \mult_22/S2_15_12  ( .A(\mult_22/ab[15][12] ), .B(
        \mult_22/CARRYB[14][12] ), .CI(\mult_22/SUMB[14][13] ), .CO(
        \mult_22/CARRYB[15][12] ), .S(\mult_22/SUMB[15][12] ) );
  FA_X1 \mult_22/S2_15_11  ( .A(\mult_22/ab[15][11] ), .B(
        \mult_22/CARRYB[14][11] ), .CI(\mult_22/SUMB[14][12] ), .CO(
        \mult_22/CARRYB[15][11] ), .S(\mult_22/SUMB[15][11] ) );
  FA_X1 \mult_22/S2_15_10  ( .A(\mult_22/ab[15][10] ), .B(
        \mult_22/CARRYB[14][10] ), .CI(\mult_22/SUMB[14][11] ), .CO(
        \mult_22/CARRYB[15][10] ), .S(\mult_22/SUMB[15][10] ) );
  FA_X1 \mult_22/S2_15_9  ( .A(\mult_22/ab[15][9] ), .B(
        \mult_22/CARRYB[14][9] ), .CI(\mult_22/SUMB[14][10] ), .CO(
        \mult_22/CARRYB[15][9] ), .S(\mult_22/SUMB[15][9] ) );
  FA_X1 \mult_22/S2_15_8  ( .A(\mult_22/ab[15][8] ), .B(
        \mult_22/CARRYB[14][8] ), .CI(\mult_22/SUMB[14][9] ), .CO(
        \mult_22/CARRYB[15][8] ), .S(\mult_22/SUMB[15][8] ) );
  FA_X1 \mult_22/S2_15_7  ( .A(\mult_22/ab[15][7] ), .B(
        \mult_22/CARRYB[14][7] ), .CI(\mult_22/SUMB[14][8] ), .CO(
        \mult_22/CARRYB[15][7] ), .S(\mult_22/SUMB[15][7] ) );
  FA_X1 \mult_22/S2_15_6  ( .A(\mult_22/ab[15][6] ), .B(
        \mult_22/CARRYB[14][6] ), .CI(\mult_22/SUMB[14][7] ), .CO(
        \mult_22/CARRYB[15][6] ), .S(\mult_22/SUMB[15][6] ) );
  FA_X1 \mult_22/S2_15_5  ( .A(\mult_22/ab[15][5] ), .B(
        \mult_22/CARRYB[14][5] ), .CI(\mult_22/SUMB[14][6] ), .CO(
        \mult_22/CARRYB[15][5] ), .S(\mult_22/SUMB[15][5] ) );
  FA_X1 \mult_22/S2_15_4  ( .A(\mult_22/ab[15][4] ), .B(
        \mult_22/CARRYB[14][4] ), .CI(\mult_22/SUMB[14][5] ), .CO(
        \mult_22/CARRYB[15][4] ), .S(\mult_22/SUMB[15][4] ) );
  FA_X1 \mult_22/S2_15_3  ( .A(\mult_22/ab[15][3] ), .B(
        \mult_22/CARRYB[14][3] ), .CI(\mult_22/SUMB[14][4] ), .CO(
        \mult_22/CARRYB[15][3] ), .S(\mult_22/SUMB[15][3] ) );
  FA_X1 \mult_22/S2_15_2  ( .A(\mult_22/ab[15][2] ), .B(
        \mult_22/CARRYB[14][2] ), .CI(\mult_22/SUMB[14][3] ), .CO(
        \mult_22/CARRYB[15][2] ), .S(\mult_22/SUMB[15][2] ) );
  FA_X1 \mult_22/S2_15_1  ( .A(\mult_22/ab[15][1] ), .B(
        \mult_22/CARRYB[14][1] ), .CI(\mult_22/SUMB[14][2] ), .CO(
        \mult_22/CARRYB[15][1] ), .S(\mult_22/SUMB[15][1] ) );
  FA_X1 \mult_22/S1_15_0  ( .A(\mult_22/ab[15][0] ), .B(
        \mult_22/CARRYB[14][0] ), .CI(\mult_22/SUMB[14][1] ), .CO(
        \mult_22/CARRYB[15][0] ), .S(N143) );
  FA_X1 \mult_22/S3_16_62  ( .A(\mult_22/ab[16][62] ), .B(
        \mult_22/CARRYB[15][62] ), .CI(\mult_22/ab[15][63] ), .CO(
        \mult_22/CARRYB[16][62] ), .S(\mult_22/SUMB[16][62] ) );
  FA_X1 \mult_22/S2_16_61  ( .A(\mult_22/ab[16][61] ), .B(
        \mult_22/CARRYB[15][61] ), .CI(\mult_22/SUMB[15][62] ), .CO(
        \mult_22/CARRYB[16][61] ), .S(\mult_22/SUMB[16][61] ) );
  FA_X1 \mult_22/S2_16_60  ( .A(\mult_22/ab[16][60] ), .B(
        \mult_22/CARRYB[15][60] ), .CI(\mult_22/SUMB[15][61] ), .CO(
        \mult_22/CARRYB[16][60] ), .S(\mult_22/SUMB[16][60] ) );
  FA_X1 \mult_22/S2_16_59  ( .A(\mult_22/ab[16][59] ), .B(
        \mult_22/CARRYB[15][59] ), .CI(\mult_22/SUMB[15][60] ), .CO(
        \mult_22/CARRYB[16][59] ), .S(\mult_22/SUMB[16][59] ) );
  FA_X1 \mult_22/S2_16_58  ( .A(\mult_22/ab[16][58] ), .B(
        \mult_22/CARRYB[15][58] ), .CI(\mult_22/SUMB[15][59] ), .CO(
        \mult_22/CARRYB[16][58] ), .S(\mult_22/SUMB[16][58] ) );
  FA_X1 \mult_22/S2_16_57  ( .A(\mult_22/ab[16][57] ), .B(
        \mult_22/CARRYB[15][57] ), .CI(\mult_22/SUMB[15][58] ), .CO(
        \mult_22/CARRYB[16][57] ), .S(\mult_22/SUMB[16][57] ) );
  FA_X1 \mult_22/S2_16_56  ( .A(\mult_22/ab[16][56] ), .B(
        \mult_22/CARRYB[15][56] ), .CI(\mult_22/SUMB[15][57] ), .CO(
        \mult_22/CARRYB[16][56] ), .S(\mult_22/SUMB[16][56] ) );
  FA_X1 \mult_22/S2_16_55  ( .A(\mult_22/ab[16][55] ), .B(
        \mult_22/CARRYB[15][55] ), .CI(\mult_22/SUMB[15][56] ), .CO(
        \mult_22/CARRYB[16][55] ), .S(\mult_22/SUMB[16][55] ) );
  FA_X1 \mult_22/S2_16_54  ( .A(\mult_22/ab[16][54] ), .B(
        \mult_22/CARRYB[15][54] ), .CI(\mult_22/SUMB[15][55] ), .CO(
        \mult_22/CARRYB[16][54] ), .S(\mult_22/SUMB[16][54] ) );
  FA_X1 \mult_22/S2_16_53  ( .A(\mult_22/ab[16][53] ), .B(
        \mult_22/CARRYB[15][53] ), .CI(\mult_22/SUMB[15][54] ), .CO(
        \mult_22/CARRYB[16][53] ), .S(\mult_22/SUMB[16][53] ) );
  FA_X1 \mult_22/S2_16_52  ( .A(\mult_22/ab[16][52] ), .B(
        \mult_22/CARRYB[15][52] ), .CI(\mult_22/SUMB[15][53] ), .CO(
        \mult_22/CARRYB[16][52] ), .S(\mult_22/SUMB[16][52] ) );
  FA_X1 \mult_22/S2_16_51  ( .A(\mult_22/ab[16][51] ), .B(
        \mult_22/CARRYB[15][51] ), .CI(\mult_22/SUMB[15][52] ), .CO(
        \mult_22/CARRYB[16][51] ), .S(\mult_22/SUMB[16][51] ) );
  FA_X1 \mult_22/S2_16_50  ( .A(\mult_22/CARRYB[15][50] ), .B(
        \mult_22/ab[16][50] ), .CI(\mult_22/SUMB[15][51] ), .CO(
        \mult_22/CARRYB[16][50] ), .S(\mult_22/SUMB[16][50] ) );
  FA_X1 \mult_22/S2_16_49  ( .A(\mult_22/ab[16][49] ), .B(
        \mult_22/CARRYB[15][49] ), .CI(\mult_22/SUMB[15][50] ), .CO(
        \mult_22/CARRYB[16][49] ), .S(\mult_22/SUMB[16][49] ) );
  FA_X1 \mult_22/S2_16_48  ( .A(\mult_22/CARRYB[15][48] ), .B(
        \mult_22/ab[16][48] ), .CI(\mult_22/SUMB[15][49] ), .CO(
        \mult_22/CARRYB[16][48] ), .S(\mult_22/SUMB[16][48] ) );
  FA_X1 \mult_22/S2_16_47  ( .A(\mult_22/ab[16][47] ), .B(
        \mult_22/CARRYB[15][47] ), .CI(\mult_22/SUMB[15][48] ), .CO(
        \mult_22/CARRYB[16][47] ), .S(\mult_22/SUMB[16][47] ) );
  FA_X1 \mult_22/S2_16_45  ( .A(\mult_22/ab[16][45] ), .B(
        \mult_22/CARRYB[15][45] ), .CI(\mult_22/SUMB[15][46] ), .CO(
        \mult_22/CARRYB[16][45] ), .S(\mult_22/SUMB[16][45] ) );
  FA_X1 \mult_22/S2_16_44  ( .A(\mult_22/ab[16][44] ), .B(
        \mult_22/CARRYB[15][44] ), .CI(\mult_22/SUMB[15][45] ), .CO(
        \mult_22/CARRYB[16][44] ), .S(\mult_22/SUMB[16][44] ) );
  FA_X1 \mult_22/S2_16_42  ( .A(\mult_22/ab[16][42] ), .B(
        \mult_22/CARRYB[15][42] ), .CI(\mult_22/SUMB[15][43] ), .CO(
        \mult_22/CARRYB[16][42] ), .S(\mult_22/SUMB[16][42] ) );
  FA_X1 \mult_22/S2_16_41  ( .A(\mult_22/ab[16][41] ), .B(
        \mult_22/CARRYB[15][41] ), .CI(\mult_22/SUMB[15][42] ), .CO(
        \mult_22/CARRYB[16][41] ), .S(\mult_22/SUMB[16][41] ) );
  FA_X1 \mult_22/S2_16_40  ( .A(\mult_22/ab[16][40] ), .B(
        \mult_22/CARRYB[15][40] ), .CI(\mult_22/SUMB[15][41] ), .CO(
        \mult_22/CARRYB[16][40] ), .S(\mult_22/SUMB[16][40] ) );
  FA_X1 \mult_22/S2_16_39  ( .A(\mult_22/ab[16][39] ), .B(
        \mult_22/CARRYB[15][39] ), .CI(\mult_22/SUMB[15][40] ), .CO(
        \mult_22/CARRYB[16][39] ), .S(\mult_22/SUMB[16][39] ) );
  FA_X1 \mult_22/S2_16_38  ( .A(\mult_22/ab[16][38] ), .B(
        \mult_22/CARRYB[15][38] ), .CI(\mult_22/SUMB[15][39] ), .CO(
        \mult_22/CARRYB[16][38] ), .S(\mult_22/SUMB[16][38] ) );
  FA_X1 \mult_22/S2_16_37  ( .A(\mult_22/ab[16][37] ), .B(
        \mult_22/CARRYB[15][37] ), .CI(\mult_22/SUMB[15][38] ), .CO(
        \mult_22/CARRYB[16][37] ), .S(\mult_22/SUMB[16][37] ) );
  FA_X1 \mult_22/S2_16_36  ( .A(\mult_22/ab[16][36] ), .B(
        \mult_22/CARRYB[15][36] ), .CI(\mult_22/SUMB[15][37] ), .CO(
        \mult_22/CARRYB[16][36] ), .S(\mult_22/SUMB[16][36] ) );
  FA_X1 \mult_22/S2_16_35  ( .A(\mult_22/ab[16][35] ), .B(
        \mult_22/CARRYB[15][35] ), .CI(\mult_22/SUMB[15][36] ), .CO(
        \mult_22/CARRYB[16][35] ), .S(\mult_22/SUMB[16][35] ) );
  FA_X1 \mult_22/S2_16_34  ( .A(\mult_22/ab[16][34] ), .B(
        \mult_22/CARRYB[15][34] ), .CI(\mult_22/SUMB[15][35] ), .CO(
        \mult_22/CARRYB[16][34] ), .S(\mult_22/SUMB[16][34] ) );
  FA_X1 \mult_22/S2_16_33  ( .A(\mult_22/ab[16][33] ), .B(
        \mult_22/CARRYB[15][33] ), .CI(\mult_22/SUMB[15][34] ), .CO(
        \mult_22/CARRYB[16][33] ), .S(\mult_22/SUMB[16][33] ) );
  FA_X1 \mult_22/S2_16_32  ( .A(\mult_22/ab[16][32] ), .B(
        \mult_22/CARRYB[15][32] ), .CI(\mult_22/SUMB[15][33] ), .CO(
        \mult_22/CARRYB[16][32] ), .S(\mult_22/SUMB[16][32] ) );
  FA_X1 \mult_22/S2_16_31  ( .A(\mult_22/ab[16][31] ), .B(
        \mult_22/CARRYB[15][31] ), .CI(\mult_22/SUMB[15][32] ), .CO(
        \mult_22/CARRYB[16][31] ), .S(\mult_22/SUMB[16][31] ) );
  FA_X1 \mult_22/S2_16_30  ( .A(\mult_22/ab[16][30] ), .B(
        \mult_22/CARRYB[15][30] ), .CI(\mult_22/SUMB[15][31] ), .CO(
        \mult_22/CARRYB[16][30] ), .S(\mult_22/SUMB[16][30] ) );
  FA_X1 \mult_22/S2_16_29  ( .A(\mult_22/ab[16][29] ), .B(
        \mult_22/CARRYB[15][29] ), .CI(\mult_22/SUMB[15][30] ), .CO(
        \mult_22/CARRYB[16][29] ), .S(\mult_22/SUMB[16][29] ) );
  FA_X1 \mult_22/S2_16_28  ( .A(\mult_22/ab[16][28] ), .B(
        \mult_22/CARRYB[15][28] ), .CI(\mult_22/SUMB[15][29] ), .CO(
        \mult_22/CARRYB[16][28] ), .S(\mult_22/SUMB[16][28] ) );
  FA_X1 \mult_22/S2_16_27  ( .A(\mult_22/ab[16][27] ), .B(
        \mult_22/CARRYB[15][27] ), .CI(\mult_22/SUMB[15][28] ), .CO(
        \mult_22/CARRYB[16][27] ), .S(\mult_22/SUMB[16][27] ) );
  FA_X1 \mult_22/S2_16_26  ( .A(\mult_22/ab[16][26] ), .B(
        \mult_22/CARRYB[15][26] ), .CI(\mult_22/SUMB[15][27] ), .CO(
        \mult_22/CARRYB[16][26] ), .S(\mult_22/SUMB[16][26] ) );
  FA_X1 \mult_22/S2_16_25  ( .A(\mult_22/ab[16][25] ), .B(
        \mult_22/CARRYB[15][25] ), .CI(\mult_22/SUMB[15][26] ), .CO(
        \mult_22/CARRYB[16][25] ), .S(\mult_22/SUMB[16][25] ) );
  FA_X1 \mult_22/S2_16_24  ( .A(\mult_22/ab[16][24] ), .B(
        \mult_22/CARRYB[15][24] ), .CI(\mult_22/SUMB[15][25] ), .CO(
        \mult_22/CARRYB[16][24] ), .S(\mult_22/SUMB[16][24] ) );
  FA_X1 \mult_22/S2_16_23  ( .A(\mult_22/ab[16][23] ), .B(
        \mult_22/CARRYB[15][23] ), .CI(\mult_22/SUMB[15][24] ), .CO(
        \mult_22/CARRYB[16][23] ), .S(\mult_22/SUMB[16][23] ) );
  FA_X1 \mult_22/S2_16_22  ( .A(\mult_22/ab[16][22] ), .B(
        \mult_22/CARRYB[15][22] ), .CI(\mult_22/SUMB[15][23] ), .CO(
        \mult_22/CARRYB[16][22] ), .S(\mult_22/SUMB[16][22] ) );
  FA_X1 \mult_22/S2_16_21  ( .A(\mult_22/ab[16][21] ), .B(
        \mult_22/CARRYB[15][21] ), .CI(\mult_22/SUMB[15][22] ), .CO(
        \mult_22/CARRYB[16][21] ), .S(\mult_22/SUMB[16][21] ) );
  FA_X1 \mult_22/S2_16_20  ( .A(\mult_22/ab[16][20] ), .B(
        \mult_22/CARRYB[15][20] ), .CI(\mult_22/SUMB[15][21] ), .CO(
        \mult_22/CARRYB[16][20] ), .S(\mult_22/SUMB[16][20] ) );
  FA_X1 \mult_22/S2_16_19  ( .A(\mult_22/ab[16][19] ), .B(
        \mult_22/CARRYB[15][19] ), .CI(\mult_22/SUMB[15][20] ), .CO(
        \mult_22/CARRYB[16][19] ), .S(\mult_22/SUMB[16][19] ) );
  FA_X1 \mult_22/S2_16_18  ( .A(\mult_22/ab[16][18] ), .B(
        \mult_22/CARRYB[15][18] ), .CI(\mult_22/SUMB[15][19] ), .CO(
        \mult_22/CARRYB[16][18] ), .S(\mult_22/SUMB[16][18] ) );
  FA_X1 \mult_22/S2_16_17  ( .A(\mult_22/ab[16][17] ), .B(
        \mult_22/CARRYB[15][17] ), .CI(\mult_22/SUMB[15][18] ), .CO(
        \mult_22/CARRYB[16][17] ), .S(\mult_22/SUMB[16][17] ) );
  FA_X1 \mult_22/S2_16_16  ( .A(\mult_22/ab[16][16] ), .B(
        \mult_22/CARRYB[15][16] ), .CI(\mult_22/SUMB[15][17] ), .CO(
        \mult_22/CARRYB[16][16] ), .S(\mult_22/SUMB[16][16] ) );
  FA_X1 \mult_22/S2_16_15  ( .A(\mult_22/ab[16][15] ), .B(
        \mult_22/CARRYB[15][15] ), .CI(\mult_22/SUMB[15][16] ), .CO(
        \mult_22/CARRYB[16][15] ), .S(\mult_22/SUMB[16][15] ) );
  FA_X1 \mult_22/S2_16_14  ( .A(\mult_22/ab[16][14] ), .B(
        \mult_22/CARRYB[15][14] ), .CI(\mult_22/SUMB[15][15] ), .CO(
        \mult_22/CARRYB[16][14] ), .S(\mult_22/SUMB[16][14] ) );
  FA_X1 \mult_22/S2_16_13  ( .A(\mult_22/ab[16][13] ), .B(
        \mult_22/CARRYB[15][13] ), .CI(\mult_22/SUMB[15][14] ), .CO(
        \mult_22/CARRYB[16][13] ), .S(\mult_22/SUMB[16][13] ) );
  FA_X1 \mult_22/S2_16_12  ( .A(\mult_22/ab[16][12] ), .B(
        \mult_22/CARRYB[15][12] ), .CI(\mult_22/SUMB[15][13] ), .CO(
        \mult_22/CARRYB[16][12] ), .S(\mult_22/SUMB[16][12] ) );
  FA_X1 \mult_22/S2_16_11  ( .A(\mult_22/ab[16][11] ), .B(
        \mult_22/CARRYB[15][11] ), .CI(\mult_22/SUMB[15][12] ), .CO(
        \mult_22/CARRYB[16][11] ), .S(\mult_22/SUMB[16][11] ) );
  FA_X1 \mult_22/S2_16_10  ( .A(\mult_22/ab[16][10] ), .B(
        \mult_22/CARRYB[15][10] ), .CI(\mult_22/SUMB[15][11] ), .CO(
        \mult_22/CARRYB[16][10] ), .S(\mult_22/SUMB[16][10] ) );
  FA_X1 \mult_22/S2_16_9  ( .A(\mult_22/ab[16][9] ), .B(
        \mult_22/CARRYB[15][9] ), .CI(\mult_22/SUMB[15][10] ), .CO(
        \mult_22/CARRYB[16][9] ), .S(\mult_22/SUMB[16][9] ) );
  FA_X1 \mult_22/S2_16_8  ( .A(\mult_22/ab[16][8] ), .B(
        \mult_22/CARRYB[15][8] ), .CI(\mult_22/SUMB[15][9] ), .CO(
        \mult_22/CARRYB[16][8] ), .S(\mult_22/SUMB[16][8] ) );
  FA_X1 \mult_22/S2_16_7  ( .A(\mult_22/ab[16][7] ), .B(
        \mult_22/CARRYB[15][7] ), .CI(\mult_22/SUMB[15][8] ), .CO(
        \mult_22/CARRYB[16][7] ), .S(\mult_22/SUMB[16][7] ) );
  FA_X1 \mult_22/S2_16_6  ( .A(\mult_22/ab[16][6] ), .B(
        \mult_22/CARRYB[15][6] ), .CI(\mult_22/SUMB[15][7] ), .CO(
        \mult_22/CARRYB[16][6] ), .S(\mult_22/SUMB[16][6] ) );
  FA_X1 \mult_22/S2_16_5  ( .A(\mult_22/ab[16][5] ), .B(
        \mult_22/CARRYB[15][5] ), .CI(\mult_22/SUMB[15][6] ), .CO(
        \mult_22/CARRYB[16][5] ), .S(\mult_22/SUMB[16][5] ) );
  FA_X1 \mult_22/S2_16_4  ( .A(\mult_22/ab[16][4] ), .B(
        \mult_22/CARRYB[15][4] ), .CI(\mult_22/SUMB[15][5] ), .CO(
        \mult_22/CARRYB[16][4] ), .S(\mult_22/SUMB[16][4] ) );
  FA_X1 \mult_22/S2_16_3  ( .A(\mult_22/ab[16][3] ), .B(
        \mult_22/CARRYB[15][3] ), .CI(\mult_22/SUMB[15][4] ), .CO(
        \mult_22/CARRYB[16][3] ), .S(\mult_22/SUMB[16][3] ) );
  FA_X1 \mult_22/S2_16_2  ( .A(\mult_22/ab[16][2] ), .B(
        \mult_22/CARRYB[15][2] ), .CI(\mult_22/SUMB[15][3] ), .CO(
        \mult_22/CARRYB[16][2] ), .S(\mult_22/SUMB[16][2] ) );
  FA_X1 \mult_22/S2_16_1  ( .A(\mult_22/ab[16][1] ), .B(
        \mult_22/CARRYB[15][1] ), .CI(\mult_22/SUMB[15][2] ), .CO(
        \mult_22/CARRYB[16][1] ), .S(\mult_22/SUMB[16][1] ) );
  FA_X1 \mult_22/S1_16_0  ( .A(\mult_22/ab[16][0] ), .B(
        \mult_22/CARRYB[15][0] ), .CI(\mult_22/SUMB[15][1] ), .CO(
        \mult_22/CARRYB[16][0] ), .S(N144) );
  FA_X1 \mult_22/S3_17_62  ( .A(\mult_22/ab[17][62] ), .B(
        \mult_22/CARRYB[16][62] ), .CI(\mult_22/ab[16][63] ), .CO(
        \mult_22/CARRYB[17][62] ), .S(\mult_22/SUMB[17][62] ) );
  FA_X1 \mult_22/S2_17_61  ( .A(\mult_22/ab[17][61] ), .B(
        \mult_22/CARRYB[16][61] ), .CI(\mult_22/SUMB[16][62] ), .CO(
        \mult_22/CARRYB[17][61] ), .S(\mult_22/SUMB[17][61] ) );
  FA_X1 \mult_22/S2_17_60  ( .A(\mult_22/ab[17][60] ), .B(
        \mult_22/CARRYB[16][60] ), .CI(\mult_22/SUMB[16][61] ), .CO(
        \mult_22/CARRYB[17][60] ), .S(\mult_22/SUMB[17][60] ) );
  FA_X1 \mult_22/S2_17_59  ( .A(\mult_22/ab[17][59] ), .B(
        \mult_22/CARRYB[16][59] ), .CI(\mult_22/SUMB[16][60] ), .CO(
        \mult_22/CARRYB[17][59] ), .S(\mult_22/SUMB[17][59] ) );
  FA_X1 \mult_22/S2_17_58  ( .A(\mult_22/ab[17][58] ), .B(
        \mult_22/CARRYB[16][58] ), .CI(\mult_22/SUMB[16][59] ), .CO(
        \mult_22/CARRYB[17][58] ), .S(\mult_22/SUMB[17][58] ) );
  FA_X1 \mult_22/S2_17_57  ( .A(\mult_22/ab[17][57] ), .B(
        \mult_22/CARRYB[16][57] ), .CI(\mult_22/SUMB[16][58] ), .CO(
        \mult_22/CARRYB[17][57] ), .S(\mult_22/SUMB[17][57] ) );
  FA_X1 \mult_22/S2_17_56  ( .A(\mult_22/ab[17][56] ), .B(
        \mult_22/CARRYB[16][56] ), .CI(\mult_22/SUMB[16][57] ), .CO(
        \mult_22/CARRYB[17][56] ), .S(\mult_22/SUMB[17][56] ) );
  FA_X1 \mult_22/S2_17_55  ( .A(\mult_22/ab[17][55] ), .B(
        \mult_22/CARRYB[16][55] ), .CI(\mult_22/SUMB[16][56] ), .CO(
        \mult_22/CARRYB[17][55] ), .S(\mult_22/SUMB[17][55] ) );
  FA_X1 \mult_22/S2_17_54  ( .A(\mult_22/ab[17][54] ), .B(
        \mult_22/CARRYB[16][54] ), .CI(\mult_22/SUMB[16][55] ), .CO(
        \mult_22/CARRYB[17][54] ), .S(\mult_22/SUMB[17][54] ) );
  FA_X1 \mult_22/S2_17_53  ( .A(\mult_22/ab[17][53] ), .B(
        \mult_22/CARRYB[16][53] ), .CI(\mult_22/SUMB[16][54] ), .CO(
        \mult_22/CARRYB[17][53] ), .S(\mult_22/SUMB[17][53] ) );
  FA_X1 \mult_22/S2_17_52  ( .A(\mult_22/ab[17][52] ), .B(
        \mult_22/CARRYB[16][52] ), .CI(\mult_22/SUMB[16][53] ), .CO(
        \mult_22/CARRYB[17][52] ), .S(\mult_22/SUMB[17][52] ) );
  FA_X1 \mult_22/S2_17_51  ( .A(\mult_22/ab[17][51] ), .B(
        \mult_22/CARRYB[16][51] ), .CI(\mult_22/SUMB[16][52] ), .CO(
        \mult_22/CARRYB[17][51] ), .S(\mult_22/SUMB[17][51] ) );
  FA_X1 \mult_22/S2_17_50  ( .A(\mult_22/CARRYB[16][50] ), .B(
        \mult_22/ab[17][50] ), .CI(\mult_22/SUMB[16][51] ), .CO(
        \mult_22/CARRYB[17][50] ), .S(\mult_22/SUMB[17][50] ) );
  FA_X1 \mult_22/S2_17_49  ( .A(\mult_22/ab[17][49] ), .B(
        \mult_22/CARRYB[16][49] ), .CI(\mult_22/SUMB[16][50] ), .CO(
        \mult_22/CARRYB[17][49] ), .S(\mult_22/SUMB[17][49] ) );
  FA_X1 \mult_22/S2_17_48  ( .A(\mult_22/CARRYB[16][48] ), .B(
        \mult_22/ab[17][48] ), .CI(\mult_22/SUMB[16][49] ), .CO(
        \mult_22/CARRYB[17][48] ), .S(\mult_22/SUMB[17][48] ) );
  FA_X1 \mult_22/S2_17_47  ( .A(\mult_22/ab[17][47] ), .B(
        \mult_22/CARRYB[16][47] ), .CI(\mult_22/SUMB[16][48] ), .CO(
        \mult_22/CARRYB[17][47] ), .S(\mult_22/SUMB[17][47] ) );
  FA_X1 \mult_22/S2_17_45  ( .A(\mult_22/ab[17][45] ), .B(
        \mult_22/CARRYB[16][45] ), .CI(\mult_22/SUMB[16][46] ), .CO(
        \mult_22/CARRYB[17][45] ), .S(\mult_22/SUMB[17][45] ) );
  FA_X1 \mult_22/S2_17_44  ( .A(\mult_22/ab[17][44] ), .B(
        \mult_22/CARRYB[16][44] ), .CI(\mult_22/SUMB[16][45] ), .CO(
        \mult_22/CARRYB[17][44] ), .S(\mult_22/SUMB[17][44] ) );
  FA_X1 \mult_22/S2_17_43  ( .A(\mult_22/ab[17][43] ), .B(
        \mult_22/CARRYB[16][43] ), .CI(\mult_22/SUMB[16][44] ), .CO(
        \mult_22/CARRYB[17][43] ), .S(\mult_22/SUMB[17][43] ) );
  FA_X1 \mult_22/S2_17_41  ( .A(\mult_22/ab[17][41] ), .B(
        \mult_22/CARRYB[16][41] ), .CI(\mult_22/SUMB[16][42] ), .CO(
        \mult_22/CARRYB[17][41] ), .S(\mult_22/SUMB[17][41] ) );
  FA_X1 \mult_22/S2_17_40  ( .A(\mult_22/ab[17][40] ), .B(
        \mult_22/CARRYB[16][40] ), .CI(\mult_22/SUMB[16][41] ), .CO(
        \mult_22/CARRYB[17][40] ), .S(\mult_22/SUMB[17][40] ) );
  FA_X1 \mult_22/S2_17_39  ( .A(\mult_22/ab[17][39] ), .B(
        \mult_22/CARRYB[16][39] ), .CI(\mult_22/SUMB[16][40] ), .CO(
        \mult_22/CARRYB[17][39] ), .S(\mult_22/SUMB[17][39] ) );
  FA_X1 \mult_22/S2_17_38  ( .A(\mult_22/ab[17][38] ), .B(
        \mult_22/CARRYB[16][38] ), .CI(\mult_22/SUMB[16][39] ), .CO(
        \mult_22/CARRYB[17][38] ), .S(\mult_22/SUMB[17][38] ) );
  FA_X1 \mult_22/S2_17_37  ( .A(\mult_22/ab[17][37] ), .B(
        \mult_22/CARRYB[16][37] ), .CI(\mult_22/SUMB[16][38] ), .CO(
        \mult_22/CARRYB[17][37] ), .S(\mult_22/SUMB[17][37] ) );
  FA_X1 \mult_22/S2_17_36  ( .A(\mult_22/ab[17][36] ), .B(
        \mult_22/CARRYB[16][36] ), .CI(\mult_22/SUMB[16][37] ), .CO(
        \mult_22/CARRYB[17][36] ), .S(\mult_22/SUMB[17][36] ) );
  FA_X1 \mult_22/S2_17_35  ( .A(\mult_22/ab[17][35] ), .B(
        \mult_22/CARRYB[16][35] ), .CI(\mult_22/SUMB[16][36] ), .CO(
        \mult_22/CARRYB[17][35] ), .S(\mult_22/SUMB[17][35] ) );
  FA_X1 \mult_22/S2_17_34  ( .A(\mult_22/ab[17][34] ), .B(
        \mult_22/CARRYB[16][34] ), .CI(\mult_22/SUMB[16][35] ), .CO(
        \mult_22/CARRYB[17][34] ), .S(\mult_22/SUMB[17][34] ) );
  FA_X1 \mult_22/S2_17_33  ( .A(\mult_22/ab[17][33] ), .B(
        \mult_22/CARRYB[16][33] ), .CI(\mult_22/SUMB[16][34] ), .CO(
        \mult_22/CARRYB[17][33] ), .S(\mult_22/SUMB[17][33] ) );
  FA_X1 \mult_22/S2_17_32  ( .A(\mult_22/ab[17][32] ), .B(
        \mult_22/CARRYB[16][32] ), .CI(\mult_22/SUMB[16][33] ), .CO(
        \mult_22/CARRYB[17][32] ), .S(\mult_22/SUMB[17][32] ) );
  FA_X1 \mult_22/S2_17_31  ( .A(\mult_22/ab[17][31] ), .B(
        \mult_22/CARRYB[16][31] ), .CI(\mult_22/SUMB[16][32] ), .CO(
        \mult_22/CARRYB[17][31] ), .S(\mult_22/SUMB[17][31] ) );
  FA_X1 \mult_22/S2_17_30  ( .A(\mult_22/ab[17][30] ), .B(
        \mult_22/CARRYB[16][30] ), .CI(\mult_22/SUMB[16][31] ), .CO(
        \mult_22/CARRYB[17][30] ), .S(\mult_22/SUMB[17][30] ) );
  FA_X1 \mult_22/S2_17_29  ( .A(\mult_22/ab[17][29] ), .B(
        \mult_22/CARRYB[16][29] ), .CI(\mult_22/SUMB[16][30] ), .CO(
        \mult_22/CARRYB[17][29] ), .S(\mult_22/SUMB[17][29] ) );
  FA_X1 \mult_22/S2_17_28  ( .A(\mult_22/ab[17][28] ), .B(
        \mult_22/CARRYB[16][28] ), .CI(\mult_22/SUMB[16][29] ), .CO(
        \mult_22/CARRYB[17][28] ), .S(\mult_22/SUMB[17][28] ) );
  FA_X1 \mult_22/S2_17_27  ( .A(\mult_22/ab[17][27] ), .B(
        \mult_22/CARRYB[16][27] ), .CI(\mult_22/SUMB[16][28] ), .CO(
        \mult_22/CARRYB[17][27] ), .S(\mult_22/SUMB[17][27] ) );
  FA_X1 \mult_22/S2_17_26  ( .A(\mult_22/ab[17][26] ), .B(
        \mult_22/CARRYB[16][26] ), .CI(\mult_22/SUMB[16][27] ), .CO(
        \mult_22/CARRYB[17][26] ), .S(\mult_22/SUMB[17][26] ) );
  FA_X1 \mult_22/S2_17_25  ( .A(\mult_22/ab[17][25] ), .B(
        \mult_22/CARRYB[16][25] ), .CI(\mult_22/SUMB[16][26] ), .CO(
        \mult_22/CARRYB[17][25] ), .S(\mult_22/SUMB[17][25] ) );
  FA_X1 \mult_22/S2_17_24  ( .A(\mult_22/ab[17][24] ), .B(
        \mult_22/CARRYB[16][24] ), .CI(\mult_22/SUMB[16][25] ), .CO(
        \mult_22/CARRYB[17][24] ), .S(\mult_22/SUMB[17][24] ) );
  FA_X1 \mult_22/S2_17_23  ( .A(\mult_22/ab[17][23] ), .B(
        \mult_22/CARRYB[16][23] ), .CI(\mult_22/SUMB[16][24] ), .CO(
        \mult_22/CARRYB[17][23] ), .S(\mult_22/SUMB[17][23] ) );
  FA_X1 \mult_22/S2_17_22  ( .A(\mult_22/ab[17][22] ), .B(
        \mult_22/CARRYB[16][22] ), .CI(\mult_22/SUMB[16][23] ), .CO(
        \mult_22/CARRYB[17][22] ), .S(\mult_22/SUMB[17][22] ) );
  FA_X1 \mult_22/S2_17_21  ( .A(\mult_22/ab[17][21] ), .B(
        \mult_22/CARRYB[16][21] ), .CI(\mult_22/SUMB[16][22] ), .CO(
        \mult_22/CARRYB[17][21] ), .S(\mult_22/SUMB[17][21] ) );
  FA_X1 \mult_22/S2_17_20  ( .A(\mult_22/ab[17][20] ), .B(
        \mult_22/CARRYB[16][20] ), .CI(\mult_22/SUMB[16][21] ), .CO(
        \mult_22/CARRYB[17][20] ), .S(\mult_22/SUMB[17][20] ) );
  FA_X1 \mult_22/S2_17_19  ( .A(\mult_22/ab[17][19] ), .B(
        \mult_22/CARRYB[16][19] ), .CI(\mult_22/SUMB[16][20] ), .CO(
        \mult_22/CARRYB[17][19] ), .S(\mult_22/SUMB[17][19] ) );
  FA_X1 \mult_22/S2_17_18  ( .A(\mult_22/ab[17][18] ), .B(
        \mult_22/CARRYB[16][18] ), .CI(\mult_22/SUMB[16][19] ), .CO(
        \mult_22/CARRYB[17][18] ), .S(\mult_22/SUMB[17][18] ) );
  FA_X1 \mult_22/S2_17_17  ( .A(\mult_22/ab[17][17] ), .B(
        \mult_22/CARRYB[16][17] ), .CI(\mult_22/SUMB[16][18] ), .CO(
        \mult_22/CARRYB[17][17] ), .S(\mult_22/SUMB[17][17] ) );
  FA_X1 \mult_22/S2_17_16  ( .A(\mult_22/ab[17][16] ), .B(
        \mult_22/CARRYB[16][16] ), .CI(\mult_22/SUMB[16][17] ), .CO(
        \mult_22/CARRYB[17][16] ), .S(\mult_22/SUMB[17][16] ) );
  FA_X1 \mult_22/S2_17_15  ( .A(\mult_22/ab[17][15] ), .B(
        \mult_22/CARRYB[16][15] ), .CI(\mult_22/SUMB[16][16] ), .CO(
        \mult_22/CARRYB[17][15] ), .S(\mult_22/SUMB[17][15] ) );
  FA_X1 \mult_22/S2_17_14  ( .A(\mult_22/ab[17][14] ), .B(
        \mult_22/CARRYB[16][14] ), .CI(\mult_22/SUMB[16][15] ), .CO(
        \mult_22/CARRYB[17][14] ), .S(\mult_22/SUMB[17][14] ) );
  FA_X1 \mult_22/S2_17_13  ( .A(\mult_22/ab[17][13] ), .B(
        \mult_22/CARRYB[16][13] ), .CI(\mult_22/SUMB[16][14] ), .CO(
        \mult_22/CARRYB[17][13] ), .S(\mult_22/SUMB[17][13] ) );
  FA_X1 \mult_22/S2_17_12  ( .A(\mult_22/ab[17][12] ), .B(
        \mult_22/CARRYB[16][12] ), .CI(\mult_22/SUMB[16][13] ), .CO(
        \mult_22/CARRYB[17][12] ), .S(\mult_22/SUMB[17][12] ) );
  FA_X1 \mult_22/S2_17_11  ( .A(\mult_22/ab[17][11] ), .B(
        \mult_22/CARRYB[16][11] ), .CI(\mult_22/SUMB[16][12] ), .CO(
        \mult_22/CARRYB[17][11] ), .S(\mult_22/SUMB[17][11] ) );
  FA_X1 \mult_22/S2_17_10  ( .A(\mult_22/ab[17][10] ), .B(
        \mult_22/CARRYB[16][10] ), .CI(\mult_22/SUMB[16][11] ), .CO(
        \mult_22/CARRYB[17][10] ), .S(\mult_22/SUMB[17][10] ) );
  FA_X1 \mult_22/S2_17_9  ( .A(\mult_22/ab[17][9] ), .B(
        \mult_22/CARRYB[16][9] ), .CI(\mult_22/SUMB[16][10] ), .CO(
        \mult_22/CARRYB[17][9] ), .S(\mult_22/SUMB[17][9] ) );
  FA_X1 \mult_22/S2_17_8  ( .A(\mult_22/ab[17][8] ), .B(
        \mult_22/CARRYB[16][8] ), .CI(\mult_22/SUMB[16][9] ), .CO(
        \mult_22/CARRYB[17][8] ), .S(\mult_22/SUMB[17][8] ) );
  FA_X1 \mult_22/S2_17_7  ( .A(\mult_22/ab[17][7] ), .B(
        \mult_22/CARRYB[16][7] ), .CI(\mult_22/SUMB[16][8] ), .CO(
        \mult_22/CARRYB[17][7] ), .S(\mult_22/SUMB[17][7] ) );
  FA_X1 \mult_22/S2_17_6  ( .A(\mult_22/ab[17][6] ), .B(
        \mult_22/CARRYB[16][6] ), .CI(\mult_22/SUMB[16][7] ), .CO(
        \mult_22/CARRYB[17][6] ), .S(\mult_22/SUMB[17][6] ) );
  FA_X1 \mult_22/S2_17_5  ( .A(\mult_22/ab[17][5] ), .B(
        \mult_22/CARRYB[16][5] ), .CI(\mult_22/SUMB[16][6] ), .CO(
        \mult_22/CARRYB[17][5] ), .S(\mult_22/SUMB[17][5] ) );
  FA_X1 \mult_22/S2_17_4  ( .A(\mult_22/ab[17][4] ), .B(
        \mult_22/CARRYB[16][4] ), .CI(\mult_22/SUMB[16][5] ), .CO(
        \mult_22/CARRYB[17][4] ), .S(\mult_22/SUMB[17][4] ) );
  FA_X1 \mult_22/S2_17_3  ( .A(\mult_22/ab[17][3] ), .B(
        \mult_22/CARRYB[16][3] ), .CI(\mult_22/SUMB[16][4] ), .CO(
        \mult_22/CARRYB[17][3] ), .S(\mult_22/SUMB[17][3] ) );
  FA_X1 \mult_22/S2_17_2  ( .A(\mult_22/ab[17][2] ), .B(
        \mult_22/CARRYB[16][2] ), .CI(\mult_22/SUMB[16][3] ), .CO(
        \mult_22/CARRYB[17][2] ), .S(\mult_22/SUMB[17][2] ) );
  FA_X1 \mult_22/S2_17_1  ( .A(\mult_22/ab[17][1] ), .B(
        \mult_22/CARRYB[16][1] ), .CI(\mult_22/SUMB[16][2] ), .CO(
        \mult_22/CARRYB[17][1] ), .S(\mult_22/SUMB[17][1] ) );
  FA_X1 \mult_22/S1_17_0  ( .A(\mult_22/ab[17][0] ), .B(
        \mult_22/CARRYB[16][0] ), .CI(\mult_22/SUMB[16][1] ), .CO(
        \mult_22/CARRYB[17][0] ), .S(N145) );
  FA_X1 \mult_22/S3_18_62  ( .A(\mult_22/ab[18][62] ), .B(
        \mult_22/CARRYB[17][62] ), .CI(\mult_22/ab[17][63] ), .CO(
        \mult_22/CARRYB[18][62] ), .S(\mult_22/SUMB[18][62] ) );
  FA_X1 \mult_22/S2_18_61  ( .A(\mult_22/ab[18][61] ), .B(
        \mult_22/CARRYB[17][61] ), .CI(\mult_22/SUMB[17][62] ), .CO(
        \mult_22/CARRYB[18][61] ), .S(\mult_22/SUMB[18][61] ) );
  FA_X1 \mult_22/S2_18_60  ( .A(\mult_22/ab[18][60] ), .B(
        \mult_22/CARRYB[17][60] ), .CI(\mult_22/SUMB[17][61] ), .CO(
        \mult_22/CARRYB[18][60] ), .S(\mult_22/SUMB[18][60] ) );
  FA_X1 \mult_22/S2_18_59  ( .A(\mult_22/ab[18][59] ), .B(
        \mult_22/CARRYB[17][59] ), .CI(\mult_22/SUMB[17][60] ), .CO(
        \mult_22/CARRYB[18][59] ), .S(\mult_22/SUMB[18][59] ) );
  FA_X1 \mult_22/S2_18_58  ( .A(\mult_22/ab[18][58] ), .B(
        \mult_22/CARRYB[17][58] ), .CI(\mult_22/SUMB[17][59] ), .CO(
        \mult_22/CARRYB[18][58] ), .S(\mult_22/SUMB[18][58] ) );
  FA_X1 \mult_22/S2_18_57  ( .A(\mult_22/ab[18][57] ), .B(
        \mult_22/CARRYB[17][57] ), .CI(\mult_22/SUMB[17][58] ), .CO(
        \mult_22/CARRYB[18][57] ), .S(\mult_22/SUMB[18][57] ) );
  FA_X1 \mult_22/S2_18_56  ( .A(\mult_22/ab[18][56] ), .B(
        \mult_22/CARRYB[17][56] ), .CI(\mult_22/SUMB[17][57] ), .CO(
        \mult_22/CARRYB[18][56] ), .S(\mult_22/SUMB[18][56] ) );
  FA_X1 \mult_22/S2_18_55  ( .A(\mult_22/ab[18][55] ), .B(
        \mult_22/CARRYB[17][55] ), .CI(\mult_22/SUMB[17][56] ), .CO(
        \mult_22/CARRYB[18][55] ), .S(\mult_22/SUMB[18][55] ) );
  FA_X1 \mult_22/S2_18_54  ( .A(\mult_22/ab[18][54] ), .B(
        \mult_22/CARRYB[17][54] ), .CI(\mult_22/SUMB[17][55] ), .CO(
        \mult_22/CARRYB[18][54] ), .S(\mult_22/SUMB[18][54] ) );
  FA_X1 \mult_22/S2_18_53  ( .A(\mult_22/ab[18][53] ), .B(
        \mult_22/CARRYB[17][53] ), .CI(\mult_22/SUMB[17][54] ), .CO(
        \mult_22/CARRYB[18][53] ), .S(\mult_22/SUMB[18][53] ) );
  FA_X1 \mult_22/S2_18_52  ( .A(\mult_22/ab[18][52] ), .B(
        \mult_22/CARRYB[17][52] ), .CI(\mult_22/SUMB[17][53] ), .CO(
        \mult_22/CARRYB[18][52] ), .S(\mult_22/SUMB[18][52] ) );
  FA_X1 \mult_22/S2_18_51  ( .A(\mult_22/ab[18][51] ), .B(
        \mult_22/CARRYB[17][51] ), .CI(\mult_22/SUMB[17][52] ), .CO(
        \mult_22/CARRYB[18][51] ), .S(\mult_22/SUMB[18][51] ) );
  FA_X1 \mult_22/S2_18_50  ( .A(\mult_22/ab[18][50] ), .B(
        \mult_22/CARRYB[17][50] ), .CI(\mult_22/SUMB[17][51] ), .CO(
        \mult_22/CARRYB[18][50] ), .S(\mult_22/SUMB[18][50] ) );
  FA_X1 \mult_22/S2_18_49  ( .A(\mult_22/ab[18][49] ), .B(
        \mult_22/CARRYB[17][49] ), .CI(\mult_22/SUMB[17][50] ), .CO(
        \mult_22/CARRYB[18][49] ), .S(\mult_22/SUMB[18][49] ) );
  FA_X1 \mult_22/S2_18_48  ( .A(\mult_22/CARRYB[17][48] ), .B(
        \mult_22/ab[18][48] ), .CI(\mult_22/SUMB[17][49] ), .CO(
        \mult_22/CARRYB[18][48] ), .S(\mult_22/SUMB[18][48] ) );
  FA_X1 \mult_22/S2_18_47  ( .A(\mult_22/CARRYB[17][47] ), .B(
        \mult_22/ab[18][47] ), .CI(\mult_22/SUMB[17][48] ), .CO(
        \mult_22/CARRYB[18][47] ), .S(\mult_22/SUMB[18][47] ) );
  FA_X1 \mult_22/S2_18_44  ( .A(\mult_22/ab[18][44] ), .B(
        \mult_22/CARRYB[17][44] ), .CI(\mult_22/SUMB[17][45] ), .CO(
        \mult_22/CARRYB[18][44] ), .S(\mult_22/SUMB[18][44] ) );
  FA_X1 \mult_22/S2_18_41  ( .A(\mult_22/ab[18][41] ), .B(
        \mult_22/CARRYB[17][41] ), .CI(\mult_22/SUMB[17][42] ), .CO(
        \mult_22/CARRYB[18][41] ), .S(\mult_22/SUMB[18][41] ) );
  FA_X1 \mult_22/S2_18_39  ( .A(\mult_22/ab[18][39] ), .B(
        \mult_22/CARRYB[17][39] ), .CI(\mult_22/SUMB[17][40] ), .CO(
        \mult_22/CARRYB[18][39] ), .S(\mult_22/SUMB[18][39] ) );
  FA_X1 \mult_22/S2_18_38  ( .A(\mult_22/ab[18][38] ), .B(
        \mult_22/CARRYB[17][38] ), .CI(\mult_22/SUMB[17][39] ), .CO(
        \mult_22/CARRYB[18][38] ), .S(\mult_22/SUMB[18][38] ) );
  FA_X1 \mult_22/S2_18_37  ( .A(\mult_22/ab[18][37] ), .B(
        \mult_22/CARRYB[17][37] ), .CI(\mult_22/SUMB[17][38] ), .CO(
        \mult_22/CARRYB[18][37] ), .S(\mult_22/SUMB[18][37] ) );
  FA_X1 \mult_22/S2_18_36  ( .A(\mult_22/ab[18][36] ), .B(
        \mult_22/CARRYB[17][36] ), .CI(\mult_22/SUMB[17][37] ), .CO(
        \mult_22/CARRYB[18][36] ), .S(\mult_22/SUMB[18][36] ) );
  FA_X1 \mult_22/S2_18_35  ( .A(\mult_22/ab[18][35] ), .B(
        \mult_22/CARRYB[17][35] ), .CI(\mult_22/SUMB[17][36] ), .CO(
        \mult_22/CARRYB[18][35] ), .S(\mult_22/SUMB[18][35] ) );
  FA_X1 \mult_22/S2_18_34  ( .A(\mult_22/ab[18][34] ), .B(
        \mult_22/CARRYB[17][34] ), .CI(\mult_22/SUMB[17][35] ), .CO(
        \mult_22/CARRYB[18][34] ), .S(\mult_22/SUMB[18][34] ) );
  FA_X1 \mult_22/S2_18_33  ( .A(\mult_22/ab[18][33] ), .B(
        \mult_22/CARRYB[17][33] ), .CI(\mult_22/SUMB[17][34] ), .CO(
        \mult_22/CARRYB[18][33] ), .S(\mult_22/SUMB[18][33] ) );
  FA_X1 \mult_22/S2_18_32  ( .A(\mult_22/ab[18][32] ), .B(
        \mult_22/CARRYB[17][32] ), .CI(\mult_22/SUMB[17][33] ), .CO(
        \mult_22/CARRYB[18][32] ), .S(\mult_22/SUMB[18][32] ) );
  FA_X1 \mult_22/S2_18_31  ( .A(\mult_22/ab[18][31] ), .B(
        \mult_22/CARRYB[17][31] ), .CI(\mult_22/SUMB[17][32] ), .CO(
        \mult_22/CARRYB[18][31] ), .S(\mult_22/SUMB[18][31] ) );
  FA_X1 \mult_22/S2_18_30  ( .A(\mult_22/ab[18][30] ), .B(
        \mult_22/CARRYB[17][30] ), .CI(\mult_22/SUMB[17][31] ), .CO(
        \mult_22/CARRYB[18][30] ), .S(\mult_22/SUMB[18][30] ) );
  FA_X1 \mult_22/S2_18_29  ( .A(\mult_22/ab[18][29] ), .B(
        \mult_22/CARRYB[17][29] ), .CI(\mult_22/SUMB[17][30] ), .CO(
        \mult_22/CARRYB[18][29] ), .S(\mult_22/SUMB[18][29] ) );
  FA_X1 \mult_22/S2_18_28  ( .A(\mult_22/ab[18][28] ), .B(
        \mult_22/CARRYB[17][28] ), .CI(\mult_22/SUMB[17][29] ), .CO(
        \mult_22/CARRYB[18][28] ), .S(\mult_22/SUMB[18][28] ) );
  FA_X1 \mult_22/S2_18_27  ( .A(\mult_22/ab[18][27] ), .B(
        \mult_22/CARRYB[17][27] ), .CI(\mult_22/SUMB[17][28] ), .CO(
        \mult_22/CARRYB[18][27] ), .S(\mult_22/SUMB[18][27] ) );
  FA_X1 \mult_22/S2_18_26  ( .A(\mult_22/ab[18][26] ), .B(
        \mult_22/CARRYB[17][26] ), .CI(\mult_22/SUMB[17][27] ), .CO(
        \mult_22/CARRYB[18][26] ), .S(\mult_22/SUMB[18][26] ) );
  FA_X1 \mult_22/S2_18_25  ( .A(\mult_22/ab[18][25] ), .B(
        \mult_22/CARRYB[17][25] ), .CI(\mult_22/SUMB[17][26] ), .CO(
        \mult_22/CARRYB[18][25] ), .S(\mult_22/SUMB[18][25] ) );
  FA_X1 \mult_22/S2_18_24  ( .A(\mult_22/ab[18][24] ), .B(
        \mult_22/CARRYB[17][24] ), .CI(\mult_22/SUMB[17][25] ), .CO(
        \mult_22/CARRYB[18][24] ), .S(\mult_22/SUMB[18][24] ) );
  FA_X1 \mult_22/S2_18_23  ( .A(\mult_22/ab[18][23] ), .B(
        \mult_22/CARRYB[17][23] ), .CI(\mult_22/SUMB[17][24] ), .CO(
        \mult_22/CARRYB[18][23] ), .S(\mult_22/SUMB[18][23] ) );
  FA_X1 \mult_22/S2_18_22  ( .A(\mult_22/ab[18][22] ), .B(
        \mult_22/CARRYB[17][22] ), .CI(\mult_22/SUMB[17][23] ), .CO(
        \mult_22/CARRYB[18][22] ), .S(\mult_22/SUMB[18][22] ) );
  FA_X1 \mult_22/S2_18_21  ( .A(\mult_22/ab[18][21] ), .B(
        \mult_22/CARRYB[17][21] ), .CI(\mult_22/SUMB[17][22] ), .CO(
        \mult_22/CARRYB[18][21] ), .S(\mult_22/SUMB[18][21] ) );
  FA_X1 \mult_22/S2_18_20  ( .A(\mult_22/ab[18][20] ), .B(
        \mult_22/CARRYB[17][20] ), .CI(\mult_22/SUMB[17][21] ), .CO(
        \mult_22/CARRYB[18][20] ), .S(\mult_22/SUMB[18][20] ) );
  FA_X1 \mult_22/S2_18_19  ( .A(\mult_22/ab[18][19] ), .B(
        \mult_22/CARRYB[17][19] ), .CI(\mult_22/SUMB[17][20] ), .CO(
        \mult_22/CARRYB[18][19] ), .S(\mult_22/SUMB[18][19] ) );
  FA_X1 \mult_22/S2_18_18  ( .A(\mult_22/ab[18][18] ), .B(
        \mult_22/CARRYB[17][18] ), .CI(\mult_22/SUMB[17][19] ), .CO(
        \mult_22/CARRYB[18][18] ), .S(\mult_22/SUMB[18][18] ) );
  FA_X1 \mult_22/S2_18_17  ( .A(\mult_22/ab[18][17] ), .B(
        \mult_22/CARRYB[17][17] ), .CI(\mult_22/SUMB[17][18] ), .CO(
        \mult_22/CARRYB[18][17] ), .S(\mult_22/SUMB[18][17] ) );
  FA_X1 \mult_22/S2_18_16  ( .A(\mult_22/ab[18][16] ), .B(
        \mult_22/CARRYB[17][16] ), .CI(\mult_22/SUMB[17][17] ), .CO(
        \mult_22/CARRYB[18][16] ), .S(\mult_22/SUMB[18][16] ) );
  FA_X1 \mult_22/S2_18_15  ( .A(\mult_22/ab[18][15] ), .B(
        \mult_22/CARRYB[17][15] ), .CI(\mult_22/SUMB[17][16] ), .CO(
        \mult_22/CARRYB[18][15] ), .S(\mult_22/SUMB[18][15] ) );
  FA_X1 \mult_22/S2_18_14  ( .A(\mult_22/ab[18][14] ), .B(
        \mult_22/CARRYB[17][14] ), .CI(\mult_22/SUMB[17][15] ), .CO(
        \mult_22/CARRYB[18][14] ), .S(\mult_22/SUMB[18][14] ) );
  FA_X1 \mult_22/S2_18_13  ( .A(\mult_22/ab[18][13] ), .B(
        \mult_22/CARRYB[17][13] ), .CI(\mult_22/SUMB[17][14] ), .CO(
        \mult_22/CARRYB[18][13] ), .S(\mult_22/SUMB[18][13] ) );
  FA_X1 \mult_22/S2_18_12  ( .A(\mult_22/ab[18][12] ), .B(
        \mult_22/CARRYB[17][12] ), .CI(\mult_22/SUMB[17][13] ), .CO(
        \mult_22/CARRYB[18][12] ), .S(\mult_22/SUMB[18][12] ) );
  FA_X1 \mult_22/S2_18_11  ( .A(\mult_22/ab[18][11] ), .B(
        \mult_22/CARRYB[17][11] ), .CI(\mult_22/SUMB[17][12] ), .CO(
        \mult_22/CARRYB[18][11] ), .S(\mult_22/SUMB[18][11] ) );
  FA_X1 \mult_22/S2_18_10  ( .A(\mult_22/ab[18][10] ), .B(
        \mult_22/CARRYB[17][10] ), .CI(\mult_22/SUMB[17][11] ), .CO(
        \mult_22/CARRYB[18][10] ), .S(\mult_22/SUMB[18][10] ) );
  FA_X1 \mult_22/S2_18_9  ( .A(\mult_22/ab[18][9] ), .B(
        \mult_22/CARRYB[17][9] ), .CI(\mult_22/SUMB[17][10] ), .CO(
        \mult_22/CARRYB[18][9] ), .S(\mult_22/SUMB[18][9] ) );
  FA_X1 \mult_22/S2_18_8  ( .A(\mult_22/ab[18][8] ), .B(
        \mult_22/CARRYB[17][8] ), .CI(\mult_22/SUMB[17][9] ), .CO(
        \mult_22/CARRYB[18][8] ), .S(\mult_22/SUMB[18][8] ) );
  FA_X1 \mult_22/S2_18_7  ( .A(\mult_22/ab[18][7] ), .B(
        \mult_22/CARRYB[17][7] ), .CI(\mult_22/SUMB[17][8] ), .CO(
        \mult_22/CARRYB[18][7] ), .S(\mult_22/SUMB[18][7] ) );
  FA_X1 \mult_22/S2_18_6  ( .A(\mult_22/ab[18][6] ), .B(
        \mult_22/CARRYB[17][6] ), .CI(\mult_22/SUMB[17][7] ), .CO(
        \mult_22/CARRYB[18][6] ), .S(\mult_22/SUMB[18][6] ) );
  FA_X1 \mult_22/S2_18_5  ( .A(\mult_22/ab[18][5] ), .B(
        \mult_22/CARRYB[17][5] ), .CI(\mult_22/SUMB[17][6] ), .CO(
        \mult_22/CARRYB[18][5] ), .S(\mult_22/SUMB[18][5] ) );
  FA_X1 \mult_22/S2_18_4  ( .A(\mult_22/ab[18][4] ), .B(
        \mult_22/CARRYB[17][4] ), .CI(\mult_22/SUMB[17][5] ), .CO(
        \mult_22/CARRYB[18][4] ), .S(\mult_22/SUMB[18][4] ) );
  FA_X1 \mult_22/S2_18_3  ( .A(\mult_22/ab[18][3] ), .B(
        \mult_22/CARRYB[17][3] ), .CI(\mult_22/SUMB[17][4] ), .CO(
        \mult_22/CARRYB[18][3] ), .S(\mult_22/SUMB[18][3] ) );
  FA_X1 \mult_22/S2_18_2  ( .A(\mult_22/ab[18][2] ), .B(
        \mult_22/CARRYB[17][2] ), .CI(\mult_22/SUMB[17][3] ), .CO(
        \mult_22/CARRYB[18][2] ), .S(\mult_22/SUMB[18][2] ) );
  FA_X1 \mult_22/S2_18_1  ( .A(\mult_22/ab[18][1] ), .B(
        \mult_22/CARRYB[17][1] ), .CI(\mult_22/SUMB[17][2] ), .CO(
        \mult_22/CARRYB[18][1] ), .S(\mult_22/SUMB[18][1] ) );
  FA_X1 \mult_22/S1_18_0  ( .A(\mult_22/ab[18][0] ), .B(
        \mult_22/CARRYB[17][0] ), .CI(\mult_22/SUMB[17][1] ), .CO(
        \mult_22/CARRYB[18][0] ), .S(N146) );
  FA_X1 \mult_22/S3_19_62  ( .A(\mult_22/ab[19][62] ), .B(
        \mult_22/CARRYB[18][62] ), .CI(\mult_22/ab[18][63] ), .CO(
        \mult_22/CARRYB[19][62] ), .S(\mult_22/SUMB[19][62] ) );
  FA_X1 \mult_22/S2_19_61  ( .A(\mult_22/ab[19][61] ), .B(
        \mult_22/CARRYB[18][61] ), .CI(\mult_22/SUMB[18][62] ), .CO(
        \mult_22/CARRYB[19][61] ), .S(\mult_22/SUMB[19][61] ) );
  FA_X1 \mult_22/S2_19_60  ( .A(\mult_22/ab[19][60] ), .B(
        \mult_22/CARRYB[18][60] ), .CI(\mult_22/SUMB[18][61] ), .CO(
        \mult_22/CARRYB[19][60] ), .S(\mult_22/SUMB[19][60] ) );
  FA_X1 \mult_22/S2_19_59  ( .A(\mult_22/ab[19][59] ), .B(
        \mult_22/CARRYB[18][59] ), .CI(\mult_22/SUMB[18][60] ), .CO(
        \mult_22/CARRYB[19][59] ), .S(\mult_22/SUMB[19][59] ) );
  FA_X1 \mult_22/S2_19_58  ( .A(\mult_22/ab[19][58] ), .B(
        \mult_22/CARRYB[18][58] ), .CI(\mult_22/SUMB[18][59] ), .CO(
        \mult_22/CARRYB[19][58] ), .S(\mult_22/SUMB[19][58] ) );
  FA_X1 \mult_22/S2_19_57  ( .A(\mult_22/ab[19][57] ), .B(
        \mult_22/CARRYB[18][57] ), .CI(\mult_22/SUMB[18][58] ), .CO(
        \mult_22/CARRYB[19][57] ), .S(\mult_22/SUMB[19][57] ) );
  FA_X1 \mult_22/S2_19_56  ( .A(\mult_22/ab[19][56] ), .B(
        \mult_22/CARRYB[18][56] ), .CI(\mult_22/SUMB[18][57] ), .CO(
        \mult_22/CARRYB[19][56] ), .S(\mult_22/SUMB[19][56] ) );
  FA_X1 \mult_22/S2_19_55  ( .A(\mult_22/ab[19][55] ), .B(
        \mult_22/CARRYB[18][55] ), .CI(\mult_22/SUMB[18][56] ), .CO(
        \mult_22/CARRYB[19][55] ), .S(\mult_22/SUMB[19][55] ) );
  FA_X1 \mult_22/S2_19_54  ( .A(\mult_22/ab[19][54] ), .B(
        \mult_22/CARRYB[18][54] ), .CI(\mult_22/SUMB[18][55] ), .CO(
        \mult_22/CARRYB[19][54] ), .S(\mult_22/SUMB[19][54] ) );
  FA_X1 \mult_22/S2_19_53  ( .A(\mult_22/ab[19][53] ), .B(
        \mult_22/CARRYB[18][53] ), .CI(\mult_22/SUMB[18][54] ), .CO(
        \mult_22/CARRYB[19][53] ), .S(\mult_22/SUMB[19][53] ) );
  FA_X1 \mult_22/S2_19_52  ( .A(\mult_22/ab[19][52] ), .B(
        \mult_22/CARRYB[18][52] ), .CI(\mult_22/SUMB[18][53] ), .CO(
        \mult_22/CARRYB[19][52] ), .S(\mult_22/SUMB[19][52] ) );
  FA_X1 \mult_22/S2_19_51  ( .A(\mult_22/ab[19][51] ), .B(
        \mult_22/CARRYB[18][51] ), .CI(\mult_22/SUMB[18][52] ), .CO(
        \mult_22/CARRYB[19][51] ), .S(\mult_22/SUMB[19][51] ) );
  FA_X1 \mult_22/S2_19_50  ( .A(\mult_22/ab[19][50] ), .B(
        \mult_22/CARRYB[18][50] ), .CI(\mult_22/SUMB[18][51] ), .CO(
        \mult_22/CARRYB[19][50] ), .S(\mult_22/SUMB[19][50] ) );
  FA_X1 \mult_22/S2_19_49  ( .A(\mult_22/ab[19][49] ), .B(
        \mult_22/CARRYB[18][49] ), .CI(\mult_22/SUMB[18][50] ), .CO(
        \mult_22/CARRYB[19][49] ), .S(\mult_22/SUMB[19][49] ) );
  FA_X1 \mult_22/S2_19_48  ( .A(\mult_22/CARRYB[18][48] ), .B(
        \mult_22/ab[19][48] ), .CI(\mult_22/SUMB[18][49] ), .CO(
        \mult_22/CARRYB[19][48] ), .S(\mult_22/SUMB[19][48] ) );
  FA_X1 \mult_22/S2_19_47  ( .A(\mult_22/ab[19][47] ), .B(
        \mult_22/CARRYB[18][47] ), .CI(\mult_22/SUMB[18][48] ), .CO(
        \mult_22/CARRYB[19][47] ), .S(\mult_22/SUMB[19][47] ) );
  FA_X1 \mult_22/S2_19_46  ( .A(\mult_22/ab[19][46] ), .B(
        \mult_22/CARRYB[18][46] ), .CI(\mult_22/SUMB[18][47] ), .CO(
        \mult_22/CARRYB[19][46] ), .S(\mult_22/SUMB[19][46] ) );
  FA_X1 \mult_22/S2_19_44  ( .A(\mult_22/ab[19][44] ), .B(
        \mult_22/CARRYB[18][44] ), .CI(\mult_22/SUMB[18][45] ), .CO(
        \mult_22/CARRYB[19][44] ), .S(\mult_22/SUMB[19][44] ) );
  FA_X1 \mult_22/S2_19_43  ( .A(\mult_22/ab[19][43] ), .B(
        \mult_22/CARRYB[18][43] ), .CI(\mult_22/SUMB[18][44] ), .CO(
        \mult_22/CARRYB[19][43] ), .S(\mult_22/SUMB[19][43] ) );
  FA_X1 \mult_22/S2_19_40  ( .A(\mult_22/SUMB[18][41] ), .B(
        \mult_22/ab[19][40] ), .CI(\mult_22/CARRYB[18][40] ), .CO(
        \mult_22/CARRYB[19][40] ), .S(\mult_22/SUMB[19][40] ) );
  FA_X1 \mult_22/S2_19_39  ( .A(\mult_22/ab[19][39] ), .B(
        \mult_22/CARRYB[18][39] ), .CI(\mult_22/SUMB[18][40] ), .CO(
        \mult_22/CARRYB[19][39] ), .S(\mult_22/SUMB[19][39] ) );
  FA_X1 \mult_22/S2_19_38  ( .A(\mult_22/ab[19][38] ), .B(
        \mult_22/CARRYB[18][38] ), .CI(\mult_22/SUMB[18][39] ), .CO(
        \mult_22/CARRYB[19][38] ), .S(\mult_22/SUMB[19][38] ) );
  FA_X1 \mult_22/S2_19_37  ( .A(\mult_22/ab[19][37] ), .B(
        \mult_22/CARRYB[18][37] ), .CI(\mult_22/SUMB[18][38] ), .CO(
        \mult_22/CARRYB[19][37] ), .S(\mult_22/SUMB[19][37] ) );
  FA_X1 \mult_22/S2_19_36  ( .A(\mult_22/ab[19][36] ), .B(
        \mult_22/CARRYB[18][36] ), .CI(\mult_22/SUMB[18][37] ), .CO(
        \mult_22/CARRYB[19][36] ), .S(\mult_22/SUMB[19][36] ) );
  FA_X1 \mult_22/S2_19_35  ( .A(\mult_22/ab[19][35] ), .B(
        \mult_22/CARRYB[18][35] ), .CI(\mult_22/SUMB[18][36] ), .CO(
        \mult_22/CARRYB[19][35] ), .S(\mult_22/SUMB[19][35] ) );
  FA_X1 \mult_22/S2_19_34  ( .A(\mult_22/ab[19][34] ), .B(
        \mult_22/CARRYB[18][34] ), .CI(\mult_22/SUMB[18][35] ), .CO(
        \mult_22/CARRYB[19][34] ), .S(\mult_22/SUMB[19][34] ) );
  FA_X1 \mult_22/S2_19_33  ( .A(\mult_22/ab[19][33] ), .B(
        \mult_22/CARRYB[18][33] ), .CI(\mult_22/SUMB[18][34] ), .CO(
        \mult_22/CARRYB[19][33] ), .S(\mult_22/SUMB[19][33] ) );
  FA_X1 \mult_22/S2_19_32  ( .A(\mult_22/ab[19][32] ), .B(
        \mult_22/CARRYB[18][32] ), .CI(\mult_22/SUMB[18][33] ), .CO(
        \mult_22/CARRYB[19][32] ), .S(\mult_22/SUMB[19][32] ) );
  FA_X1 \mult_22/S2_19_31  ( .A(\mult_22/ab[19][31] ), .B(
        \mult_22/CARRYB[18][31] ), .CI(\mult_22/SUMB[18][32] ), .CO(
        \mult_22/CARRYB[19][31] ), .S(\mult_22/SUMB[19][31] ) );
  FA_X1 \mult_22/S2_19_30  ( .A(\mult_22/ab[19][30] ), .B(
        \mult_22/CARRYB[18][30] ), .CI(\mult_22/SUMB[18][31] ), .CO(
        \mult_22/CARRYB[19][30] ), .S(\mult_22/SUMB[19][30] ) );
  FA_X1 \mult_22/S2_19_29  ( .A(\mult_22/ab[19][29] ), .B(
        \mult_22/CARRYB[18][29] ), .CI(\mult_22/SUMB[18][30] ), .CO(
        \mult_22/CARRYB[19][29] ), .S(\mult_22/SUMB[19][29] ) );
  FA_X1 \mult_22/S2_19_28  ( .A(\mult_22/ab[19][28] ), .B(
        \mult_22/CARRYB[18][28] ), .CI(\mult_22/SUMB[18][29] ), .CO(
        \mult_22/CARRYB[19][28] ), .S(\mult_22/SUMB[19][28] ) );
  FA_X1 \mult_22/S2_19_27  ( .A(\mult_22/ab[19][27] ), .B(
        \mult_22/CARRYB[18][27] ), .CI(\mult_22/SUMB[18][28] ), .CO(
        \mult_22/CARRYB[19][27] ), .S(\mult_22/SUMB[19][27] ) );
  FA_X1 \mult_22/S2_19_26  ( .A(\mult_22/ab[19][26] ), .B(
        \mult_22/CARRYB[18][26] ), .CI(\mult_22/SUMB[18][27] ), .CO(
        \mult_22/CARRYB[19][26] ), .S(\mult_22/SUMB[19][26] ) );
  FA_X1 \mult_22/S2_19_25  ( .A(\mult_22/ab[19][25] ), .B(
        \mult_22/CARRYB[18][25] ), .CI(\mult_22/SUMB[18][26] ), .CO(
        \mult_22/CARRYB[19][25] ), .S(\mult_22/SUMB[19][25] ) );
  FA_X1 \mult_22/S2_19_24  ( .A(\mult_22/ab[19][24] ), .B(
        \mult_22/CARRYB[18][24] ), .CI(\mult_22/SUMB[18][25] ), .CO(
        \mult_22/CARRYB[19][24] ), .S(\mult_22/SUMB[19][24] ) );
  FA_X1 \mult_22/S2_19_23  ( .A(\mult_22/ab[19][23] ), .B(
        \mult_22/CARRYB[18][23] ), .CI(\mult_22/SUMB[18][24] ), .CO(
        \mult_22/CARRYB[19][23] ), .S(\mult_22/SUMB[19][23] ) );
  FA_X1 \mult_22/S2_19_22  ( .A(\mult_22/ab[19][22] ), .B(
        \mult_22/CARRYB[18][22] ), .CI(\mult_22/SUMB[18][23] ), .CO(
        \mult_22/CARRYB[19][22] ), .S(\mult_22/SUMB[19][22] ) );
  FA_X1 \mult_22/S2_19_21  ( .A(\mult_22/ab[19][21] ), .B(
        \mult_22/CARRYB[18][21] ), .CI(\mult_22/SUMB[18][22] ), .CO(
        \mult_22/CARRYB[19][21] ), .S(\mult_22/SUMB[19][21] ) );
  FA_X1 \mult_22/S2_19_20  ( .A(\mult_22/ab[19][20] ), .B(
        \mult_22/CARRYB[18][20] ), .CI(\mult_22/SUMB[18][21] ), .CO(
        \mult_22/CARRYB[19][20] ), .S(\mult_22/SUMB[19][20] ) );
  FA_X1 \mult_22/S2_19_19  ( .A(\mult_22/ab[19][19] ), .B(
        \mult_22/CARRYB[18][19] ), .CI(\mult_22/SUMB[18][20] ), .CO(
        \mult_22/CARRYB[19][19] ), .S(\mult_22/SUMB[19][19] ) );
  FA_X1 \mult_22/S2_19_18  ( .A(\mult_22/ab[19][18] ), .B(
        \mult_22/CARRYB[18][18] ), .CI(\mult_22/SUMB[18][19] ), .CO(
        \mult_22/CARRYB[19][18] ), .S(\mult_22/SUMB[19][18] ) );
  FA_X1 \mult_22/S2_19_17  ( .A(\mult_22/ab[19][17] ), .B(
        \mult_22/CARRYB[18][17] ), .CI(\mult_22/SUMB[18][18] ), .CO(
        \mult_22/CARRYB[19][17] ), .S(\mult_22/SUMB[19][17] ) );
  FA_X1 \mult_22/S2_19_16  ( .A(\mult_22/ab[19][16] ), .B(
        \mult_22/CARRYB[18][16] ), .CI(\mult_22/SUMB[18][17] ), .CO(
        \mult_22/CARRYB[19][16] ), .S(\mult_22/SUMB[19][16] ) );
  FA_X1 \mult_22/S2_19_15  ( .A(\mult_22/ab[19][15] ), .B(
        \mult_22/CARRYB[18][15] ), .CI(\mult_22/SUMB[18][16] ), .CO(
        \mult_22/CARRYB[19][15] ), .S(\mult_22/SUMB[19][15] ) );
  FA_X1 \mult_22/S2_19_14  ( .A(\mult_22/ab[19][14] ), .B(
        \mult_22/CARRYB[18][14] ), .CI(\mult_22/SUMB[18][15] ), .CO(
        \mult_22/CARRYB[19][14] ), .S(\mult_22/SUMB[19][14] ) );
  FA_X1 \mult_22/S2_19_13  ( .A(\mult_22/ab[19][13] ), .B(
        \mult_22/CARRYB[18][13] ), .CI(\mult_22/SUMB[18][14] ), .CO(
        \mult_22/CARRYB[19][13] ), .S(\mult_22/SUMB[19][13] ) );
  FA_X1 \mult_22/S2_19_12  ( .A(\mult_22/ab[19][12] ), .B(
        \mult_22/CARRYB[18][12] ), .CI(\mult_22/SUMB[18][13] ), .CO(
        \mult_22/CARRYB[19][12] ), .S(\mult_22/SUMB[19][12] ) );
  FA_X1 \mult_22/S2_19_11  ( .A(\mult_22/ab[19][11] ), .B(
        \mult_22/CARRYB[18][11] ), .CI(\mult_22/SUMB[18][12] ), .CO(
        \mult_22/CARRYB[19][11] ), .S(\mult_22/SUMB[19][11] ) );
  FA_X1 \mult_22/S2_19_10  ( .A(\mult_22/ab[19][10] ), .B(
        \mult_22/CARRYB[18][10] ), .CI(\mult_22/SUMB[18][11] ), .CO(
        \mult_22/CARRYB[19][10] ), .S(\mult_22/SUMB[19][10] ) );
  FA_X1 \mult_22/S2_19_9  ( .A(\mult_22/ab[19][9] ), .B(
        \mult_22/CARRYB[18][9] ), .CI(\mult_22/SUMB[18][10] ), .CO(
        \mult_22/CARRYB[19][9] ), .S(\mult_22/SUMB[19][9] ) );
  FA_X1 \mult_22/S2_19_8  ( .A(\mult_22/ab[19][8] ), .B(
        \mult_22/CARRYB[18][8] ), .CI(\mult_22/SUMB[18][9] ), .CO(
        \mult_22/CARRYB[19][8] ), .S(\mult_22/SUMB[19][8] ) );
  FA_X1 \mult_22/S2_19_7  ( .A(\mult_22/ab[19][7] ), .B(
        \mult_22/CARRYB[18][7] ), .CI(\mult_22/SUMB[18][8] ), .CO(
        \mult_22/CARRYB[19][7] ), .S(\mult_22/SUMB[19][7] ) );
  FA_X1 \mult_22/S2_19_6  ( .A(\mult_22/ab[19][6] ), .B(
        \mult_22/CARRYB[18][6] ), .CI(\mult_22/SUMB[18][7] ), .CO(
        \mult_22/CARRYB[19][6] ), .S(\mult_22/SUMB[19][6] ) );
  FA_X1 \mult_22/S2_19_5  ( .A(\mult_22/ab[19][5] ), .B(
        \mult_22/CARRYB[18][5] ), .CI(\mult_22/SUMB[18][6] ), .CO(
        \mult_22/CARRYB[19][5] ), .S(\mult_22/SUMB[19][5] ) );
  FA_X1 \mult_22/S2_19_4  ( .A(\mult_22/ab[19][4] ), .B(
        \mult_22/CARRYB[18][4] ), .CI(\mult_22/SUMB[18][5] ), .CO(
        \mult_22/CARRYB[19][4] ), .S(\mult_22/SUMB[19][4] ) );
  FA_X1 \mult_22/S2_19_3  ( .A(\mult_22/ab[19][3] ), .B(
        \mult_22/CARRYB[18][3] ), .CI(\mult_22/SUMB[18][4] ), .CO(
        \mult_22/CARRYB[19][3] ), .S(\mult_22/SUMB[19][3] ) );
  FA_X1 \mult_22/S2_19_2  ( .A(\mult_22/ab[19][2] ), .B(
        \mult_22/CARRYB[18][2] ), .CI(\mult_22/SUMB[18][3] ), .CO(
        \mult_22/CARRYB[19][2] ), .S(\mult_22/SUMB[19][2] ) );
  FA_X1 \mult_22/S2_19_1  ( .A(\mult_22/ab[19][1] ), .B(
        \mult_22/CARRYB[18][1] ), .CI(\mult_22/SUMB[18][2] ), .CO(
        \mult_22/CARRYB[19][1] ), .S(\mult_22/SUMB[19][1] ) );
  FA_X1 \mult_22/S1_19_0  ( .A(\mult_22/ab[19][0] ), .B(
        \mult_22/CARRYB[18][0] ), .CI(\mult_22/SUMB[18][1] ), .CO(
        \mult_22/CARRYB[19][0] ), .S(N147) );
  FA_X1 \mult_22/S3_20_62  ( .A(\mult_22/ab[20][62] ), .B(
        \mult_22/CARRYB[19][62] ), .CI(\mult_22/ab[19][63] ), .CO(
        \mult_22/CARRYB[20][62] ), .S(\mult_22/SUMB[20][62] ) );
  FA_X1 \mult_22/S2_20_61  ( .A(\mult_22/ab[20][61] ), .B(
        \mult_22/CARRYB[19][61] ), .CI(\mult_22/SUMB[19][62] ), .CO(
        \mult_22/CARRYB[20][61] ), .S(\mult_22/SUMB[20][61] ) );
  FA_X1 \mult_22/S2_20_60  ( .A(\mult_22/ab[20][60] ), .B(
        \mult_22/CARRYB[19][60] ), .CI(\mult_22/SUMB[19][61] ), .CO(
        \mult_22/CARRYB[20][60] ), .S(\mult_22/SUMB[20][60] ) );
  FA_X1 \mult_22/S2_20_59  ( .A(\mult_22/ab[20][59] ), .B(
        \mult_22/CARRYB[19][59] ), .CI(\mult_22/SUMB[19][60] ), .CO(
        \mult_22/CARRYB[20][59] ), .S(\mult_22/SUMB[20][59] ) );
  FA_X1 \mult_22/S2_20_58  ( .A(\mult_22/ab[20][58] ), .B(
        \mult_22/CARRYB[19][58] ), .CI(\mult_22/SUMB[19][59] ), .CO(
        \mult_22/CARRYB[20][58] ), .S(\mult_22/SUMB[20][58] ) );
  FA_X1 \mult_22/S2_20_57  ( .A(\mult_22/ab[20][57] ), .B(
        \mult_22/CARRYB[19][57] ), .CI(\mult_22/SUMB[19][58] ), .CO(
        \mult_22/CARRYB[20][57] ), .S(\mult_22/SUMB[20][57] ) );
  FA_X1 \mult_22/S2_20_56  ( .A(\mult_22/ab[20][56] ), .B(
        \mult_22/CARRYB[19][56] ), .CI(\mult_22/SUMB[19][57] ), .CO(
        \mult_22/CARRYB[20][56] ), .S(\mult_22/SUMB[20][56] ) );
  FA_X1 \mult_22/S2_20_55  ( .A(\mult_22/ab[20][55] ), .B(
        \mult_22/CARRYB[19][55] ), .CI(\mult_22/SUMB[19][56] ), .CO(
        \mult_22/CARRYB[20][55] ), .S(\mult_22/SUMB[20][55] ) );
  FA_X1 \mult_22/S2_20_54  ( .A(\mult_22/ab[20][54] ), .B(
        \mult_22/CARRYB[19][54] ), .CI(\mult_22/SUMB[19][55] ), .CO(
        \mult_22/CARRYB[20][54] ), .S(\mult_22/SUMB[20][54] ) );
  FA_X1 \mult_22/S2_20_53  ( .A(\mult_22/ab[20][53] ), .B(
        \mult_22/CARRYB[19][53] ), .CI(\mult_22/SUMB[19][54] ), .CO(
        \mult_22/CARRYB[20][53] ), .S(\mult_22/SUMB[20][53] ) );
  FA_X1 \mult_22/S2_20_52  ( .A(\mult_22/ab[20][52] ), .B(
        \mult_22/CARRYB[19][52] ), .CI(\mult_22/SUMB[19][53] ), .CO(
        \mult_22/CARRYB[20][52] ), .S(\mult_22/SUMB[20][52] ) );
  FA_X1 \mult_22/S2_20_51  ( .A(\mult_22/ab[20][51] ), .B(
        \mult_22/CARRYB[19][51] ), .CI(\mult_22/SUMB[19][52] ), .CO(
        \mult_22/CARRYB[20][51] ), .S(\mult_22/SUMB[20][51] ) );
  FA_X1 \mult_22/S2_20_50  ( .A(\mult_22/ab[20][50] ), .B(
        \mult_22/CARRYB[19][50] ), .CI(\mult_22/SUMB[19][51] ), .CO(
        \mult_22/CARRYB[20][50] ), .S(\mult_22/SUMB[20][50] ) );
  FA_X1 \mult_22/S2_20_49  ( .A(\mult_22/ab[20][49] ), .B(
        \mult_22/CARRYB[19][49] ), .CI(\mult_22/SUMB[19][50] ), .CO(
        \mult_22/CARRYB[20][49] ), .S(\mult_22/SUMB[20][49] ) );
  FA_X1 \mult_22/S2_20_48  ( .A(\mult_22/ab[20][48] ), .B(
        \mult_22/CARRYB[19][48] ), .CI(\mult_22/SUMB[19][49] ), .CO(
        \mult_22/CARRYB[20][48] ), .S(\mult_22/SUMB[20][48] ) );
  FA_X1 \mult_22/S2_20_47  ( .A(\mult_22/ab[20][47] ), .B(
        \mult_22/CARRYB[19][47] ), .CI(\mult_22/SUMB[19][48] ), .CO(
        \mult_22/CARRYB[20][47] ), .S(\mult_22/SUMB[20][47] ) );
  FA_X1 \mult_22/S2_20_46  ( .A(\mult_22/CARRYB[19][46] ), .B(
        \mult_22/ab[20][46] ), .CI(\mult_22/SUMB[19][47] ), .CO(
        \mult_22/CARRYB[20][46] ), .S(\mult_22/SUMB[20][46] ) );
  FA_X1 \mult_22/S2_20_45  ( .A(\mult_22/ab[20][45] ), .B(
        \mult_22/CARRYB[19][45] ), .CI(\mult_22/SUMB[19][46] ), .CO(
        \mult_22/CARRYB[20][45] ), .S(\mult_22/SUMB[20][45] ) );
  FA_X1 \mult_22/S2_20_43  ( .A(\mult_22/CARRYB[19][43] ), .B(
        \mult_22/ab[20][43] ), .CI(\mult_22/SUMB[19][44] ), .CO(
        \mult_22/CARRYB[20][43] ), .S(\mult_22/SUMB[20][43] ) );
  FA_X1 \mult_22/S2_20_42  ( .A(\mult_22/ab[20][42] ), .B(
        \mult_22/CARRYB[19][42] ), .CI(\mult_22/SUMB[19][43] ), .CO(
        \mult_22/CARRYB[20][42] ), .S(\mult_22/SUMB[20][42] ) );
  FA_X1 \mult_22/S2_20_41  ( .A(\mult_22/ab[20][41] ), .B(
        \mult_22/CARRYB[19][41] ), .CI(\mult_22/SUMB[19][42] ), .CO(
        \mult_22/CARRYB[20][41] ), .S(\mult_22/SUMB[20][41] ) );
  FA_X1 \mult_22/S2_20_40  ( .A(\mult_22/ab[20][40] ), .B(
        \mult_22/CARRYB[19][40] ), .CI(\mult_22/SUMB[19][41] ), .CO(
        \mult_22/CARRYB[20][40] ), .S(\mult_22/SUMB[20][40] ) );
  FA_X1 \mult_22/S2_20_39  ( .A(\mult_22/ab[20][39] ), .B(
        \mult_22/CARRYB[19][39] ), .CI(\mult_22/SUMB[19][40] ), .CO(
        \mult_22/CARRYB[20][39] ), .S(\mult_22/SUMB[20][39] ) );
  FA_X1 \mult_22/S2_20_37  ( .A(\mult_22/ab[20][37] ), .B(
        \mult_22/CARRYB[19][37] ), .CI(\mult_22/SUMB[19][38] ), .CO(
        \mult_22/CARRYB[20][37] ), .S(\mult_22/SUMB[20][37] ) );
  FA_X1 \mult_22/S2_20_36  ( .A(\mult_22/ab[20][36] ), .B(
        \mult_22/CARRYB[19][36] ), .CI(\mult_22/SUMB[19][37] ), .CO(
        \mult_22/CARRYB[20][36] ), .S(\mult_22/SUMB[20][36] ) );
  FA_X1 \mult_22/S2_20_35  ( .A(\mult_22/ab[20][35] ), .B(
        \mult_22/CARRYB[19][35] ), .CI(\mult_22/SUMB[19][36] ), .CO(
        \mult_22/CARRYB[20][35] ), .S(\mult_22/SUMB[20][35] ) );
  FA_X1 \mult_22/S2_20_34  ( .A(\mult_22/ab[20][34] ), .B(
        \mult_22/CARRYB[19][34] ), .CI(\mult_22/SUMB[19][35] ), .CO(
        \mult_22/CARRYB[20][34] ), .S(\mult_22/SUMB[20][34] ) );
  FA_X1 \mult_22/S2_20_33  ( .A(\mult_22/ab[20][33] ), .B(
        \mult_22/CARRYB[19][33] ), .CI(\mult_22/SUMB[19][34] ), .CO(
        \mult_22/CARRYB[20][33] ), .S(\mult_22/SUMB[20][33] ) );
  FA_X1 \mult_22/S2_20_32  ( .A(\mult_22/ab[20][32] ), .B(
        \mult_22/CARRYB[19][32] ), .CI(\mult_22/SUMB[19][33] ), .CO(
        \mult_22/CARRYB[20][32] ), .S(\mult_22/SUMB[20][32] ) );
  FA_X1 \mult_22/S2_20_31  ( .A(\mult_22/ab[20][31] ), .B(
        \mult_22/CARRYB[19][31] ), .CI(\mult_22/SUMB[19][32] ), .CO(
        \mult_22/CARRYB[20][31] ), .S(\mult_22/SUMB[20][31] ) );
  FA_X1 \mult_22/S2_20_30  ( .A(\mult_22/ab[20][30] ), .B(
        \mult_22/CARRYB[19][30] ), .CI(\mult_22/SUMB[19][31] ), .CO(
        \mult_22/CARRYB[20][30] ), .S(\mult_22/SUMB[20][30] ) );
  FA_X1 \mult_22/S2_20_29  ( .A(\mult_22/ab[20][29] ), .B(
        \mult_22/CARRYB[19][29] ), .CI(\mult_22/SUMB[19][30] ), .CO(
        \mult_22/CARRYB[20][29] ), .S(\mult_22/SUMB[20][29] ) );
  FA_X1 \mult_22/S2_20_28  ( .A(\mult_22/ab[20][28] ), .B(
        \mult_22/CARRYB[19][28] ), .CI(\mult_22/SUMB[19][29] ), .CO(
        \mult_22/CARRYB[20][28] ), .S(\mult_22/SUMB[20][28] ) );
  FA_X1 \mult_22/S2_20_27  ( .A(\mult_22/ab[20][27] ), .B(
        \mult_22/CARRYB[19][27] ), .CI(\mult_22/SUMB[19][28] ), .CO(
        \mult_22/CARRYB[20][27] ), .S(\mult_22/SUMB[20][27] ) );
  FA_X1 \mult_22/S2_20_26  ( .A(\mult_22/ab[20][26] ), .B(
        \mult_22/CARRYB[19][26] ), .CI(\mult_22/SUMB[19][27] ), .CO(
        \mult_22/CARRYB[20][26] ), .S(\mult_22/SUMB[20][26] ) );
  FA_X1 \mult_22/S2_20_25  ( .A(\mult_22/ab[20][25] ), .B(
        \mult_22/CARRYB[19][25] ), .CI(\mult_22/SUMB[19][26] ), .CO(
        \mult_22/CARRYB[20][25] ), .S(\mult_22/SUMB[20][25] ) );
  FA_X1 \mult_22/S2_20_24  ( .A(\mult_22/ab[20][24] ), .B(
        \mult_22/CARRYB[19][24] ), .CI(\mult_22/SUMB[19][25] ), .CO(
        \mult_22/CARRYB[20][24] ), .S(\mult_22/SUMB[20][24] ) );
  FA_X1 \mult_22/S2_20_23  ( .A(\mult_22/ab[20][23] ), .B(
        \mult_22/CARRYB[19][23] ), .CI(\mult_22/SUMB[19][24] ), .CO(
        \mult_22/CARRYB[20][23] ), .S(\mult_22/SUMB[20][23] ) );
  FA_X1 \mult_22/S2_20_22  ( .A(\mult_22/ab[20][22] ), .B(
        \mult_22/CARRYB[19][22] ), .CI(\mult_22/SUMB[19][23] ), .CO(
        \mult_22/CARRYB[20][22] ), .S(\mult_22/SUMB[20][22] ) );
  FA_X1 \mult_22/S2_20_21  ( .A(\mult_22/ab[20][21] ), .B(
        \mult_22/CARRYB[19][21] ), .CI(\mult_22/SUMB[19][22] ), .CO(
        \mult_22/CARRYB[20][21] ), .S(\mult_22/SUMB[20][21] ) );
  FA_X1 \mult_22/S2_20_20  ( .A(\mult_22/ab[20][20] ), .B(
        \mult_22/CARRYB[19][20] ), .CI(\mult_22/SUMB[19][21] ), .CO(
        \mult_22/CARRYB[20][20] ), .S(\mult_22/SUMB[20][20] ) );
  FA_X1 \mult_22/S2_20_19  ( .A(\mult_22/ab[20][19] ), .B(
        \mult_22/CARRYB[19][19] ), .CI(\mult_22/SUMB[19][20] ), .CO(
        \mult_22/CARRYB[20][19] ), .S(\mult_22/SUMB[20][19] ) );
  FA_X1 \mult_22/S2_20_18  ( .A(\mult_22/ab[20][18] ), .B(
        \mult_22/CARRYB[19][18] ), .CI(\mult_22/SUMB[19][19] ), .CO(
        \mult_22/CARRYB[20][18] ), .S(\mult_22/SUMB[20][18] ) );
  FA_X1 \mult_22/S2_20_17  ( .A(\mult_22/ab[20][17] ), .B(
        \mult_22/CARRYB[19][17] ), .CI(\mult_22/SUMB[19][18] ), .CO(
        \mult_22/CARRYB[20][17] ), .S(\mult_22/SUMB[20][17] ) );
  FA_X1 \mult_22/S2_20_16  ( .A(\mult_22/ab[20][16] ), .B(
        \mult_22/CARRYB[19][16] ), .CI(\mult_22/SUMB[19][17] ), .CO(
        \mult_22/CARRYB[20][16] ), .S(\mult_22/SUMB[20][16] ) );
  FA_X1 \mult_22/S2_20_15  ( .A(\mult_22/ab[20][15] ), .B(
        \mult_22/CARRYB[19][15] ), .CI(\mult_22/SUMB[19][16] ), .CO(
        \mult_22/CARRYB[20][15] ), .S(\mult_22/SUMB[20][15] ) );
  FA_X1 \mult_22/S2_20_14  ( .A(\mult_22/ab[20][14] ), .B(
        \mult_22/CARRYB[19][14] ), .CI(\mult_22/SUMB[19][15] ), .CO(
        \mult_22/CARRYB[20][14] ), .S(\mult_22/SUMB[20][14] ) );
  FA_X1 \mult_22/S2_20_13  ( .A(\mult_22/ab[20][13] ), .B(
        \mult_22/CARRYB[19][13] ), .CI(\mult_22/SUMB[19][14] ), .CO(
        \mult_22/CARRYB[20][13] ), .S(\mult_22/SUMB[20][13] ) );
  FA_X1 \mult_22/S2_20_12  ( .A(\mult_22/ab[20][12] ), .B(
        \mult_22/CARRYB[19][12] ), .CI(\mult_22/SUMB[19][13] ), .CO(
        \mult_22/CARRYB[20][12] ), .S(\mult_22/SUMB[20][12] ) );
  FA_X1 \mult_22/S2_20_11  ( .A(\mult_22/ab[20][11] ), .B(
        \mult_22/CARRYB[19][11] ), .CI(\mult_22/SUMB[19][12] ), .CO(
        \mult_22/CARRYB[20][11] ), .S(\mult_22/SUMB[20][11] ) );
  FA_X1 \mult_22/S2_20_10  ( .A(\mult_22/ab[20][10] ), .B(
        \mult_22/CARRYB[19][10] ), .CI(\mult_22/SUMB[19][11] ), .CO(
        \mult_22/CARRYB[20][10] ), .S(\mult_22/SUMB[20][10] ) );
  FA_X1 \mult_22/S2_20_9  ( .A(\mult_22/ab[20][9] ), .B(
        \mult_22/CARRYB[19][9] ), .CI(\mult_22/SUMB[19][10] ), .CO(
        \mult_22/CARRYB[20][9] ), .S(\mult_22/SUMB[20][9] ) );
  FA_X1 \mult_22/S2_20_8  ( .A(\mult_22/ab[20][8] ), .B(
        \mult_22/CARRYB[19][8] ), .CI(\mult_22/SUMB[19][9] ), .CO(
        \mult_22/CARRYB[20][8] ), .S(\mult_22/SUMB[20][8] ) );
  FA_X1 \mult_22/S2_20_7  ( .A(\mult_22/ab[20][7] ), .B(
        \mult_22/CARRYB[19][7] ), .CI(\mult_22/SUMB[19][8] ), .CO(
        \mult_22/CARRYB[20][7] ), .S(\mult_22/SUMB[20][7] ) );
  FA_X1 \mult_22/S2_20_6  ( .A(\mult_22/ab[20][6] ), .B(
        \mult_22/CARRYB[19][6] ), .CI(\mult_22/SUMB[19][7] ), .CO(
        \mult_22/CARRYB[20][6] ), .S(\mult_22/SUMB[20][6] ) );
  FA_X1 \mult_22/S2_20_5  ( .A(\mult_22/ab[20][5] ), .B(
        \mult_22/CARRYB[19][5] ), .CI(\mult_22/SUMB[19][6] ), .CO(
        \mult_22/CARRYB[20][5] ), .S(\mult_22/SUMB[20][5] ) );
  FA_X1 \mult_22/S2_20_4  ( .A(\mult_22/ab[20][4] ), .B(
        \mult_22/CARRYB[19][4] ), .CI(\mult_22/SUMB[19][5] ), .CO(
        \mult_22/CARRYB[20][4] ), .S(\mult_22/SUMB[20][4] ) );
  FA_X1 \mult_22/S2_20_3  ( .A(\mult_22/ab[20][3] ), .B(
        \mult_22/CARRYB[19][3] ), .CI(\mult_22/SUMB[19][4] ), .CO(
        \mult_22/CARRYB[20][3] ), .S(\mult_22/SUMB[20][3] ) );
  FA_X1 \mult_22/S2_20_2  ( .A(\mult_22/ab[20][2] ), .B(
        \mult_22/CARRYB[19][2] ), .CI(\mult_22/SUMB[19][3] ), .CO(
        \mult_22/CARRYB[20][2] ), .S(\mult_22/SUMB[20][2] ) );
  FA_X1 \mult_22/S2_20_1  ( .A(\mult_22/ab[20][1] ), .B(
        \mult_22/CARRYB[19][1] ), .CI(\mult_22/SUMB[19][2] ), .CO(
        \mult_22/CARRYB[20][1] ), .S(\mult_22/SUMB[20][1] ) );
  FA_X1 \mult_22/S1_20_0  ( .A(\mult_22/ab[20][0] ), .B(
        \mult_22/CARRYB[19][0] ), .CI(\mult_22/SUMB[19][1] ), .CO(
        \mult_22/CARRYB[20][0] ), .S(N148) );
  FA_X1 \mult_22/S3_21_62  ( .A(\mult_22/ab[21][62] ), .B(
        \mult_22/CARRYB[20][62] ), .CI(\mult_22/ab[20][63] ), .CO(
        \mult_22/CARRYB[21][62] ), .S(\mult_22/SUMB[21][62] ) );
  FA_X1 \mult_22/S2_21_61  ( .A(\mult_22/ab[21][61] ), .B(
        \mult_22/CARRYB[20][61] ), .CI(\mult_22/SUMB[20][62] ), .CO(
        \mult_22/CARRYB[21][61] ), .S(\mult_22/SUMB[21][61] ) );
  FA_X1 \mult_22/S2_21_60  ( .A(\mult_22/ab[21][60] ), .B(
        \mult_22/CARRYB[20][60] ), .CI(\mult_22/SUMB[20][61] ), .CO(
        \mult_22/CARRYB[21][60] ), .S(\mult_22/SUMB[21][60] ) );
  FA_X1 \mult_22/S2_21_59  ( .A(\mult_22/ab[21][59] ), .B(
        \mult_22/CARRYB[20][59] ), .CI(\mult_22/SUMB[20][60] ), .CO(
        \mult_22/CARRYB[21][59] ), .S(\mult_22/SUMB[21][59] ) );
  FA_X1 \mult_22/S2_21_58  ( .A(\mult_22/ab[21][58] ), .B(
        \mult_22/CARRYB[20][58] ), .CI(\mult_22/SUMB[20][59] ), .CO(
        \mult_22/CARRYB[21][58] ), .S(\mult_22/SUMB[21][58] ) );
  FA_X1 \mult_22/S2_21_57  ( .A(\mult_22/ab[21][57] ), .B(
        \mult_22/CARRYB[20][57] ), .CI(\mult_22/SUMB[20][58] ), .CO(
        \mult_22/CARRYB[21][57] ), .S(\mult_22/SUMB[21][57] ) );
  FA_X1 \mult_22/S2_21_56  ( .A(\mult_22/ab[21][56] ), .B(
        \mult_22/CARRYB[20][56] ), .CI(\mult_22/SUMB[20][57] ), .CO(
        \mult_22/CARRYB[21][56] ), .S(\mult_22/SUMB[21][56] ) );
  FA_X1 \mult_22/S2_21_55  ( .A(\mult_22/ab[21][55] ), .B(
        \mult_22/CARRYB[20][55] ), .CI(\mult_22/SUMB[20][56] ), .CO(
        \mult_22/CARRYB[21][55] ), .S(\mult_22/SUMB[21][55] ) );
  FA_X1 \mult_22/S2_21_54  ( .A(\mult_22/ab[21][54] ), .B(
        \mult_22/CARRYB[20][54] ), .CI(\mult_22/SUMB[20][55] ), .CO(
        \mult_22/CARRYB[21][54] ), .S(\mult_22/SUMB[21][54] ) );
  FA_X1 \mult_22/S2_21_53  ( .A(\mult_22/ab[21][53] ), .B(
        \mult_22/CARRYB[20][53] ), .CI(\mult_22/SUMB[20][54] ), .CO(
        \mult_22/CARRYB[21][53] ), .S(\mult_22/SUMB[21][53] ) );
  FA_X1 \mult_22/S2_21_52  ( .A(\mult_22/ab[21][52] ), .B(
        \mult_22/CARRYB[20][52] ), .CI(\mult_22/SUMB[20][53] ), .CO(
        \mult_22/CARRYB[21][52] ), .S(\mult_22/SUMB[21][52] ) );
  FA_X1 \mult_22/S2_21_51  ( .A(\mult_22/ab[21][51] ), .B(
        \mult_22/CARRYB[20][51] ), .CI(\mult_22/SUMB[20][52] ), .CO(
        \mult_22/CARRYB[21][51] ), .S(\mult_22/SUMB[21][51] ) );
  FA_X1 \mult_22/S2_21_50  ( .A(\mult_22/ab[21][50] ), .B(
        \mult_22/CARRYB[20][50] ), .CI(\mult_22/SUMB[20][51] ), .CO(
        \mult_22/CARRYB[21][50] ), .S(\mult_22/SUMB[21][50] ) );
  FA_X1 \mult_22/S2_21_49  ( .A(\mult_22/ab[21][49] ), .B(
        \mult_22/CARRYB[20][49] ), .CI(\mult_22/SUMB[20][50] ), .CO(
        \mult_22/CARRYB[21][49] ), .S(\mult_22/SUMB[21][49] ) );
  FA_X1 \mult_22/S2_21_48  ( .A(\mult_22/ab[21][48] ), .B(
        \mult_22/CARRYB[20][48] ), .CI(\mult_22/SUMB[20][49] ), .CO(
        \mult_22/CARRYB[21][48] ), .S(\mult_22/SUMB[21][48] ) );
  FA_X1 \mult_22/S2_21_47  ( .A(\mult_22/ab[21][47] ), .B(
        \mult_22/CARRYB[20][47] ), .CI(\mult_22/SUMB[20][48] ), .CO(
        \mult_22/CARRYB[21][47] ), .S(\mult_22/SUMB[21][47] ) );
  FA_X1 \mult_22/S2_21_46  ( .A(\mult_22/CARRYB[20][46] ), .B(
        \mult_22/ab[21][46] ), .CI(\mult_22/SUMB[20][47] ), .CO(
        \mult_22/CARRYB[21][46] ), .S(\mult_22/SUMB[21][46] ) );
  FA_X1 \mult_22/S2_21_45  ( .A(\mult_22/ab[21][45] ), .B(
        \mult_22/CARRYB[20][45] ), .CI(\mult_22/SUMB[20][46] ), .CO(
        \mult_22/CARRYB[21][45] ), .S(\mult_22/SUMB[21][45] ) );
  FA_X1 \mult_22/S2_21_42  ( .A(\mult_22/ab[21][42] ), .B(
        \mult_22/CARRYB[20][42] ), .CI(\mult_22/SUMB[20][43] ), .CO(
        \mult_22/CARRYB[21][42] ), .S(\mult_22/SUMB[21][42] ) );
  FA_X1 \mult_22/S2_21_41  ( .A(\mult_22/ab[21][41] ), .B(
        \mult_22/CARRYB[20][41] ), .CI(\mult_22/SUMB[20][42] ), .CO(
        \mult_22/CARRYB[21][41] ), .S(\mult_22/SUMB[21][41] ) );
  FA_X1 \mult_22/S2_21_40  ( .A(\mult_22/ab[21][40] ), .B(
        \mult_22/CARRYB[20][40] ), .CI(\mult_22/SUMB[20][41] ), .CO(
        \mult_22/CARRYB[21][40] ), .S(\mult_22/SUMB[21][40] ) );
  FA_X1 \mult_22/S2_21_39  ( .A(\mult_22/ab[21][39] ), .B(
        \mult_22/CARRYB[20][39] ), .CI(\mult_22/SUMB[20][40] ), .CO(
        \mult_22/CARRYB[21][39] ), .S(\mult_22/SUMB[21][39] ) );
  FA_X1 \mult_22/S2_21_37  ( .A(\mult_22/ab[21][37] ), .B(
        \mult_22/CARRYB[20][37] ), .CI(\mult_22/SUMB[20][38] ), .CO(
        \mult_22/CARRYB[21][37] ), .S(\mult_22/SUMB[21][37] ) );
  FA_X1 \mult_22/S2_21_35  ( .A(\mult_22/ab[21][35] ), .B(
        \mult_22/CARRYB[20][35] ), .CI(\mult_22/SUMB[20][36] ), .CO(
        \mult_22/CARRYB[21][35] ), .S(\mult_22/SUMB[21][35] ) );
  FA_X1 \mult_22/S2_21_34  ( .A(\mult_22/ab[21][34] ), .B(
        \mult_22/CARRYB[20][34] ), .CI(\mult_22/SUMB[20][35] ), .CO(
        \mult_22/CARRYB[21][34] ), .S(\mult_22/SUMB[21][34] ) );
  FA_X1 \mult_22/S2_21_33  ( .A(\mult_22/ab[21][33] ), .B(
        \mult_22/CARRYB[20][33] ), .CI(\mult_22/SUMB[20][34] ), .CO(
        \mult_22/CARRYB[21][33] ), .S(\mult_22/SUMB[21][33] ) );
  FA_X1 \mult_22/S2_21_32  ( .A(\mult_22/ab[21][32] ), .B(
        \mult_22/CARRYB[20][32] ), .CI(\mult_22/SUMB[20][33] ), .CO(
        \mult_22/CARRYB[21][32] ), .S(\mult_22/SUMB[21][32] ) );
  FA_X1 \mult_22/S2_21_31  ( .A(\mult_22/ab[21][31] ), .B(
        \mult_22/CARRYB[20][31] ), .CI(\mult_22/SUMB[20][32] ), .CO(
        \mult_22/CARRYB[21][31] ), .S(\mult_22/SUMB[21][31] ) );
  FA_X1 \mult_22/S2_21_30  ( .A(\mult_22/ab[21][30] ), .B(
        \mult_22/CARRYB[20][30] ), .CI(\mult_22/SUMB[20][31] ), .CO(
        \mult_22/CARRYB[21][30] ), .S(\mult_22/SUMB[21][30] ) );
  FA_X1 \mult_22/S2_21_29  ( .A(\mult_22/ab[21][29] ), .B(
        \mult_22/CARRYB[20][29] ), .CI(\mult_22/SUMB[20][30] ), .CO(
        \mult_22/CARRYB[21][29] ), .S(\mult_22/SUMB[21][29] ) );
  FA_X1 \mult_22/S2_21_28  ( .A(\mult_22/ab[21][28] ), .B(
        \mult_22/CARRYB[20][28] ), .CI(\mult_22/SUMB[20][29] ), .CO(
        \mult_22/CARRYB[21][28] ), .S(\mult_22/SUMB[21][28] ) );
  FA_X1 \mult_22/S2_21_27  ( .A(\mult_22/ab[21][27] ), .B(
        \mult_22/CARRYB[20][27] ), .CI(\mult_22/SUMB[20][28] ), .CO(
        \mult_22/CARRYB[21][27] ), .S(\mult_22/SUMB[21][27] ) );
  FA_X1 \mult_22/S2_21_26  ( .A(\mult_22/ab[21][26] ), .B(
        \mult_22/CARRYB[20][26] ), .CI(\mult_22/SUMB[20][27] ), .CO(
        \mult_22/CARRYB[21][26] ), .S(\mult_22/SUMB[21][26] ) );
  FA_X1 \mult_22/S2_21_25  ( .A(\mult_22/ab[21][25] ), .B(
        \mult_22/CARRYB[20][25] ), .CI(\mult_22/SUMB[20][26] ), .CO(
        \mult_22/CARRYB[21][25] ), .S(\mult_22/SUMB[21][25] ) );
  FA_X1 \mult_22/S2_21_24  ( .A(\mult_22/ab[21][24] ), .B(
        \mult_22/CARRYB[20][24] ), .CI(\mult_22/SUMB[20][25] ), .CO(
        \mult_22/CARRYB[21][24] ), .S(\mult_22/SUMB[21][24] ) );
  FA_X1 \mult_22/S2_21_23  ( .A(\mult_22/ab[21][23] ), .B(
        \mult_22/CARRYB[20][23] ), .CI(\mult_22/SUMB[20][24] ), .CO(
        \mult_22/CARRYB[21][23] ), .S(\mult_22/SUMB[21][23] ) );
  FA_X1 \mult_22/S2_21_22  ( .A(\mult_22/ab[21][22] ), .B(
        \mult_22/CARRYB[20][22] ), .CI(\mult_22/SUMB[20][23] ), .CO(
        \mult_22/CARRYB[21][22] ), .S(\mult_22/SUMB[21][22] ) );
  FA_X1 \mult_22/S2_21_21  ( .A(\mult_22/ab[21][21] ), .B(
        \mult_22/CARRYB[20][21] ), .CI(\mult_22/SUMB[20][22] ), .CO(
        \mult_22/CARRYB[21][21] ), .S(\mult_22/SUMB[21][21] ) );
  FA_X1 \mult_22/S2_21_20  ( .A(\mult_22/ab[21][20] ), .B(
        \mult_22/CARRYB[20][20] ), .CI(\mult_22/SUMB[20][21] ), .CO(
        \mult_22/CARRYB[21][20] ), .S(\mult_22/SUMB[21][20] ) );
  FA_X1 \mult_22/S2_21_19  ( .A(\mult_22/ab[21][19] ), .B(
        \mult_22/CARRYB[20][19] ), .CI(\mult_22/SUMB[20][20] ), .CO(
        \mult_22/CARRYB[21][19] ), .S(\mult_22/SUMB[21][19] ) );
  FA_X1 \mult_22/S2_21_18  ( .A(\mult_22/ab[21][18] ), .B(
        \mult_22/CARRYB[20][18] ), .CI(\mult_22/SUMB[20][19] ), .CO(
        \mult_22/CARRYB[21][18] ), .S(\mult_22/SUMB[21][18] ) );
  FA_X1 \mult_22/S2_21_17  ( .A(\mult_22/ab[21][17] ), .B(
        \mult_22/CARRYB[20][17] ), .CI(\mult_22/SUMB[20][18] ), .CO(
        \mult_22/CARRYB[21][17] ), .S(\mult_22/SUMB[21][17] ) );
  FA_X1 \mult_22/S2_21_16  ( .A(\mult_22/ab[21][16] ), .B(
        \mult_22/CARRYB[20][16] ), .CI(\mult_22/SUMB[20][17] ), .CO(
        \mult_22/CARRYB[21][16] ), .S(\mult_22/SUMB[21][16] ) );
  FA_X1 \mult_22/S2_21_15  ( .A(\mult_22/ab[21][15] ), .B(
        \mult_22/CARRYB[20][15] ), .CI(\mult_22/SUMB[20][16] ), .CO(
        \mult_22/CARRYB[21][15] ), .S(\mult_22/SUMB[21][15] ) );
  FA_X1 \mult_22/S2_21_14  ( .A(\mult_22/ab[21][14] ), .B(
        \mult_22/CARRYB[20][14] ), .CI(\mult_22/SUMB[20][15] ), .CO(
        \mult_22/CARRYB[21][14] ), .S(\mult_22/SUMB[21][14] ) );
  FA_X1 \mult_22/S2_21_13  ( .A(\mult_22/ab[21][13] ), .B(
        \mult_22/CARRYB[20][13] ), .CI(\mult_22/SUMB[20][14] ), .CO(
        \mult_22/CARRYB[21][13] ), .S(\mult_22/SUMB[21][13] ) );
  FA_X1 \mult_22/S2_21_12  ( .A(\mult_22/ab[21][12] ), .B(
        \mult_22/CARRYB[20][12] ), .CI(\mult_22/SUMB[20][13] ), .CO(
        \mult_22/CARRYB[21][12] ), .S(\mult_22/SUMB[21][12] ) );
  FA_X1 \mult_22/S2_21_11  ( .A(\mult_22/ab[21][11] ), .B(
        \mult_22/CARRYB[20][11] ), .CI(\mult_22/SUMB[20][12] ), .CO(
        \mult_22/CARRYB[21][11] ), .S(\mult_22/SUMB[21][11] ) );
  FA_X1 \mult_22/S2_21_10  ( .A(\mult_22/ab[21][10] ), .B(
        \mult_22/CARRYB[20][10] ), .CI(\mult_22/SUMB[20][11] ), .CO(
        \mult_22/CARRYB[21][10] ), .S(\mult_22/SUMB[21][10] ) );
  FA_X1 \mult_22/S2_21_9  ( .A(\mult_22/ab[21][9] ), .B(
        \mult_22/CARRYB[20][9] ), .CI(\mult_22/SUMB[20][10] ), .CO(
        \mult_22/CARRYB[21][9] ), .S(\mult_22/SUMB[21][9] ) );
  FA_X1 \mult_22/S2_21_8  ( .A(\mult_22/ab[21][8] ), .B(
        \mult_22/CARRYB[20][8] ), .CI(\mult_22/SUMB[20][9] ), .CO(
        \mult_22/CARRYB[21][8] ), .S(\mult_22/SUMB[21][8] ) );
  FA_X1 \mult_22/S2_21_7  ( .A(\mult_22/ab[21][7] ), .B(
        \mult_22/CARRYB[20][7] ), .CI(\mult_22/SUMB[20][8] ), .CO(
        \mult_22/CARRYB[21][7] ), .S(\mult_22/SUMB[21][7] ) );
  FA_X1 \mult_22/S2_21_6  ( .A(\mult_22/ab[21][6] ), .B(
        \mult_22/CARRYB[20][6] ), .CI(\mult_22/SUMB[20][7] ), .CO(
        \mult_22/CARRYB[21][6] ), .S(\mult_22/SUMB[21][6] ) );
  FA_X1 \mult_22/S2_21_5  ( .A(\mult_22/ab[21][5] ), .B(
        \mult_22/CARRYB[20][5] ), .CI(\mult_22/SUMB[20][6] ), .CO(
        \mult_22/CARRYB[21][5] ), .S(\mult_22/SUMB[21][5] ) );
  FA_X1 \mult_22/S2_21_4  ( .A(\mult_22/ab[21][4] ), .B(
        \mult_22/CARRYB[20][4] ), .CI(\mult_22/SUMB[20][5] ), .CO(
        \mult_22/CARRYB[21][4] ), .S(\mult_22/SUMB[21][4] ) );
  FA_X1 \mult_22/S2_21_3  ( .A(\mult_22/ab[21][3] ), .B(
        \mult_22/CARRYB[20][3] ), .CI(\mult_22/SUMB[20][4] ), .CO(
        \mult_22/CARRYB[21][3] ), .S(\mult_22/SUMB[21][3] ) );
  FA_X1 \mult_22/S2_21_2  ( .A(\mult_22/ab[21][2] ), .B(
        \mult_22/CARRYB[20][2] ), .CI(\mult_22/SUMB[20][3] ), .CO(
        \mult_22/CARRYB[21][2] ), .S(\mult_22/SUMB[21][2] ) );
  FA_X1 \mult_22/S2_21_1  ( .A(\mult_22/ab[21][1] ), .B(
        \mult_22/CARRYB[20][1] ), .CI(\mult_22/SUMB[20][2] ), .CO(
        \mult_22/CARRYB[21][1] ), .S(\mult_22/SUMB[21][1] ) );
  FA_X1 \mult_22/S1_21_0  ( .A(\mult_22/ab[21][0] ), .B(
        \mult_22/CARRYB[20][0] ), .CI(\mult_22/SUMB[20][1] ), .CO(
        \mult_22/CARRYB[21][0] ), .S(N149) );
  FA_X1 \mult_22/S3_22_62  ( .A(\mult_22/ab[22][62] ), .B(
        \mult_22/CARRYB[21][62] ), .CI(\mult_22/ab[21][63] ), .CO(
        \mult_22/CARRYB[22][62] ), .S(\mult_22/SUMB[22][62] ) );
  FA_X1 \mult_22/S2_22_61  ( .A(\mult_22/ab[22][61] ), .B(
        \mult_22/CARRYB[21][61] ), .CI(\mult_22/SUMB[21][62] ), .CO(
        \mult_22/CARRYB[22][61] ), .S(\mult_22/SUMB[22][61] ) );
  FA_X1 \mult_22/S2_22_60  ( .A(\mult_22/ab[22][60] ), .B(
        \mult_22/CARRYB[21][60] ), .CI(\mult_22/SUMB[21][61] ), .CO(
        \mult_22/CARRYB[22][60] ), .S(\mult_22/SUMB[22][60] ) );
  FA_X1 \mult_22/S2_22_59  ( .A(\mult_22/ab[22][59] ), .B(
        \mult_22/CARRYB[21][59] ), .CI(\mult_22/SUMB[21][60] ), .CO(
        \mult_22/CARRYB[22][59] ), .S(\mult_22/SUMB[22][59] ) );
  FA_X1 \mult_22/S2_22_58  ( .A(\mult_22/ab[22][58] ), .B(
        \mult_22/CARRYB[21][58] ), .CI(\mult_22/SUMB[21][59] ), .CO(
        \mult_22/CARRYB[22][58] ), .S(\mult_22/SUMB[22][58] ) );
  FA_X1 \mult_22/S2_22_57  ( .A(\mult_22/ab[22][57] ), .B(
        \mult_22/CARRYB[21][57] ), .CI(\mult_22/SUMB[21][58] ), .CO(
        \mult_22/CARRYB[22][57] ), .S(\mult_22/SUMB[22][57] ) );
  FA_X1 \mult_22/S2_22_56  ( .A(\mult_22/ab[22][56] ), .B(
        \mult_22/CARRYB[21][56] ), .CI(\mult_22/SUMB[21][57] ), .CO(
        \mult_22/CARRYB[22][56] ), .S(\mult_22/SUMB[22][56] ) );
  FA_X1 \mult_22/S2_22_55  ( .A(\mult_22/ab[22][55] ), .B(
        \mult_22/CARRYB[21][55] ), .CI(\mult_22/SUMB[21][56] ), .CO(
        \mult_22/CARRYB[22][55] ), .S(\mult_22/SUMB[22][55] ) );
  FA_X1 \mult_22/S2_22_54  ( .A(\mult_22/ab[22][54] ), .B(
        \mult_22/CARRYB[21][54] ), .CI(\mult_22/SUMB[21][55] ), .CO(
        \mult_22/CARRYB[22][54] ), .S(\mult_22/SUMB[22][54] ) );
  FA_X1 \mult_22/S2_22_53  ( .A(\mult_22/ab[22][53] ), .B(
        \mult_22/CARRYB[21][53] ), .CI(\mult_22/SUMB[21][54] ), .CO(
        \mult_22/CARRYB[22][53] ), .S(\mult_22/SUMB[22][53] ) );
  FA_X1 \mult_22/S2_22_52  ( .A(\mult_22/ab[22][52] ), .B(
        \mult_22/CARRYB[21][52] ), .CI(\mult_22/SUMB[21][53] ), .CO(
        \mult_22/CARRYB[22][52] ), .S(\mult_22/SUMB[22][52] ) );
  FA_X1 \mult_22/S2_22_51  ( .A(\mult_22/ab[22][51] ), .B(
        \mult_22/CARRYB[21][51] ), .CI(\mult_22/SUMB[21][52] ), .CO(
        \mult_22/CARRYB[22][51] ), .S(\mult_22/SUMB[22][51] ) );
  FA_X1 \mult_22/S2_22_50  ( .A(\mult_22/ab[22][50] ), .B(
        \mult_22/CARRYB[21][50] ), .CI(\mult_22/SUMB[21][51] ), .CO(
        \mult_22/CARRYB[22][50] ), .S(\mult_22/SUMB[22][50] ) );
  FA_X1 \mult_22/S2_22_49  ( .A(\mult_22/ab[22][49] ), .B(
        \mult_22/CARRYB[21][49] ), .CI(\mult_22/SUMB[21][50] ), .CO(
        \mult_22/CARRYB[22][49] ), .S(\mult_22/SUMB[22][49] ) );
  FA_X1 \mult_22/S2_22_48  ( .A(\mult_22/ab[22][48] ), .B(
        \mult_22/CARRYB[21][48] ), .CI(\mult_22/SUMB[21][49] ), .CO(
        \mult_22/CARRYB[22][48] ), .S(\mult_22/SUMB[22][48] ) );
  FA_X1 \mult_22/S2_22_47  ( .A(\mult_22/ab[22][47] ), .B(
        \mult_22/CARRYB[21][47] ), .CI(\mult_22/SUMB[21][48] ), .CO(
        \mult_22/CARRYB[22][47] ), .S(\mult_22/SUMB[22][47] ) );
  FA_X1 \mult_22/S2_22_46  ( .A(\mult_22/ab[22][46] ), .B(
        \mult_22/CARRYB[21][46] ), .CI(\mult_22/SUMB[21][47] ), .CO(
        \mult_22/CARRYB[22][46] ), .S(\mult_22/SUMB[22][46] ) );
  FA_X1 \mult_22/S2_22_45  ( .A(\mult_22/ab[22][45] ), .B(
        \mult_22/CARRYB[21][45] ), .CI(\mult_22/SUMB[21][46] ), .CO(
        \mult_22/CARRYB[22][45] ), .S(\mult_22/SUMB[22][45] ) );
  FA_X1 \mult_22/S2_22_44  ( .A(\mult_22/CARRYB[21][44] ), .B(
        \mult_22/ab[22][44] ), .CI(\mult_22/SUMB[21][45] ), .CO(
        \mult_22/CARRYB[22][44] ), .S(\mult_22/SUMB[22][44] ) );
  FA_X1 \mult_22/S2_22_43  ( .A(\mult_22/ab[22][43] ), .B(
        \mult_22/CARRYB[21][43] ), .CI(\mult_22/SUMB[21][44] ), .CO(
        \mult_22/CARRYB[22][43] ), .S(\mult_22/SUMB[22][43] ) );
  FA_X1 \mult_22/S2_22_42  ( .A(\mult_22/ab[22][42] ), .B(
        \mult_22/CARRYB[21][42] ), .CI(\mult_22/SUMB[21][43] ), .CO(
        \mult_22/CARRYB[22][42] ), .S(\mult_22/SUMB[22][42] ) );
  FA_X1 \mult_22/S2_22_41  ( .A(\mult_22/ab[22][41] ), .B(
        \mult_22/CARRYB[21][41] ), .CI(\mult_22/SUMB[21][42] ), .CO(
        \mult_22/CARRYB[22][41] ), .S(\mult_22/SUMB[22][41] ) );
  FA_X1 \mult_22/S2_22_40  ( .A(\mult_22/ab[22][40] ), .B(
        \mult_22/CARRYB[21][40] ), .CI(\mult_22/SUMB[21][41] ), .CO(
        \mult_22/CARRYB[22][40] ), .S(\mult_22/SUMB[22][40] ) );
  FA_X1 \mult_22/S2_22_39  ( .A(\mult_22/CARRYB[21][39] ), .B(
        \mult_22/ab[22][39] ), .CI(\mult_22/SUMB[21][40] ), .CO(
        \mult_22/CARRYB[22][39] ), .S(\mult_22/SUMB[22][39] ) );
  FA_X1 \mult_22/S2_22_37  ( .A(\mult_22/ab[22][37] ), .B(
        \mult_22/CARRYB[21][37] ), .CI(\mult_22/SUMB[21][38] ), .CO(
        \mult_22/CARRYB[22][37] ), .S(\mult_22/SUMB[22][37] ) );
  FA_X1 \mult_22/S2_22_36  ( .A(\mult_22/ab[22][36] ), .B(
        \mult_22/CARRYB[21][36] ), .CI(\mult_22/SUMB[21][37] ), .CO(
        \mult_22/CARRYB[22][36] ), .S(\mult_22/SUMB[22][36] ) );
  FA_X1 \mult_22/S2_22_35  ( .A(\mult_22/ab[22][35] ), .B(
        \mult_22/CARRYB[21][35] ), .CI(\mult_22/SUMB[21][36] ), .CO(
        \mult_22/CARRYB[22][35] ), .S(\mult_22/SUMB[22][35] ) );
  FA_X1 \mult_22/S2_22_34  ( .A(\mult_22/ab[22][34] ), .B(
        \mult_22/CARRYB[21][34] ), .CI(\mult_22/SUMB[21][35] ), .CO(
        \mult_22/CARRYB[22][34] ), .S(\mult_22/SUMB[22][34] ) );
  FA_X1 \mult_22/S2_22_33  ( .A(\mult_22/ab[22][33] ), .B(
        \mult_22/CARRYB[21][33] ), .CI(\mult_22/SUMB[21][34] ), .CO(
        \mult_22/CARRYB[22][33] ), .S(\mult_22/SUMB[22][33] ) );
  FA_X1 \mult_22/S2_22_32  ( .A(\mult_22/ab[22][32] ), .B(
        \mult_22/CARRYB[21][32] ), .CI(\mult_22/SUMB[21][33] ), .CO(
        \mult_22/CARRYB[22][32] ), .S(\mult_22/SUMB[22][32] ) );
  FA_X1 \mult_22/S2_22_31  ( .A(\mult_22/ab[22][31] ), .B(
        \mult_22/CARRYB[21][31] ), .CI(\mult_22/SUMB[21][32] ), .CO(
        \mult_22/CARRYB[22][31] ), .S(\mult_22/SUMB[22][31] ) );
  FA_X1 \mult_22/S2_22_30  ( .A(\mult_22/ab[22][30] ), .B(
        \mult_22/CARRYB[21][30] ), .CI(\mult_22/SUMB[21][31] ), .CO(
        \mult_22/CARRYB[22][30] ), .S(\mult_22/SUMB[22][30] ) );
  FA_X1 \mult_22/S2_22_29  ( .A(\mult_22/ab[22][29] ), .B(
        \mult_22/CARRYB[21][29] ), .CI(\mult_22/SUMB[21][30] ), .CO(
        \mult_22/CARRYB[22][29] ), .S(\mult_22/SUMB[22][29] ) );
  FA_X1 \mult_22/S2_22_28  ( .A(\mult_22/ab[22][28] ), .B(
        \mult_22/CARRYB[21][28] ), .CI(\mult_22/SUMB[21][29] ), .CO(
        \mult_22/CARRYB[22][28] ), .S(\mult_22/SUMB[22][28] ) );
  FA_X1 \mult_22/S2_22_27  ( .A(\mult_22/ab[22][27] ), .B(
        \mult_22/CARRYB[21][27] ), .CI(\mult_22/SUMB[21][28] ), .CO(
        \mult_22/CARRYB[22][27] ), .S(\mult_22/SUMB[22][27] ) );
  FA_X1 \mult_22/S2_22_26  ( .A(\mult_22/ab[22][26] ), .B(
        \mult_22/CARRYB[21][26] ), .CI(\mult_22/SUMB[21][27] ), .CO(
        \mult_22/CARRYB[22][26] ), .S(\mult_22/SUMB[22][26] ) );
  FA_X1 \mult_22/S2_22_25  ( .A(\mult_22/ab[22][25] ), .B(
        \mult_22/CARRYB[21][25] ), .CI(\mult_22/SUMB[21][26] ), .CO(
        \mult_22/CARRYB[22][25] ), .S(\mult_22/SUMB[22][25] ) );
  FA_X1 \mult_22/S2_22_24  ( .A(\mult_22/ab[22][24] ), .B(
        \mult_22/CARRYB[21][24] ), .CI(\mult_22/SUMB[21][25] ), .CO(
        \mult_22/CARRYB[22][24] ), .S(\mult_22/SUMB[22][24] ) );
  FA_X1 \mult_22/S2_22_23  ( .A(\mult_22/ab[22][23] ), .B(
        \mult_22/CARRYB[21][23] ), .CI(\mult_22/SUMB[21][24] ), .CO(
        \mult_22/CARRYB[22][23] ), .S(\mult_22/SUMB[22][23] ) );
  FA_X1 \mult_22/S2_22_22  ( .A(\mult_22/ab[22][22] ), .B(
        \mult_22/CARRYB[21][22] ), .CI(\mult_22/SUMB[21][23] ), .CO(
        \mult_22/CARRYB[22][22] ), .S(\mult_22/SUMB[22][22] ) );
  FA_X1 \mult_22/S2_22_21  ( .A(\mult_22/ab[22][21] ), .B(
        \mult_22/CARRYB[21][21] ), .CI(\mult_22/SUMB[21][22] ), .CO(
        \mult_22/CARRYB[22][21] ), .S(\mult_22/SUMB[22][21] ) );
  FA_X1 \mult_22/S2_22_20  ( .A(\mult_22/ab[22][20] ), .B(
        \mult_22/CARRYB[21][20] ), .CI(\mult_22/SUMB[21][21] ), .CO(
        \mult_22/CARRYB[22][20] ), .S(\mult_22/SUMB[22][20] ) );
  FA_X1 \mult_22/S2_22_19  ( .A(\mult_22/ab[22][19] ), .B(
        \mult_22/CARRYB[21][19] ), .CI(\mult_22/SUMB[21][20] ), .CO(
        \mult_22/CARRYB[22][19] ), .S(\mult_22/SUMB[22][19] ) );
  FA_X1 \mult_22/S2_22_18  ( .A(\mult_22/ab[22][18] ), .B(
        \mult_22/CARRYB[21][18] ), .CI(\mult_22/SUMB[21][19] ), .CO(
        \mult_22/CARRYB[22][18] ), .S(\mult_22/SUMB[22][18] ) );
  FA_X1 \mult_22/S2_22_17  ( .A(\mult_22/ab[22][17] ), .B(
        \mult_22/CARRYB[21][17] ), .CI(\mult_22/SUMB[21][18] ), .CO(
        \mult_22/CARRYB[22][17] ), .S(\mult_22/SUMB[22][17] ) );
  FA_X1 \mult_22/S2_22_16  ( .A(\mult_22/ab[22][16] ), .B(
        \mult_22/CARRYB[21][16] ), .CI(\mult_22/SUMB[21][17] ), .CO(
        \mult_22/CARRYB[22][16] ), .S(\mult_22/SUMB[22][16] ) );
  FA_X1 \mult_22/S2_22_15  ( .A(\mult_22/ab[22][15] ), .B(
        \mult_22/CARRYB[21][15] ), .CI(\mult_22/SUMB[21][16] ), .CO(
        \mult_22/CARRYB[22][15] ), .S(\mult_22/SUMB[22][15] ) );
  FA_X1 \mult_22/S2_22_14  ( .A(\mult_22/ab[22][14] ), .B(
        \mult_22/CARRYB[21][14] ), .CI(\mult_22/SUMB[21][15] ), .CO(
        \mult_22/CARRYB[22][14] ), .S(\mult_22/SUMB[22][14] ) );
  FA_X1 \mult_22/S2_22_13  ( .A(\mult_22/ab[22][13] ), .B(
        \mult_22/CARRYB[21][13] ), .CI(\mult_22/SUMB[21][14] ), .CO(
        \mult_22/CARRYB[22][13] ), .S(\mult_22/SUMB[22][13] ) );
  FA_X1 \mult_22/S2_22_12  ( .A(\mult_22/ab[22][12] ), .B(
        \mult_22/CARRYB[21][12] ), .CI(\mult_22/SUMB[21][13] ), .CO(
        \mult_22/CARRYB[22][12] ), .S(\mult_22/SUMB[22][12] ) );
  FA_X1 \mult_22/S2_22_11  ( .A(\mult_22/ab[22][11] ), .B(
        \mult_22/CARRYB[21][11] ), .CI(\mult_22/SUMB[21][12] ), .CO(
        \mult_22/CARRYB[22][11] ), .S(\mult_22/SUMB[22][11] ) );
  FA_X1 \mult_22/S2_22_10  ( .A(\mult_22/ab[22][10] ), .B(
        \mult_22/CARRYB[21][10] ), .CI(\mult_22/SUMB[21][11] ), .CO(
        \mult_22/CARRYB[22][10] ), .S(\mult_22/SUMB[22][10] ) );
  FA_X1 \mult_22/S2_22_9  ( .A(\mult_22/ab[22][9] ), .B(
        \mult_22/CARRYB[21][9] ), .CI(\mult_22/SUMB[21][10] ), .CO(
        \mult_22/CARRYB[22][9] ), .S(\mult_22/SUMB[22][9] ) );
  FA_X1 \mult_22/S2_22_8  ( .A(\mult_22/ab[22][8] ), .B(
        \mult_22/CARRYB[21][8] ), .CI(\mult_22/SUMB[21][9] ), .CO(
        \mult_22/CARRYB[22][8] ), .S(\mult_22/SUMB[22][8] ) );
  FA_X1 \mult_22/S2_22_7  ( .A(\mult_22/ab[22][7] ), .B(
        \mult_22/CARRYB[21][7] ), .CI(\mult_22/SUMB[21][8] ), .CO(
        \mult_22/CARRYB[22][7] ), .S(\mult_22/SUMB[22][7] ) );
  FA_X1 \mult_22/S2_22_6  ( .A(\mult_22/ab[22][6] ), .B(
        \mult_22/CARRYB[21][6] ), .CI(\mult_22/SUMB[21][7] ), .CO(
        \mult_22/CARRYB[22][6] ), .S(\mult_22/SUMB[22][6] ) );
  FA_X1 \mult_22/S2_22_5  ( .A(\mult_22/ab[22][5] ), .B(
        \mult_22/CARRYB[21][5] ), .CI(\mult_22/SUMB[21][6] ), .CO(
        \mult_22/CARRYB[22][5] ), .S(\mult_22/SUMB[22][5] ) );
  FA_X1 \mult_22/S2_22_4  ( .A(\mult_22/ab[22][4] ), .B(
        \mult_22/CARRYB[21][4] ), .CI(\mult_22/SUMB[21][5] ), .CO(
        \mult_22/CARRYB[22][4] ), .S(\mult_22/SUMB[22][4] ) );
  FA_X1 \mult_22/S2_22_3  ( .A(\mult_22/ab[22][3] ), .B(
        \mult_22/CARRYB[21][3] ), .CI(\mult_22/SUMB[21][4] ), .CO(
        \mult_22/CARRYB[22][3] ), .S(\mult_22/SUMB[22][3] ) );
  FA_X1 \mult_22/S2_22_2  ( .A(\mult_22/ab[22][2] ), .B(
        \mult_22/CARRYB[21][2] ), .CI(\mult_22/SUMB[21][3] ), .CO(
        \mult_22/CARRYB[22][2] ), .S(\mult_22/SUMB[22][2] ) );
  FA_X1 \mult_22/S2_22_1  ( .A(\mult_22/ab[22][1] ), .B(
        \mult_22/CARRYB[21][1] ), .CI(\mult_22/SUMB[21][2] ), .CO(
        \mult_22/CARRYB[22][1] ), .S(\mult_22/SUMB[22][1] ) );
  FA_X1 \mult_22/S1_22_0  ( .A(\mult_22/ab[22][0] ), .B(
        \mult_22/CARRYB[21][0] ), .CI(\mult_22/SUMB[21][1] ), .CO(
        \mult_22/CARRYB[22][0] ), .S(N150) );
  FA_X1 \mult_22/S3_23_62  ( .A(\mult_22/ab[23][62] ), .B(
        \mult_22/CARRYB[22][62] ), .CI(\mult_22/ab[22][63] ), .CO(
        \mult_22/CARRYB[23][62] ), .S(\mult_22/SUMB[23][62] ) );
  FA_X1 \mult_22/S2_23_61  ( .A(\mult_22/ab[23][61] ), .B(
        \mult_22/CARRYB[22][61] ), .CI(\mult_22/SUMB[22][62] ), .CO(
        \mult_22/CARRYB[23][61] ), .S(\mult_22/SUMB[23][61] ) );
  FA_X1 \mult_22/S2_23_60  ( .A(\mult_22/ab[23][60] ), .B(
        \mult_22/CARRYB[22][60] ), .CI(\mult_22/SUMB[22][61] ), .CO(
        \mult_22/CARRYB[23][60] ), .S(\mult_22/SUMB[23][60] ) );
  FA_X1 \mult_22/S2_23_59  ( .A(\mult_22/ab[23][59] ), .B(
        \mult_22/CARRYB[22][59] ), .CI(\mult_22/SUMB[22][60] ), .CO(
        \mult_22/CARRYB[23][59] ), .S(\mult_22/SUMB[23][59] ) );
  FA_X1 \mult_22/S2_23_58  ( .A(\mult_22/ab[23][58] ), .B(
        \mult_22/CARRYB[22][58] ), .CI(\mult_22/SUMB[22][59] ), .CO(
        \mult_22/CARRYB[23][58] ), .S(\mult_22/SUMB[23][58] ) );
  FA_X1 \mult_22/S2_23_57  ( .A(\mult_22/ab[23][57] ), .B(
        \mult_22/CARRYB[22][57] ), .CI(\mult_22/SUMB[22][58] ), .CO(
        \mult_22/CARRYB[23][57] ), .S(\mult_22/SUMB[23][57] ) );
  FA_X1 \mult_22/S2_23_56  ( .A(\mult_22/ab[23][56] ), .B(
        \mult_22/CARRYB[22][56] ), .CI(\mult_22/SUMB[22][57] ), .CO(
        \mult_22/CARRYB[23][56] ), .S(\mult_22/SUMB[23][56] ) );
  FA_X1 \mult_22/S2_23_55  ( .A(\mult_22/ab[23][55] ), .B(
        \mult_22/CARRYB[22][55] ), .CI(\mult_22/SUMB[22][56] ), .CO(
        \mult_22/CARRYB[23][55] ), .S(\mult_22/SUMB[23][55] ) );
  FA_X1 \mult_22/S2_23_54  ( .A(\mult_22/ab[23][54] ), .B(
        \mult_22/CARRYB[22][54] ), .CI(\mult_22/SUMB[22][55] ), .CO(
        \mult_22/CARRYB[23][54] ), .S(\mult_22/SUMB[23][54] ) );
  FA_X1 \mult_22/S2_23_53  ( .A(\mult_22/ab[23][53] ), .B(
        \mult_22/CARRYB[22][53] ), .CI(\mult_22/SUMB[22][54] ), .CO(
        \mult_22/CARRYB[23][53] ), .S(\mult_22/SUMB[23][53] ) );
  FA_X1 \mult_22/S2_23_52  ( .A(\mult_22/ab[23][52] ), .B(
        \mult_22/CARRYB[22][52] ), .CI(\mult_22/SUMB[22][53] ), .CO(
        \mult_22/CARRYB[23][52] ), .S(\mult_22/SUMB[23][52] ) );
  FA_X1 \mult_22/S2_23_51  ( .A(\mult_22/ab[23][51] ), .B(
        \mult_22/CARRYB[22][51] ), .CI(\mult_22/SUMB[22][52] ), .CO(
        \mult_22/CARRYB[23][51] ), .S(\mult_22/SUMB[23][51] ) );
  FA_X1 \mult_22/S2_23_50  ( .A(\mult_22/ab[23][50] ), .B(
        \mult_22/CARRYB[22][50] ), .CI(\mult_22/SUMB[22][51] ), .CO(
        \mult_22/CARRYB[23][50] ), .S(\mult_22/SUMB[23][50] ) );
  FA_X1 \mult_22/S2_23_49  ( .A(\mult_22/ab[23][49] ), .B(
        \mult_22/CARRYB[22][49] ), .CI(\mult_22/SUMB[22][50] ), .CO(
        \mult_22/CARRYB[23][49] ), .S(\mult_22/SUMB[23][49] ) );
  FA_X1 \mult_22/S2_23_48  ( .A(\mult_22/ab[23][48] ), .B(
        \mult_22/CARRYB[22][48] ), .CI(\mult_22/SUMB[22][49] ), .CO(
        \mult_22/CARRYB[23][48] ), .S(\mult_22/SUMB[23][48] ) );
  FA_X1 \mult_22/S2_23_47  ( .A(\mult_22/ab[23][47] ), .B(
        \mult_22/CARRYB[22][47] ), .CI(\mult_22/SUMB[22][48] ), .CO(
        \mult_22/CARRYB[23][47] ), .S(\mult_22/SUMB[23][47] ) );
  FA_X1 \mult_22/S2_23_46  ( .A(\mult_22/ab[23][46] ), .B(
        \mult_22/CARRYB[22][46] ), .CI(\mult_22/SUMB[22][47] ), .CO(
        \mult_22/CARRYB[23][46] ), .S(\mult_22/SUMB[23][46] ) );
  FA_X1 \mult_22/S2_23_45  ( .A(\mult_22/ab[23][45] ), .B(
        \mult_22/CARRYB[22][45] ), .CI(\mult_22/SUMB[22][46] ), .CO(
        \mult_22/CARRYB[23][45] ), .S(\mult_22/SUMB[23][45] ) );
  FA_X1 \mult_22/S2_23_44  ( .A(\mult_22/CARRYB[22][44] ), .B(
        \mult_22/ab[23][44] ), .CI(\mult_22/SUMB[22][45] ), .CO(
        \mult_22/CARRYB[23][44] ), .S(\mult_22/SUMB[23][44] ) );
  FA_X1 \mult_22/S2_23_43  ( .A(\mult_22/ab[23][43] ), .B(
        \mult_22/CARRYB[22][43] ), .CI(\mult_22/SUMB[22][44] ), .CO(
        \mult_22/CARRYB[23][43] ), .S(\mult_22/SUMB[23][43] ) );
  FA_X1 \mult_22/S2_23_42  ( .A(\mult_22/ab[23][42] ), .B(
        \mult_22/CARRYB[22][42] ), .CI(\mult_22/SUMB[22][43] ), .CO(
        \mult_22/CARRYB[23][42] ), .S(\mult_22/SUMB[23][42] ) );
  FA_X1 \mult_22/S2_23_41  ( .A(\mult_22/CARRYB[22][41] ), .B(
        \mult_22/ab[23][41] ), .CI(\mult_22/SUMB[22][42] ), .CO(
        \mult_22/CARRYB[23][41] ), .S(\mult_22/SUMB[23][41] ) );
  FA_X1 \mult_22/S2_23_40  ( .A(\mult_22/ab[23][40] ), .B(
        \mult_22/CARRYB[22][40] ), .CI(\mult_22/SUMB[22][41] ), .CO(
        \mult_22/CARRYB[23][40] ), .S(\mult_22/SUMB[23][40] ) );
  FA_X1 \mult_22/S2_23_39  ( .A(\mult_22/ab[23][39] ), .B(
        \mult_22/CARRYB[22][39] ), .CI(\mult_22/SUMB[22][40] ), .CO(
        \mult_22/CARRYB[23][39] ), .S(\mult_22/SUMB[23][39] ) );
  FA_X1 \mult_22/S2_23_38  ( .A(\mult_22/SUMB[22][39] ), .B(
        \mult_22/ab[23][38] ), .CI(\mult_22/CARRYB[22][38] ), .CO(
        \mult_22/CARRYB[23][38] ), .S(\mult_22/SUMB[23][38] ) );
  FA_X1 \mult_22/S2_23_36  ( .A(\mult_22/ab[23][36] ), .B(
        \mult_22/CARRYB[22][36] ), .CI(\mult_22/SUMB[22][37] ), .CO(
        \mult_22/CARRYB[23][36] ), .S(\mult_22/SUMB[23][36] ) );
  FA_X1 \mult_22/S2_23_35  ( .A(\mult_22/ab[23][35] ), .B(
        \mult_22/CARRYB[22][35] ), .CI(\mult_22/SUMB[22][36] ), .CO(
        \mult_22/CARRYB[23][35] ), .S(\mult_22/SUMB[23][35] ) );
  FA_X1 \mult_22/S2_23_34  ( .A(\mult_22/ab[23][34] ), .B(
        \mult_22/CARRYB[22][34] ), .CI(\mult_22/SUMB[22][35] ), .CO(
        \mult_22/CARRYB[23][34] ), .S(\mult_22/SUMB[23][34] ) );
  FA_X1 \mult_22/S2_23_33  ( .A(\mult_22/ab[23][33] ), .B(
        \mult_22/CARRYB[22][33] ), .CI(\mult_22/SUMB[22][34] ), .CO(
        \mult_22/CARRYB[23][33] ), .S(\mult_22/SUMB[23][33] ) );
  FA_X1 \mult_22/S2_23_32  ( .A(\mult_22/ab[23][32] ), .B(
        \mult_22/CARRYB[22][32] ), .CI(\mult_22/SUMB[22][33] ), .CO(
        \mult_22/CARRYB[23][32] ), .S(\mult_22/SUMB[23][32] ) );
  FA_X1 \mult_22/S2_23_31  ( .A(\mult_22/ab[23][31] ), .B(
        \mult_22/CARRYB[22][31] ), .CI(\mult_22/SUMB[22][32] ), .CO(
        \mult_22/CARRYB[23][31] ), .S(\mult_22/SUMB[23][31] ) );
  FA_X1 \mult_22/S2_23_30  ( .A(\mult_22/ab[23][30] ), .B(
        \mult_22/CARRYB[22][30] ), .CI(\mult_22/SUMB[22][31] ), .CO(
        \mult_22/CARRYB[23][30] ), .S(\mult_22/SUMB[23][30] ) );
  FA_X1 \mult_22/S2_23_29  ( .A(\mult_22/ab[23][29] ), .B(
        \mult_22/CARRYB[22][29] ), .CI(\mult_22/SUMB[22][30] ), .CO(
        \mult_22/CARRYB[23][29] ), .S(\mult_22/SUMB[23][29] ) );
  FA_X1 \mult_22/S2_23_28  ( .A(\mult_22/ab[23][28] ), .B(
        \mult_22/CARRYB[22][28] ), .CI(\mult_22/SUMB[22][29] ), .CO(
        \mult_22/CARRYB[23][28] ), .S(\mult_22/SUMB[23][28] ) );
  FA_X1 \mult_22/S2_23_27  ( .A(\mult_22/ab[23][27] ), .B(
        \mult_22/CARRYB[22][27] ), .CI(\mult_22/SUMB[22][28] ), .CO(
        \mult_22/CARRYB[23][27] ), .S(\mult_22/SUMB[23][27] ) );
  FA_X1 \mult_22/S2_23_26  ( .A(\mult_22/ab[23][26] ), .B(
        \mult_22/CARRYB[22][26] ), .CI(\mult_22/SUMB[22][27] ), .CO(
        \mult_22/CARRYB[23][26] ), .S(\mult_22/SUMB[23][26] ) );
  FA_X1 \mult_22/S2_23_25  ( .A(\mult_22/ab[23][25] ), .B(
        \mult_22/CARRYB[22][25] ), .CI(\mult_22/SUMB[22][26] ), .CO(
        \mult_22/CARRYB[23][25] ), .S(\mult_22/SUMB[23][25] ) );
  FA_X1 \mult_22/S2_23_24  ( .A(\mult_22/ab[23][24] ), .B(
        \mult_22/CARRYB[22][24] ), .CI(\mult_22/SUMB[22][25] ), .CO(
        \mult_22/CARRYB[23][24] ), .S(\mult_22/SUMB[23][24] ) );
  FA_X1 \mult_22/S2_23_23  ( .A(\mult_22/ab[23][23] ), .B(
        \mult_22/CARRYB[22][23] ), .CI(\mult_22/SUMB[22][24] ), .CO(
        \mult_22/CARRYB[23][23] ), .S(\mult_22/SUMB[23][23] ) );
  FA_X1 \mult_22/S2_23_22  ( .A(\mult_22/ab[23][22] ), .B(
        \mult_22/CARRYB[22][22] ), .CI(\mult_22/SUMB[22][23] ), .CO(
        \mult_22/CARRYB[23][22] ), .S(\mult_22/SUMB[23][22] ) );
  FA_X1 \mult_22/S2_23_21  ( .A(\mult_22/ab[23][21] ), .B(
        \mult_22/CARRYB[22][21] ), .CI(\mult_22/SUMB[22][22] ), .CO(
        \mult_22/CARRYB[23][21] ), .S(\mult_22/SUMB[23][21] ) );
  FA_X1 \mult_22/S2_23_20  ( .A(\mult_22/ab[23][20] ), .B(
        \mult_22/CARRYB[22][20] ), .CI(\mult_22/SUMB[22][21] ), .CO(
        \mult_22/CARRYB[23][20] ), .S(\mult_22/SUMB[23][20] ) );
  FA_X1 \mult_22/S2_23_19  ( .A(\mult_22/ab[23][19] ), .B(
        \mult_22/CARRYB[22][19] ), .CI(\mult_22/SUMB[22][20] ), .CO(
        \mult_22/CARRYB[23][19] ), .S(\mult_22/SUMB[23][19] ) );
  FA_X1 \mult_22/S2_23_18  ( .A(\mult_22/ab[23][18] ), .B(
        \mult_22/CARRYB[22][18] ), .CI(\mult_22/SUMB[22][19] ), .CO(
        \mult_22/CARRYB[23][18] ), .S(\mult_22/SUMB[23][18] ) );
  FA_X1 \mult_22/S2_23_17  ( .A(\mult_22/ab[23][17] ), .B(
        \mult_22/CARRYB[22][17] ), .CI(\mult_22/SUMB[22][18] ), .CO(
        \mult_22/CARRYB[23][17] ), .S(\mult_22/SUMB[23][17] ) );
  FA_X1 \mult_22/S2_23_16  ( .A(\mult_22/ab[23][16] ), .B(
        \mult_22/CARRYB[22][16] ), .CI(\mult_22/SUMB[22][17] ), .CO(
        \mult_22/CARRYB[23][16] ), .S(\mult_22/SUMB[23][16] ) );
  FA_X1 \mult_22/S2_23_15  ( .A(\mult_22/ab[23][15] ), .B(
        \mult_22/CARRYB[22][15] ), .CI(\mult_22/SUMB[22][16] ), .CO(
        \mult_22/CARRYB[23][15] ), .S(\mult_22/SUMB[23][15] ) );
  FA_X1 \mult_22/S2_23_14  ( .A(\mult_22/ab[23][14] ), .B(
        \mult_22/CARRYB[22][14] ), .CI(\mult_22/SUMB[22][15] ), .CO(
        \mult_22/CARRYB[23][14] ), .S(\mult_22/SUMB[23][14] ) );
  FA_X1 \mult_22/S2_23_13  ( .A(\mult_22/ab[23][13] ), .B(
        \mult_22/CARRYB[22][13] ), .CI(\mult_22/SUMB[22][14] ), .CO(
        \mult_22/CARRYB[23][13] ), .S(\mult_22/SUMB[23][13] ) );
  FA_X1 \mult_22/S2_23_12  ( .A(\mult_22/ab[23][12] ), .B(
        \mult_22/CARRYB[22][12] ), .CI(\mult_22/SUMB[22][13] ), .CO(
        \mult_22/CARRYB[23][12] ), .S(\mult_22/SUMB[23][12] ) );
  FA_X1 \mult_22/S2_23_11  ( .A(\mult_22/ab[23][11] ), .B(
        \mult_22/CARRYB[22][11] ), .CI(\mult_22/SUMB[22][12] ), .CO(
        \mult_22/CARRYB[23][11] ), .S(\mult_22/SUMB[23][11] ) );
  FA_X1 \mult_22/S2_23_10  ( .A(\mult_22/ab[23][10] ), .B(
        \mult_22/CARRYB[22][10] ), .CI(\mult_22/SUMB[22][11] ), .CO(
        \mult_22/CARRYB[23][10] ), .S(\mult_22/SUMB[23][10] ) );
  FA_X1 \mult_22/S2_23_9  ( .A(\mult_22/ab[23][9] ), .B(
        \mult_22/CARRYB[22][9] ), .CI(\mult_22/SUMB[22][10] ), .CO(
        \mult_22/CARRYB[23][9] ), .S(\mult_22/SUMB[23][9] ) );
  FA_X1 \mult_22/S2_23_8  ( .A(\mult_22/ab[23][8] ), .B(
        \mult_22/CARRYB[22][8] ), .CI(\mult_22/SUMB[22][9] ), .CO(
        \mult_22/CARRYB[23][8] ), .S(\mult_22/SUMB[23][8] ) );
  FA_X1 \mult_22/S2_23_7  ( .A(\mult_22/ab[23][7] ), .B(
        \mult_22/CARRYB[22][7] ), .CI(\mult_22/SUMB[22][8] ), .CO(
        \mult_22/CARRYB[23][7] ), .S(\mult_22/SUMB[23][7] ) );
  FA_X1 \mult_22/S2_23_6  ( .A(\mult_22/ab[23][6] ), .B(
        \mult_22/CARRYB[22][6] ), .CI(\mult_22/SUMB[22][7] ), .CO(
        \mult_22/CARRYB[23][6] ), .S(\mult_22/SUMB[23][6] ) );
  FA_X1 \mult_22/S2_23_5  ( .A(\mult_22/ab[23][5] ), .B(
        \mult_22/CARRYB[22][5] ), .CI(\mult_22/SUMB[22][6] ), .CO(
        \mult_22/CARRYB[23][5] ), .S(\mult_22/SUMB[23][5] ) );
  FA_X1 \mult_22/S2_23_4  ( .A(\mult_22/ab[23][4] ), .B(
        \mult_22/CARRYB[22][4] ), .CI(\mult_22/SUMB[22][5] ), .CO(
        \mult_22/CARRYB[23][4] ), .S(\mult_22/SUMB[23][4] ) );
  FA_X1 \mult_22/S2_23_3  ( .A(\mult_22/ab[23][3] ), .B(
        \mult_22/CARRYB[22][3] ), .CI(\mult_22/SUMB[22][4] ), .CO(
        \mult_22/CARRYB[23][3] ), .S(\mult_22/SUMB[23][3] ) );
  FA_X1 \mult_22/S2_23_2  ( .A(\mult_22/ab[23][2] ), .B(
        \mult_22/CARRYB[22][2] ), .CI(\mult_22/SUMB[22][3] ), .CO(
        \mult_22/CARRYB[23][2] ), .S(\mult_22/SUMB[23][2] ) );
  FA_X1 \mult_22/S2_23_1  ( .A(\mult_22/ab[23][1] ), .B(
        \mult_22/CARRYB[22][1] ), .CI(\mult_22/SUMB[22][2] ), .CO(
        \mult_22/CARRYB[23][1] ), .S(\mult_22/SUMB[23][1] ) );
  FA_X1 \mult_22/S1_23_0  ( .A(\mult_22/ab[23][0] ), .B(
        \mult_22/CARRYB[22][0] ), .CI(\mult_22/SUMB[22][1] ), .CO(
        \mult_22/CARRYB[23][0] ), .S(N151) );
  FA_X1 \mult_22/S3_24_62  ( .A(\mult_22/ab[24][62] ), .B(
        \mult_22/CARRYB[23][62] ), .CI(\mult_22/ab[23][63] ), .CO(
        \mult_22/CARRYB[24][62] ), .S(\mult_22/SUMB[24][62] ) );
  FA_X1 \mult_22/S2_24_61  ( .A(\mult_22/ab[24][61] ), .B(
        \mult_22/CARRYB[23][61] ), .CI(\mult_22/SUMB[23][62] ), .CO(
        \mult_22/CARRYB[24][61] ), .S(\mult_22/SUMB[24][61] ) );
  FA_X1 \mult_22/S2_24_60  ( .A(\mult_22/ab[24][60] ), .B(
        \mult_22/CARRYB[23][60] ), .CI(\mult_22/SUMB[23][61] ), .CO(
        \mult_22/CARRYB[24][60] ), .S(\mult_22/SUMB[24][60] ) );
  FA_X1 \mult_22/S2_24_59  ( .A(\mult_22/ab[24][59] ), .B(
        \mult_22/CARRYB[23][59] ), .CI(\mult_22/SUMB[23][60] ), .CO(
        \mult_22/CARRYB[24][59] ), .S(\mult_22/SUMB[24][59] ) );
  FA_X1 \mult_22/S2_24_58  ( .A(\mult_22/ab[24][58] ), .B(
        \mult_22/CARRYB[23][58] ), .CI(\mult_22/SUMB[23][59] ), .CO(
        \mult_22/CARRYB[24][58] ), .S(\mult_22/SUMB[24][58] ) );
  FA_X1 \mult_22/S2_24_57  ( .A(\mult_22/ab[24][57] ), .B(
        \mult_22/CARRYB[23][57] ), .CI(\mult_22/SUMB[23][58] ), .CO(
        \mult_22/CARRYB[24][57] ), .S(\mult_22/SUMB[24][57] ) );
  FA_X1 \mult_22/S2_24_56  ( .A(\mult_22/ab[24][56] ), .B(
        \mult_22/CARRYB[23][56] ), .CI(\mult_22/SUMB[23][57] ), .CO(
        \mult_22/CARRYB[24][56] ), .S(\mult_22/SUMB[24][56] ) );
  FA_X1 \mult_22/S2_24_55  ( .A(\mult_22/ab[24][55] ), .B(
        \mult_22/CARRYB[23][55] ), .CI(\mult_22/SUMB[23][56] ), .CO(
        \mult_22/CARRYB[24][55] ), .S(\mult_22/SUMB[24][55] ) );
  FA_X1 \mult_22/S2_24_54  ( .A(\mult_22/ab[24][54] ), .B(
        \mult_22/CARRYB[23][54] ), .CI(\mult_22/SUMB[23][55] ), .CO(
        \mult_22/CARRYB[24][54] ), .S(\mult_22/SUMB[24][54] ) );
  FA_X1 \mult_22/S2_24_53  ( .A(\mult_22/ab[24][53] ), .B(
        \mult_22/CARRYB[23][53] ), .CI(\mult_22/SUMB[23][54] ), .CO(
        \mult_22/CARRYB[24][53] ), .S(\mult_22/SUMB[24][53] ) );
  FA_X1 \mult_22/S2_24_52  ( .A(\mult_22/ab[24][52] ), .B(
        \mult_22/CARRYB[23][52] ), .CI(\mult_22/SUMB[23][53] ), .CO(
        \mult_22/CARRYB[24][52] ), .S(\mult_22/SUMB[24][52] ) );
  FA_X1 \mult_22/S2_24_51  ( .A(\mult_22/ab[24][51] ), .B(
        \mult_22/CARRYB[23][51] ), .CI(\mult_22/SUMB[23][52] ), .CO(
        \mult_22/CARRYB[24][51] ), .S(\mult_22/SUMB[24][51] ) );
  FA_X1 \mult_22/S2_24_50  ( .A(\mult_22/ab[24][50] ), .B(
        \mult_22/CARRYB[23][50] ), .CI(\mult_22/SUMB[23][51] ), .CO(
        \mult_22/CARRYB[24][50] ), .S(\mult_22/SUMB[24][50] ) );
  FA_X1 \mult_22/S2_24_49  ( .A(\mult_22/ab[24][49] ), .B(
        \mult_22/CARRYB[23][49] ), .CI(\mult_22/SUMB[23][50] ), .CO(
        \mult_22/CARRYB[24][49] ), .S(\mult_22/SUMB[24][49] ) );
  FA_X1 \mult_22/S2_24_48  ( .A(\mult_22/ab[24][48] ), .B(
        \mult_22/CARRYB[23][48] ), .CI(\mult_22/SUMB[23][49] ), .CO(
        \mult_22/CARRYB[24][48] ), .S(\mult_22/SUMB[24][48] ) );
  FA_X1 \mult_22/S2_24_47  ( .A(\mult_22/ab[24][47] ), .B(
        \mult_22/CARRYB[23][47] ), .CI(\mult_22/SUMB[23][48] ), .CO(
        \mult_22/CARRYB[24][47] ), .S(\mult_22/SUMB[24][47] ) );
  FA_X1 \mult_22/S2_24_46  ( .A(\mult_22/ab[24][46] ), .B(
        \mult_22/CARRYB[23][46] ), .CI(\mult_22/SUMB[23][47] ), .CO(
        \mult_22/CARRYB[24][46] ), .S(\mult_22/SUMB[24][46] ) );
  FA_X1 \mult_22/S2_24_45  ( .A(\mult_22/ab[24][45] ), .B(
        \mult_22/CARRYB[23][45] ), .CI(\mult_22/SUMB[23][46] ), .CO(
        \mult_22/CARRYB[24][45] ), .S(\mult_22/SUMB[24][45] ) );
  FA_X1 \mult_22/S2_24_44  ( .A(\mult_22/ab[24][44] ), .B(
        \mult_22/CARRYB[23][44] ), .CI(\mult_22/SUMB[23][45] ), .CO(
        \mult_22/CARRYB[24][44] ), .S(\mult_22/SUMB[24][44] ) );
  FA_X1 \mult_22/S2_24_43  ( .A(\mult_22/ab[24][43] ), .B(
        \mult_22/CARRYB[23][43] ), .CI(\mult_22/SUMB[23][44] ), .CO(
        \mult_22/CARRYB[24][43] ), .S(\mult_22/SUMB[24][43] ) );
  FA_X1 \mult_22/S2_24_42  ( .A(\mult_22/CARRYB[23][42] ), .B(
        \mult_22/ab[24][42] ), .CI(\mult_22/SUMB[23][43] ), .CO(
        \mult_22/CARRYB[24][42] ), .S(\mult_22/SUMB[24][42] ) );
  FA_X1 \mult_22/S2_24_40  ( .A(\mult_22/ab[24][40] ), .B(
        \mult_22/CARRYB[23][40] ), .CI(\mult_22/SUMB[23][41] ), .CO(
        \mult_22/CARRYB[24][40] ), .S(\mult_22/SUMB[24][40] ) );
  FA_X1 \mult_22/S2_24_39  ( .A(\mult_22/ab[24][39] ), .B(
        \mult_22/CARRYB[23][39] ), .CI(\mult_22/SUMB[23][40] ), .CO(
        \mult_22/CARRYB[24][39] ), .S(\mult_22/SUMB[24][39] ) );
  FA_X1 \mult_22/S2_24_38  ( .A(\mult_22/ab[24][38] ), .B(
        \mult_22/CARRYB[23][38] ), .CI(\mult_22/SUMB[23][39] ), .CO(
        \mult_22/CARRYB[24][38] ), .S(\mult_22/SUMB[24][38] ) );
  FA_X1 \mult_22/S2_24_37  ( .A(\mult_22/ab[24][37] ), .B(
        \mult_22/CARRYB[23][37] ), .CI(\mult_22/SUMB[23][38] ), .CO(
        \mult_22/CARRYB[24][37] ), .S(\mult_22/SUMB[24][37] ) );
  FA_X1 \mult_22/S2_24_36  ( .A(\mult_22/ab[24][36] ), .B(
        \mult_22/CARRYB[23][36] ), .CI(\mult_22/SUMB[23][37] ), .CO(
        \mult_22/CARRYB[24][36] ), .S(\mult_22/SUMB[24][36] ) );
  FA_X1 \mult_22/S2_24_35  ( .A(\mult_22/ab[24][35] ), .B(
        \mult_22/CARRYB[23][35] ), .CI(\mult_22/SUMB[23][36] ), .CO(
        \mult_22/CARRYB[24][35] ), .S(\mult_22/SUMB[24][35] ) );
  FA_X1 \mult_22/S2_24_34  ( .A(\mult_22/ab[24][34] ), .B(
        \mult_22/CARRYB[23][34] ), .CI(\mult_22/SUMB[23][35] ), .CO(
        \mult_22/CARRYB[24][34] ), .S(\mult_22/SUMB[24][34] ) );
  FA_X1 \mult_22/S2_24_33  ( .A(\mult_22/ab[24][33] ), .B(
        \mult_22/CARRYB[23][33] ), .CI(\mult_22/SUMB[23][34] ), .CO(
        \mult_22/CARRYB[24][33] ), .S(\mult_22/SUMB[24][33] ) );
  FA_X1 \mult_22/S2_24_31  ( .A(\mult_22/ab[24][31] ), .B(
        \mult_22/CARRYB[23][31] ), .CI(\mult_22/SUMB[23][32] ), .CO(
        \mult_22/CARRYB[24][31] ), .S(\mult_22/SUMB[24][31] ) );
  FA_X1 \mult_22/S2_24_30  ( .A(\mult_22/ab[24][30] ), .B(
        \mult_22/CARRYB[23][30] ), .CI(\mult_22/SUMB[23][31] ), .CO(
        \mult_22/CARRYB[24][30] ), .S(\mult_22/SUMB[24][30] ) );
  FA_X1 \mult_22/S2_24_29  ( .A(\mult_22/ab[24][29] ), .B(
        \mult_22/CARRYB[23][29] ), .CI(\mult_22/SUMB[23][30] ), .CO(
        \mult_22/CARRYB[24][29] ), .S(\mult_22/SUMB[24][29] ) );
  FA_X1 \mult_22/S2_24_28  ( .A(\mult_22/ab[24][28] ), .B(
        \mult_22/CARRYB[23][28] ), .CI(\mult_22/SUMB[23][29] ), .CO(
        \mult_22/CARRYB[24][28] ), .S(\mult_22/SUMB[24][28] ) );
  FA_X1 \mult_22/S2_24_27  ( .A(\mult_22/ab[24][27] ), .B(
        \mult_22/CARRYB[23][27] ), .CI(\mult_22/SUMB[23][28] ), .CO(
        \mult_22/CARRYB[24][27] ), .S(\mult_22/SUMB[24][27] ) );
  FA_X1 \mult_22/S2_24_26  ( .A(\mult_22/ab[24][26] ), .B(
        \mult_22/CARRYB[23][26] ), .CI(\mult_22/SUMB[23][27] ), .CO(
        \mult_22/CARRYB[24][26] ), .S(\mult_22/SUMB[24][26] ) );
  FA_X1 \mult_22/S2_24_25  ( .A(\mult_22/ab[24][25] ), .B(
        \mult_22/CARRYB[23][25] ), .CI(\mult_22/SUMB[23][26] ), .CO(
        \mult_22/CARRYB[24][25] ), .S(\mult_22/SUMB[24][25] ) );
  FA_X1 \mult_22/S2_24_24  ( .A(\mult_22/ab[24][24] ), .B(
        \mult_22/CARRYB[23][24] ), .CI(\mult_22/SUMB[23][25] ), .CO(
        \mult_22/CARRYB[24][24] ), .S(\mult_22/SUMB[24][24] ) );
  FA_X1 \mult_22/S2_24_23  ( .A(\mult_22/ab[24][23] ), .B(
        \mult_22/CARRYB[23][23] ), .CI(\mult_22/SUMB[23][24] ), .CO(
        \mult_22/CARRYB[24][23] ), .S(\mult_22/SUMB[24][23] ) );
  FA_X1 \mult_22/S2_24_22  ( .A(\mult_22/ab[24][22] ), .B(
        \mult_22/CARRYB[23][22] ), .CI(\mult_22/SUMB[23][23] ), .CO(
        \mult_22/CARRYB[24][22] ), .S(\mult_22/SUMB[24][22] ) );
  FA_X1 \mult_22/S2_24_21  ( .A(\mult_22/ab[24][21] ), .B(
        \mult_22/CARRYB[23][21] ), .CI(\mult_22/SUMB[23][22] ), .CO(
        \mult_22/CARRYB[24][21] ), .S(\mult_22/SUMB[24][21] ) );
  FA_X1 \mult_22/S2_24_20  ( .A(\mult_22/ab[24][20] ), .B(
        \mult_22/CARRYB[23][20] ), .CI(\mult_22/SUMB[23][21] ), .CO(
        \mult_22/CARRYB[24][20] ), .S(\mult_22/SUMB[24][20] ) );
  FA_X1 \mult_22/S2_24_19  ( .A(\mult_22/ab[24][19] ), .B(
        \mult_22/CARRYB[23][19] ), .CI(\mult_22/SUMB[23][20] ), .CO(
        \mult_22/CARRYB[24][19] ), .S(\mult_22/SUMB[24][19] ) );
  FA_X1 \mult_22/S2_24_18  ( .A(\mult_22/ab[24][18] ), .B(
        \mult_22/CARRYB[23][18] ), .CI(\mult_22/SUMB[23][19] ), .CO(
        \mult_22/CARRYB[24][18] ), .S(\mult_22/SUMB[24][18] ) );
  FA_X1 \mult_22/S2_24_17  ( .A(\mult_22/ab[24][17] ), .B(
        \mult_22/CARRYB[23][17] ), .CI(\mult_22/SUMB[23][18] ), .CO(
        \mult_22/CARRYB[24][17] ), .S(\mult_22/SUMB[24][17] ) );
  FA_X1 \mult_22/S2_24_16  ( .A(\mult_22/ab[24][16] ), .B(
        \mult_22/CARRYB[23][16] ), .CI(\mult_22/SUMB[23][17] ), .CO(
        \mult_22/CARRYB[24][16] ), .S(\mult_22/SUMB[24][16] ) );
  FA_X1 \mult_22/S2_24_15  ( .A(\mult_22/ab[24][15] ), .B(
        \mult_22/CARRYB[23][15] ), .CI(\mult_22/SUMB[23][16] ), .CO(
        \mult_22/CARRYB[24][15] ), .S(\mult_22/SUMB[24][15] ) );
  FA_X1 \mult_22/S2_24_14  ( .A(\mult_22/ab[24][14] ), .B(
        \mult_22/CARRYB[23][14] ), .CI(\mult_22/SUMB[23][15] ), .CO(
        \mult_22/CARRYB[24][14] ), .S(\mult_22/SUMB[24][14] ) );
  FA_X1 \mult_22/S2_24_13  ( .A(\mult_22/ab[24][13] ), .B(
        \mult_22/CARRYB[23][13] ), .CI(\mult_22/SUMB[23][14] ), .CO(
        \mult_22/CARRYB[24][13] ), .S(\mult_22/SUMB[24][13] ) );
  FA_X1 \mult_22/S2_24_12  ( .A(\mult_22/ab[24][12] ), .B(
        \mult_22/CARRYB[23][12] ), .CI(\mult_22/SUMB[23][13] ), .CO(
        \mult_22/CARRYB[24][12] ), .S(\mult_22/SUMB[24][12] ) );
  FA_X1 \mult_22/S2_24_11  ( .A(\mult_22/ab[24][11] ), .B(
        \mult_22/CARRYB[23][11] ), .CI(\mult_22/SUMB[23][12] ), .CO(
        \mult_22/CARRYB[24][11] ), .S(\mult_22/SUMB[24][11] ) );
  FA_X1 \mult_22/S2_24_10  ( .A(\mult_22/ab[24][10] ), .B(
        \mult_22/CARRYB[23][10] ), .CI(\mult_22/SUMB[23][11] ), .CO(
        \mult_22/CARRYB[24][10] ), .S(\mult_22/SUMB[24][10] ) );
  FA_X1 \mult_22/S2_24_9  ( .A(\mult_22/ab[24][9] ), .B(
        \mult_22/CARRYB[23][9] ), .CI(\mult_22/SUMB[23][10] ), .CO(
        \mult_22/CARRYB[24][9] ), .S(\mult_22/SUMB[24][9] ) );
  FA_X1 \mult_22/S2_24_8  ( .A(\mult_22/ab[24][8] ), .B(
        \mult_22/CARRYB[23][8] ), .CI(\mult_22/SUMB[23][9] ), .CO(
        \mult_22/CARRYB[24][8] ), .S(\mult_22/SUMB[24][8] ) );
  FA_X1 \mult_22/S2_24_7  ( .A(\mult_22/ab[24][7] ), .B(
        \mult_22/CARRYB[23][7] ), .CI(\mult_22/SUMB[23][8] ), .CO(
        \mult_22/CARRYB[24][7] ), .S(\mult_22/SUMB[24][7] ) );
  FA_X1 \mult_22/S2_24_6  ( .A(\mult_22/ab[24][6] ), .B(
        \mult_22/CARRYB[23][6] ), .CI(\mult_22/SUMB[23][7] ), .CO(
        \mult_22/CARRYB[24][6] ), .S(\mult_22/SUMB[24][6] ) );
  FA_X1 \mult_22/S2_24_5  ( .A(\mult_22/ab[24][5] ), .B(
        \mult_22/CARRYB[23][5] ), .CI(\mult_22/SUMB[23][6] ), .CO(
        \mult_22/CARRYB[24][5] ), .S(\mult_22/SUMB[24][5] ) );
  FA_X1 \mult_22/S2_24_4  ( .A(\mult_22/ab[24][4] ), .B(
        \mult_22/CARRYB[23][4] ), .CI(\mult_22/SUMB[23][5] ), .CO(
        \mult_22/CARRYB[24][4] ), .S(\mult_22/SUMB[24][4] ) );
  FA_X1 \mult_22/S2_24_3  ( .A(\mult_22/ab[24][3] ), .B(
        \mult_22/CARRYB[23][3] ), .CI(\mult_22/SUMB[23][4] ), .CO(
        \mult_22/CARRYB[24][3] ), .S(\mult_22/SUMB[24][3] ) );
  FA_X1 \mult_22/S2_24_2  ( .A(\mult_22/ab[24][2] ), .B(
        \mult_22/CARRYB[23][2] ), .CI(\mult_22/SUMB[23][3] ), .CO(
        \mult_22/CARRYB[24][2] ), .S(\mult_22/SUMB[24][2] ) );
  FA_X1 \mult_22/S2_24_1  ( .A(\mult_22/ab[24][1] ), .B(
        \mult_22/CARRYB[23][1] ), .CI(\mult_22/SUMB[23][2] ), .CO(
        \mult_22/CARRYB[24][1] ), .S(\mult_22/SUMB[24][1] ) );
  FA_X1 \mult_22/S1_24_0  ( .A(\mult_22/ab[24][0] ), .B(
        \mult_22/CARRYB[23][0] ), .CI(\mult_22/SUMB[23][1] ), .CO(
        \mult_22/CARRYB[24][0] ), .S(N152) );
  FA_X1 \mult_22/S3_25_62  ( .A(\mult_22/ab[25][62] ), .B(
        \mult_22/CARRYB[24][62] ), .CI(\mult_22/ab[24][63] ), .CO(
        \mult_22/CARRYB[25][62] ), .S(\mult_22/SUMB[25][62] ) );
  FA_X1 \mult_22/S2_25_61  ( .A(\mult_22/ab[25][61] ), .B(
        \mult_22/CARRYB[24][61] ), .CI(\mult_22/SUMB[24][62] ), .CO(
        \mult_22/CARRYB[25][61] ), .S(\mult_22/SUMB[25][61] ) );
  FA_X1 \mult_22/S2_25_60  ( .A(\mult_22/ab[25][60] ), .B(
        \mult_22/CARRYB[24][60] ), .CI(\mult_22/SUMB[24][61] ), .CO(
        \mult_22/CARRYB[25][60] ), .S(\mult_22/SUMB[25][60] ) );
  FA_X1 \mult_22/S2_25_59  ( .A(\mult_22/ab[25][59] ), .B(
        \mult_22/CARRYB[24][59] ), .CI(\mult_22/SUMB[24][60] ), .CO(
        \mult_22/CARRYB[25][59] ), .S(\mult_22/SUMB[25][59] ) );
  FA_X1 \mult_22/S2_25_58  ( .A(\mult_22/ab[25][58] ), .B(
        \mult_22/CARRYB[24][58] ), .CI(\mult_22/SUMB[24][59] ), .CO(
        \mult_22/CARRYB[25][58] ), .S(\mult_22/SUMB[25][58] ) );
  FA_X1 \mult_22/S2_25_57  ( .A(\mult_22/ab[25][57] ), .B(
        \mult_22/CARRYB[24][57] ), .CI(\mult_22/SUMB[24][58] ), .CO(
        \mult_22/CARRYB[25][57] ), .S(\mult_22/SUMB[25][57] ) );
  FA_X1 \mult_22/S2_25_56  ( .A(\mult_22/ab[25][56] ), .B(
        \mult_22/CARRYB[24][56] ), .CI(\mult_22/SUMB[24][57] ), .CO(
        \mult_22/CARRYB[25][56] ), .S(\mult_22/SUMB[25][56] ) );
  FA_X1 \mult_22/S2_25_55  ( .A(\mult_22/ab[25][55] ), .B(
        \mult_22/CARRYB[24][55] ), .CI(\mult_22/SUMB[24][56] ), .CO(
        \mult_22/CARRYB[25][55] ), .S(\mult_22/SUMB[25][55] ) );
  FA_X1 \mult_22/S2_25_54  ( .A(\mult_22/ab[25][54] ), .B(
        \mult_22/CARRYB[24][54] ), .CI(\mult_22/SUMB[24][55] ), .CO(
        \mult_22/CARRYB[25][54] ), .S(\mult_22/SUMB[25][54] ) );
  FA_X1 \mult_22/S2_25_53  ( .A(\mult_22/ab[25][53] ), .B(
        \mult_22/CARRYB[24][53] ), .CI(\mult_22/SUMB[24][54] ), .CO(
        \mult_22/CARRYB[25][53] ), .S(\mult_22/SUMB[25][53] ) );
  FA_X1 \mult_22/S2_25_52  ( .A(\mult_22/ab[25][52] ), .B(
        \mult_22/CARRYB[24][52] ), .CI(\mult_22/SUMB[24][53] ), .CO(
        \mult_22/CARRYB[25][52] ), .S(\mult_22/SUMB[25][52] ) );
  FA_X1 \mult_22/S2_25_51  ( .A(\mult_22/ab[25][51] ), .B(
        \mult_22/CARRYB[24][51] ), .CI(\mult_22/SUMB[24][52] ), .CO(
        \mult_22/CARRYB[25][51] ), .S(\mult_22/SUMB[25][51] ) );
  FA_X1 \mult_22/S2_25_50  ( .A(\mult_22/ab[25][50] ), .B(
        \mult_22/CARRYB[24][50] ), .CI(\mult_22/SUMB[24][51] ), .CO(
        \mult_22/CARRYB[25][50] ), .S(\mult_22/SUMB[25][50] ) );
  FA_X1 \mult_22/S2_25_49  ( .A(\mult_22/ab[25][49] ), .B(
        \mult_22/CARRYB[24][49] ), .CI(\mult_22/SUMB[24][50] ), .CO(
        \mult_22/CARRYB[25][49] ), .S(\mult_22/SUMB[25][49] ) );
  FA_X1 \mult_22/S2_25_48  ( .A(\mult_22/ab[25][48] ), .B(
        \mult_22/CARRYB[24][48] ), .CI(\mult_22/SUMB[24][49] ), .CO(
        \mult_22/CARRYB[25][48] ), .S(\mult_22/SUMB[25][48] ) );
  FA_X1 \mult_22/S2_25_47  ( .A(\mult_22/ab[25][47] ), .B(
        \mult_22/CARRYB[24][47] ), .CI(\mult_22/SUMB[24][48] ), .CO(
        \mult_22/CARRYB[25][47] ), .S(\mult_22/SUMB[25][47] ) );
  FA_X1 \mult_22/S2_25_46  ( .A(\mult_22/ab[25][46] ), .B(
        \mult_22/CARRYB[24][46] ), .CI(\mult_22/SUMB[24][47] ), .CO(
        \mult_22/CARRYB[25][46] ), .S(\mult_22/SUMB[25][46] ) );
  FA_X1 \mult_22/S2_25_45  ( .A(\mult_22/ab[25][45] ), .B(
        \mult_22/CARRYB[24][45] ), .CI(\mult_22/SUMB[24][46] ), .CO(
        \mult_22/CARRYB[25][45] ), .S(\mult_22/SUMB[25][45] ) );
  FA_X1 \mult_22/S2_25_44  ( .A(\mult_22/ab[25][44] ), .B(
        \mult_22/CARRYB[24][44] ), .CI(\mult_22/SUMB[24][45] ), .CO(
        \mult_22/CARRYB[25][44] ), .S(\mult_22/SUMB[25][44] ) );
  FA_X1 \mult_22/S2_25_43  ( .A(\mult_22/ab[25][43] ), .B(
        \mult_22/CARRYB[24][43] ), .CI(\mult_22/SUMB[24][44] ), .CO(
        \mult_22/CARRYB[25][43] ), .S(\mult_22/SUMB[25][43] ) );
  FA_X1 \mult_22/S2_25_42  ( .A(\mult_22/CARRYB[24][42] ), .B(
        \mult_22/ab[25][42] ), .CI(\mult_22/SUMB[24][43] ), .CO(
        \mult_22/CARRYB[25][42] ), .S(\mult_22/SUMB[25][42] ) );
  FA_X1 \mult_22/S2_25_41  ( .A(\mult_22/ab[25][41] ), .B(
        \mult_22/CARRYB[24][41] ), .CI(\mult_22/SUMB[24][42] ), .CO(
        \mult_22/CARRYB[25][41] ), .S(\mult_22/SUMB[25][41] ) );
  FA_X1 \mult_22/S2_25_40  ( .A(\mult_22/ab[25][40] ), .B(
        \mult_22/CARRYB[24][40] ), .CI(\mult_22/SUMB[24][41] ), .CO(
        \mult_22/CARRYB[25][40] ), .S(\mult_22/SUMB[25][40] ) );
  FA_X1 \mult_22/S2_25_39  ( .A(\mult_22/CARRYB[24][39] ), .B(
        \mult_22/ab[25][39] ), .CI(\mult_22/SUMB[24][40] ), .CO(
        \mult_22/CARRYB[25][39] ), .S(\mult_22/SUMB[25][39] ) );
  FA_X1 \mult_22/S2_25_38  ( .A(\mult_22/ab[25][38] ), .B(
        \mult_22/CARRYB[24][38] ), .CI(\mult_22/SUMB[24][39] ), .CO(
        \mult_22/CARRYB[25][38] ), .S(\mult_22/SUMB[25][38] ) );
  FA_X1 \mult_22/S2_25_37  ( .A(\mult_22/ab[25][37] ), .B(
        \mult_22/CARRYB[24][37] ), .CI(\mult_22/SUMB[24][38] ), .CO(
        \mult_22/CARRYB[25][37] ), .S(\mult_22/SUMB[25][37] ) );
  FA_X1 \mult_22/S2_25_36  ( .A(\mult_22/ab[25][36] ), .B(
        \mult_22/CARRYB[24][36] ), .CI(\mult_22/SUMB[24][37] ), .CO(
        \mult_22/CARRYB[25][36] ), .S(\mult_22/SUMB[25][36] ) );
  FA_X1 \mult_22/S2_25_34  ( .A(\mult_22/ab[25][34] ), .B(
        \mult_22/CARRYB[24][34] ), .CI(\mult_22/SUMB[24][35] ), .CO(
        \mult_22/CARRYB[25][34] ), .S(\mult_22/SUMB[25][34] ) );
  FA_X1 \mult_22/S2_25_33  ( .A(\mult_22/ab[25][33] ), .B(
        \mult_22/CARRYB[24][33] ), .CI(\mult_22/SUMB[24][34] ), .CO(
        \mult_22/CARRYB[25][33] ), .S(\mult_22/SUMB[25][33] ) );
  FA_X1 \mult_22/S2_25_32  ( .A(\mult_22/ab[25][32] ), .B(
        \mult_22/CARRYB[24][32] ), .CI(\mult_22/SUMB[24][33] ), .CO(
        \mult_22/CARRYB[25][32] ), .S(\mult_22/SUMB[25][32] ) );
  FA_X1 \mult_22/S2_25_31  ( .A(\mult_22/ab[25][31] ), .B(
        \mult_22/CARRYB[24][31] ), .CI(\mult_22/SUMB[24][32] ), .CO(
        \mult_22/CARRYB[25][31] ), .S(\mult_22/SUMB[25][31] ) );
  FA_X1 \mult_22/S2_25_30  ( .A(\mult_22/ab[25][30] ), .B(
        \mult_22/CARRYB[24][30] ), .CI(\mult_22/SUMB[24][31] ), .CO(
        \mult_22/CARRYB[25][30] ), .S(\mult_22/SUMB[25][30] ) );
  FA_X1 \mult_22/S2_25_29  ( .A(\mult_22/ab[25][29] ), .B(
        \mult_22/CARRYB[24][29] ), .CI(\mult_22/SUMB[24][30] ), .CO(
        \mult_22/CARRYB[25][29] ), .S(\mult_22/SUMB[25][29] ) );
  FA_X1 \mult_22/S2_25_28  ( .A(\mult_22/ab[25][28] ), .B(
        \mult_22/CARRYB[24][28] ), .CI(\mult_22/SUMB[24][29] ), .CO(
        \mult_22/CARRYB[25][28] ), .S(\mult_22/SUMB[25][28] ) );
  FA_X1 \mult_22/S2_25_27  ( .A(\mult_22/ab[25][27] ), .B(
        \mult_22/CARRYB[24][27] ), .CI(\mult_22/SUMB[24][28] ), .CO(
        \mult_22/CARRYB[25][27] ), .S(\mult_22/SUMB[25][27] ) );
  FA_X1 \mult_22/S2_25_26  ( .A(\mult_22/ab[25][26] ), .B(
        \mult_22/CARRYB[24][26] ), .CI(\mult_22/SUMB[24][27] ), .CO(
        \mult_22/CARRYB[25][26] ), .S(\mult_22/SUMB[25][26] ) );
  FA_X1 \mult_22/S2_25_25  ( .A(\mult_22/ab[25][25] ), .B(
        \mult_22/CARRYB[24][25] ), .CI(\mult_22/SUMB[24][26] ), .CO(
        \mult_22/CARRYB[25][25] ), .S(\mult_22/SUMB[25][25] ) );
  FA_X1 \mult_22/S2_25_24  ( .A(\mult_22/ab[25][24] ), .B(
        \mult_22/CARRYB[24][24] ), .CI(\mult_22/SUMB[24][25] ), .CO(
        \mult_22/CARRYB[25][24] ), .S(\mult_22/SUMB[25][24] ) );
  FA_X1 \mult_22/S2_25_23  ( .A(\mult_22/ab[25][23] ), .B(
        \mult_22/CARRYB[24][23] ), .CI(\mult_22/SUMB[24][24] ), .CO(
        \mult_22/CARRYB[25][23] ), .S(\mult_22/SUMB[25][23] ) );
  FA_X1 \mult_22/S2_25_22  ( .A(\mult_22/ab[25][22] ), .B(
        \mult_22/CARRYB[24][22] ), .CI(\mult_22/SUMB[24][23] ), .CO(
        \mult_22/CARRYB[25][22] ), .S(\mult_22/SUMB[25][22] ) );
  FA_X1 \mult_22/S2_25_21  ( .A(\mult_22/ab[25][21] ), .B(
        \mult_22/CARRYB[24][21] ), .CI(\mult_22/SUMB[24][22] ), .CO(
        \mult_22/CARRYB[25][21] ), .S(\mult_22/SUMB[25][21] ) );
  FA_X1 \mult_22/S2_25_20  ( .A(\mult_22/ab[25][20] ), .B(
        \mult_22/CARRYB[24][20] ), .CI(\mult_22/SUMB[24][21] ), .CO(
        \mult_22/CARRYB[25][20] ), .S(\mult_22/SUMB[25][20] ) );
  FA_X1 \mult_22/S2_25_19  ( .A(\mult_22/ab[25][19] ), .B(
        \mult_22/CARRYB[24][19] ), .CI(\mult_22/SUMB[24][20] ), .CO(
        \mult_22/CARRYB[25][19] ), .S(\mult_22/SUMB[25][19] ) );
  FA_X1 \mult_22/S2_25_18  ( .A(\mult_22/ab[25][18] ), .B(
        \mult_22/CARRYB[24][18] ), .CI(\mult_22/SUMB[24][19] ), .CO(
        \mult_22/CARRYB[25][18] ), .S(\mult_22/SUMB[25][18] ) );
  FA_X1 \mult_22/S2_25_17  ( .A(\mult_22/ab[25][17] ), .B(
        \mult_22/CARRYB[24][17] ), .CI(\mult_22/SUMB[24][18] ), .CO(
        \mult_22/CARRYB[25][17] ), .S(\mult_22/SUMB[25][17] ) );
  FA_X1 \mult_22/S2_25_16  ( .A(\mult_22/ab[25][16] ), .B(
        \mult_22/CARRYB[24][16] ), .CI(\mult_22/SUMB[24][17] ), .CO(
        \mult_22/CARRYB[25][16] ), .S(\mult_22/SUMB[25][16] ) );
  FA_X1 \mult_22/S2_25_15  ( .A(\mult_22/ab[25][15] ), .B(
        \mult_22/CARRYB[24][15] ), .CI(\mult_22/SUMB[24][16] ), .CO(
        \mult_22/CARRYB[25][15] ), .S(\mult_22/SUMB[25][15] ) );
  FA_X1 \mult_22/S2_25_14  ( .A(\mult_22/ab[25][14] ), .B(
        \mult_22/CARRYB[24][14] ), .CI(\mult_22/SUMB[24][15] ), .CO(
        \mult_22/CARRYB[25][14] ), .S(\mult_22/SUMB[25][14] ) );
  FA_X1 \mult_22/S2_25_13  ( .A(\mult_22/ab[25][13] ), .B(
        \mult_22/CARRYB[24][13] ), .CI(\mult_22/SUMB[24][14] ), .CO(
        \mult_22/CARRYB[25][13] ), .S(\mult_22/SUMB[25][13] ) );
  FA_X1 \mult_22/S2_25_12  ( .A(\mult_22/ab[25][12] ), .B(
        \mult_22/CARRYB[24][12] ), .CI(\mult_22/SUMB[24][13] ), .CO(
        \mult_22/CARRYB[25][12] ), .S(\mult_22/SUMB[25][12] ) );
  FA_X1 \mult_22/S2_25_11  ( .A(\mult_22/ab[25][11] ), .B(
        \mult_22/CARRYB[24][11] ), .CI(\mult_22/SUMB[24][12] ), .CO(
        \mult_22/CARRYB[25][11] ), .S(\mult_22/SUMB[25][11] ) );
  FA_X1 \mult_22/S2_25_10  ( .A(\mult_22/ab[25][10] ), .B(
        \mult_22/CARRYB[24][10] ), .CI(\mult_22/SUMB[24][11] ), .CO(
        \mult_22/CARRYB[25][10] ), .S(\mult_22/SUMB[25][10] ) );
  FA_X1 \mult_22/S2_25_9  ( .A(\mult_22/ab[25][9] ), .B(
        \mult_22/CARRYB[24][9] ), .CI(\mult_22/SUMB[24][10] ), .CO(
        \mult_22/CARRYB[25][9] ), .S(\mult_22/SUMB[25][9] ) );
  FA_X1 \mult_22/S2_25_8  ( .A(\mult_22/ab[25][8] ), .B(
        \mult_22/CARRYB[24][8] ), .CI(\mult_22/SUMB[24][9] ), .CO(
        \mult_22/CARRYB[25][8] ), .S(\mult_22/SUMB[25][8] ) );
  FA_X1 \mult_22/S2_25_7  ( .A(\mult_22/ab[25][7] ), .B(
        \mult_22/CARRYB[24][7] ), .CI(\mult_22/SUMB[24][8] ), .CO(
        \mult_22/CARRYB[25][7] ), .S(\mult_22/SUMB[25][7] ) );
  FA_X1 \mult_22/S2_25_6  ( .A(\mult_22/ab[25][6] ), .B(
        \mult_22/CARRYB[24][6] ), .CI(\mult_22/SUMB[24][7] ), .CO(
        \mult_22/CARRYB[25][6] ), .S(\mult_22/SUMB[25][6] ) );
  FA_X1 \mult_22/S2_25_5  ( .A(\mult_22/ab[25][5] ), .B(
        \mult_22/CARRYB[24][5] ), .CI(\mult_22/SUMB[24][6] ), .CO(
        \mult_22/CARRYB[25][5] ), .S(\mult_22/SUMB[25][5] ) );
  FA_X1 \mult_22/S2_25_4  ( .A(\mult_22/ab[25][4] ), .B(
        \mult_22/CARRYB[24][4] ), .CI(\mult_22/SUMB[24][5] ), .CO(
        \mult_22/CARRYB[25][4] ), .S(\mult_22/SUMB[25][4] ) );
  FA_X1 \mult_22/S2_25_3  ( .A(\mult_22/ab[25][3] ), .B(
        \mult_22/CARRYB[24][3] ), .CI(\mult_22/SUMB[24][4] ), .CO(
        \mult_22/CARRYB[25][3] ), .S(\mult_22/SUMB[25][3] ) );
  FA_X1 \mult_22/S2_25_2  ( .A(\mult_22/ab[25][2] ), .B(
        \mult_22/CARRYB[24][2] ), .CI(\mult_22/SUMB[24][3] ), .CO(
        \mult_22/CARRYB[25][2] ), .S(\mult_22/SUMB[25][2] ) );
  FA_X1 \mult_22/S2_25_1  ( .A(\mult_22/ab[25][1] ), .B(
        \mult_22/CARRYB[24][1] ), .CI(\mult_22/SUMB[24][2] ), .CO(
        \mult_22/CARRYB[25][1] ), .S(\mult_22/SUMB[25][1] ) );
  FA_X1 \mult_22/S1_25_0  ( .A(\mult_22/ab[25][0] ), .B(
        \mult_22/CARRYB[24][0] ), .CI(\mult_22/SUMB[24][1] ), .CO(
        \mult_22/CARRYB[25][0] ), .S(N153) );
  FA_X1 \mult_22/S3_26_62  ( .A(\mult_22/ab[26][62] ), .B(
        \mult_22/CARRYB[25][62] ), .CI(\mult_22/ab[25][63] ), .CO(
        \mult_22/CARRYB[26][62] ), .S(\mult_22/SUMB[26][62] ) );
  FA_X1 \mult_22/S2_26_61  ( .A(\mult_22/ab[26][61] ), .B(
        \mult_22/CARRYB[25][61] ), .CI(\mult_22/SUMB[25][62] ), .CO(
        \mult_22/CARRYB[26][61] ), .S(\mult_22/SUMB[26][61] ) );
  FA_X1 \mult_22/S2_26_60  ( .A(\mult_22/ab[26][60] ), .B(
        \mult_22/CARRYB[25][60] ), .CI(\mult_22/SUMB[25][61] ), .CO(
        \mult_22/CARRYB[26][60] ), .S(\mult_22/SUMB[26][60] ) );
  FA_X1 \mult_22/S2_26_59  ( .A(\mult_22/ab[26][59] ), .B(
        \mult_22/CARRYB[25][59] ), .CI(\mult_22/SUMB[25][60] ), .CO(
        \mult_22/CARRYB[26][59] ), .S(\mult_22/SUMB[26][59] ) );
  FA_X1 \mult_22/S2_26_58  ( .A(\mult_22/ab[26][58] ), .B(
        \mult_22/CARRYB[25][58] ), .CI(\mult_22/SUMB[25][59] ), .CO(
        \mult_22/CARRYB[26][58] ), .S(\mult_22/SUMB[26][58] ) );
  FA_X1 \mult_22/S2_26_57  ( .A(\mult_22/ab[26][57] ), .B(
        \mult_22/CARRYB[25][57] ), .CI(\mult_22/SUMB[25][58] ), .CO(
        \mult_22/CARRYB[26][57] ), .S(\mult_22/SUMB[26][57] ) );
  FA_X1 \mult_22/S2_26_56  ( .A(\mult_22/ab[26][56] ), .B(
        \mult_22/CARRYB[25][56] ), .CI(\mult_22/SUMB[25][57] ), .CO(
        \mult_22/CARRYB[26][56] ), .S(\mult_22/SUMB[26][56] ) );
  FA_X1 \mult_22/S2_26_55  ( .A(\mult_22/ab[26][55] ), .B(
        \mult_22/CARRYB[25][55] ), .CI(\mult_22/SUMB[25][56] ), .CO(
        \mult_22/CARRYB[26][55] ), .S(\mult_22/SUMB[26][55] ) );
  FA_X1 \mult_22/S2_26_54  ( .A(\mult_22/ab[26][54] ), .B(
        \mult_22/CARRYB[25][54] ), .CI(\mult_22/SUMB[25][55] ), .CO(
        \mult_22/CARRYB[26][54] ), .S(\mult_22/SUMB[26][54] ) );
  FA_X1 \mult_22/S2_26_53  ( .A(\mult_22/ab[26][53] ), .B(
        \mult_22/CARRYB[25][53] ), .CI(\mult_22/SUMB[25][54] ), .CO(
        \mult_22/CARRYB[26][53] ), .S(\mult_22/SUMB[26][53] ) );
  FA_X1 \mult_22/S2_26_52  ( .A(\mult_22/ab[26][52] ), .B(
        \mult_22/CARRYB[25][52] ), .CI(\mult_22/SUMB[25][53] ), .CO(
        \mult_22/CARRYB[26][52] ), .S(\mult_22/SUMB[26][52] ) );
  FA_X1 \mult_22/S2_26_51  ( .A(\mult_22/ab[26][51] ), .B(
        \mult_22/CARRYB[25][51] ), .CI(\mult_22/SUMB[25][52] ), .CO(
        \mult_22/CARRYB[26][51] ), .S(\mult_22/SUMB[26][51] ) );
  FA_X1 \mult_22/S2_26_50  ( .A(\mult_22/ab[26][50] ), .B(
        \mult_22/CARRYB[25][50] ), .CI(\mult_22/SUMB[25][51] ), .CO(
        \mult_22/CARRYB[26][50] ), .S(\mult_22/SUMB[26][50] ) );
  FA_X1 \mult_22/S2_26_49  ( .A(\mult_22/ab[26][49] ), .B(
        \mult_22/CARRYB[25][49] ), .CI(\mult_22/SUMB[25][50] ), .CO(
        \mult_22/CARRYB[26][49] ), .S(\mult_22/SUMB[26][49] ) );
  FA_X1 \mult_22/S2_26_48  ( .A(\mult_22/ab[26][48] ), .B(
        \mult_22/CARRYB[25][48] ), .CI(\mult_22/SUMB[25][49] ), .CO(
        \mult_22/CARRYB[26][48] ), .S(\mult_22/SUMB[26][48] ) );
  FA_X1 \mult_22/S2_26_47  ( .A(\mult_22/ab[26][47] ), .B(
        \mult_22/CARRYB[25][47] ), .CI(\mult_22/SUMB[25][48] ), .CO(
        \mult_22/CARRYB[26][47] ), .S(\mult_22/SUMB[26][47] ) );
  FA_X1 \mult_22/S2_26_46  ( .A(\mult_22/ab[26][46] ), .B(
        \mult_22/CARRYB[25][46] ), .CI(\mult_22/SUMB[25][47] ), .CO(
        \mult_22/CARRYB[26][46] ), .S(\mult_22/SUMB[26][46] ) );
  FA_X1 \mult_22/S2_26_45  ( .A(\mult_22/ab[26][45] ), .B(
        \mult_22/CARRYB[25][45] ), .CI(\mult_22/SUMB[25][46] ), .CO(
        \mult_22/CARRYB[26][45] ), .S(\mult_22/SUMB[26][45] ) );
  FA_X1 \mult_22/S2_26_44  ( .A(\mult_22/ab[26][44] ), .B(
        \mult_22/CARRYB[25][44] ), .CI(\mult_22/SUMB[25][45] ), .CO(
        \mult_22/CARRYB[26][44] ), .S(\mult_22/SUMB[26][44] ) );
  FA_X1 \mult_22/S2_26_43  ( .A(\mult_22/ab[26][43] ), .B(
        \mult_22/CARRYB[25][43] ), .CI(\mult_22/SUMB[25][44] ), .CO(
        \mult_22/CARRYB[26][43] ), .S(\mult_22/SUMB[26][43] ) );
  FA_X1 \mult_22/S2_26_42  ( .A(\mult_22/ab[26][42] ), .B(
        \mult_22/CARRYB[25][42] ), .CI(\mult_22/SUMB[25][43] ), .CO(
        \mult_22/CARRYB[26][42] ), .S(\mult_22/SUMB[26][42] ) );
  FA_X1 \mult_22/S2_26_41  ( .A(\mult_22/ab[26][41] ), .B(
        \mult_22/CARRYB[25][41] ), .CI(\mult_22/SUMB[25][42] ), .CO(
        \mult_22/CARRYB[26][41] ), .S(\mult_22/SUMB[26][41] ) );
  FA_X1 \mult_22/S2_26_38  ( .A(\mult_22/ab[26][38] ), .B(
        \mult_22/CARRYB[25][38] ), .CI(\mult_22/SUMB[25][39] ), .CO(
        \mult_22/CARRYB[26][38] ), .S(\mult_22/SUMB[26][38] ) );
  FA_X1 \mult_22/S2_26_37  ( .A(\mult_22/ab[26][37] ), .B(
        \mult_22/CARRYB[25][37] ), .CI(\mult_22/SUMB[25][38] ), .CO(
        \mult_22/CARRYB[26][37] ), .S(\mult_22/SUMB[26][37] ) );
  FA_X1 \mult_22/S2_26_36  ( .A(\mult_22/ab[26][36] ), .B(
        \mult_22/CARRYB[25][36] ), .CI(\mult_22/SUMB[25][37] ), .CO(
        \mult_22/CARRYB[26][36] ), .S(\mult_22/SUMB[26][36] ) );
  FA_X1 \mult_22/S2_26_33  ( .A(\mult_22/ab[26][33] ), .B(
        \mult_22/CARRYB[25][33] ), .CI(\mult_22/SUMB[25][34] ), .CO(
        \mult_22/CARRYB[26][33] ), .S(\mult_22/SUMB[26][33] ) );
  FA_X1 \mult_22/S2_26_32  ( .A(\mult_22/ab[26][32] ), .B(
        \mult_22/CARRYB[25][32] ), .CI(\mult_22/SUMB[25][33] ), .CO(
        \mult_22/CARRYB[26][32] ), .S(\mult_22/SUMB[26][32] ) );
  FA_X1 \mult_22/S2_26_31  ( .A(\mult_22/ab[26][31] ), .B(
        \mult_22/CARRYB[25][31] ), .CI(\mult_22/SUMB[25][32] ), .CO(
        \mult_22/CARRYB[26][31] ), .S(\mult_22/SUMB[26][31] ) );
  FA_X1 \mult_22/S2_26_30  ( .A(\mult_22/ab[26][30] ), .B(
        \mult_22/CARRYB[25][30] ), .CI(\mult_22/SUMB[25][31] ), .CO(
        \mult_22/CARRYB[26][30] ), .S(\mult_22/SUMB[26][30] ) );
  FA_X1 \mult_22/S2_26_29  ( .A(\mult_22/ab[26][29] ), .B(
        \mult_22/CARRYB[25][29] ), .CI(\mult_22/SUMB[25][30] ), .CO(
        \mult_22/CARRYB[26][29] ), .S(\mult_22/SUMB[26][29] ) );
  FA_X1 \mult_22/S2_26_28  ( .A(\mult_22/ab[26][28] ), .B(
        \mult_22/CARRYB[25][28] ), .CI(\mult_22/SUMB[25][29] ), .CO(
        \mult_22/CARRYB[26][28] ), .S(\mult_22/SUMB[26][28] ) );
  FA_X1 \mult_22/S2_26_27  ( .A(\mult_22/ab[26][27] ), .B(
        \mult_22/CARRYB[25][27] ), .CI(\mult_22/SUMB[25][28] ), .CO(
        \mult_22/CARRYB[26][27] ), .S(\mult_22/SUMB[26][27] ) );
  FA_X1 \mult_22/S2_26_26  ( .A(\mult_22/ab[26][26] ), .B(
        \mult_22/CARRYB[25][26] ), .CI(\mult_22/SUMB[25][27] ), .CO(
        \mult_22/CARRYB[26][26] ), .S(\mult_22/SUMB[26][26] ) );
  FA_X1 \mult_22/S2_26_25  ( .A(\mult_22/ab[26][25] ), .B(
        \mult_22/CARRYB[25][25] ), .CI(\mult_22/SUMB[25][26] ), .CO(
        \mult_22/CARRYB[26][25] ), .S(\mult_22/SUMB[26][25] ) );
  FA_X1 \mult_22/S2_26_24  ( .A(\mult_22/ab[26][24] ), .B(
        \mult_22/CARRYB[25][24] ), .CI(\mult_22/SUMB[25][25] ), .CO(
        \mult_22/CARRYB[26][24] ), .S(\mult_22/SUMB[26][24] ) );
  FA_X1 \mult_22/S2_26_23  ( .A(\mult_22/ab[26][23] ), .B(
        \mult_22/CARRYB[25][23] ), .CI(\mult_22/SUMB[25][24] ), .CO(
        \mult_22/CARRYB[26][23] ), .S(\mult_22/SUMB[26][23] ) );
  FA_X1 \mult_22/S2_26_22  ( .A(\mult_22/ab[26][22] ), .B(
        \mult_22/CARRYB[25][22] ), .CI(\mult_22/SUMB[25][23] ), .CO(
        \mult_22/CARRYB[26][22] ), .S(\mult_22/SUMB[26][22] ) );
  FA_X1 \mult_22/S2_26_21  ( .A(\mult_22/ab[26][21] ), .B(
        \mult_22/CARRYB[25][21] ), .CI(\mult_22/SUMB[25][22] ), .CO(
        \mult_22/CARRYB[26][21] ), .S(\mult_22/SUMB[26][21] ) );
  FA_X1 \mult_22/S2_26_20  ( .A(\mult_22/ab[26][20] ), .B(
        \mult_22/CARRYB[25][20] ), .CI(\mult_22/SUMB[25][21] ), .CO(
        \mult_22/CARRYB[26][20] ), .S(\mult_22/SUMB[26][20] ) );
  FA_X1 \mult_22/S2_26_19  ( .A(\mult_22/ab[26][19] ), .B(
        \mult_22/CARRYB[25][19] ), .CI(\mult_22/SUMB[25][20] ), .CO(
        \mult_22/CARRYB[26][19] ), .S(\mult_22/SUMB[26][19] ) );
  FA_X1 \mult_22/S2_26_18  ( .A(\mult_22/ab[26][18] ), .B(
        \mult_22/CARRYB[25][18] ), .CI(\mult_22/SUMB[25][19] ), .CO(
        \mult_22/CARRYB[26][18] ), .S(\mult_22/SUMB[26][18] ) );
  FA_X1 \mult_22/S2_26_17  ( .A(\mult_22/ab[26][17] ), .B(
        \mult_22/CARRYB[25][17] ), .CI(\mult_22/SUMB[25][18] ), .CO(
        \mult_22/CARRYB[26][17] ), .S(\mult_22/SUMB[26][17] ) );
  FA_X1 \mult_22/S2_26_16  ( .A(\mult_22/ab[26][16] ), .B(
        \mult_22/CARRYB[25][16] ), .CI(\mult_22/SUMB[25][17] ), .CO(
        \mult_22/CARRYB[26][16] ), .S(\mult_22/SUMB[26][16] ) );
  FA_X1 \mult_22/S2_26_15  ( .A(\mult_22/ab[26][15] ), .B(
        \mult_22/CARRYB[25][15] ), .CI(\mult_22/SUMB[25][16] ), .CO(
        \mult_22/CARRYB[26][15] ), .S(\mult_22/SUMB[26][15] ) );
  FA_X1 \mult_22/S2_26_14  ( .A(\mult_22/ab[26][14] ), .B(
        \mult_22/CARRYB[25][14] ), .CI(\mult_22/SUMB[25][15] ), .CO(
        \mult_22/CARRYB[26][14] ), .S(\mult_22/SUMB[26][14] ) );
  FA_X1 \mult_22/S2_26_13  ( .A(\mult_22/ab[26][13] ), .B(
        \mult_22/CARRYB[25][13] ), .CI(\mult_22/SUMB[25][14] ), .CO(
        \mult_22/CARRYB[26][13] ), .S(\mult_22/SUMB[26][13] ) );
  FA_X1 \mult_22/S2_26_12  ( .A(\mult_22/ab[26][12] ), .B(
        \mult_22/CARRYB[25][12] ), .CI(\mult_22/SUMB[25][13] ), .CO(
        \mult_22/CARRYB[26][12] ), .S(\mult_22/SUMB[26][12] ) );
  FA_X1 \mult_22/S2_26_11  ( .A(\mult_22/ab[26][11] ), .B(
        \mult_22/CARRYB[25][11] ), .CI(\mult_22/SUMB[25][12] ), .CO(
        \mult_22/CARRYB[26][11] ), .S(\mult_22/SUMB[26][11] ) );
  FA_X1 \mult_22/S2_26_10  ( .A(\mult_22/ab[26][10] ), .B(
        \mult_22/CARRYB[25][10] ), .CI(\mult_22/SUMB[25][11] ), .CO(
        \mult_22/CARRYB[26][10] ), .S(\mult_22/SUMB[26][10] ) );
  FA_X1 \mult_22/S2_26_9  ( .A(\mult_22/ab[26][9] ), .B(
        \mult_22/CARRYB[25][9] ), .CI(\mult_22/SUMB[25][10] ), .CO(
        \mult_22/CARRYB[26][9] ), .S(\mult_22/SUMB[26][9] ) );
  FA_X1 \mult_22/S2_26_8  ( .A(\mult_22/ab[26][8] ), .B(
        \mult_22/CARRYB[25][8] ), .CI(\mult_22/SUMB[25][9] ), .CO(
        \mult_22/CARRYB[26][8] ), .S(\mult_22/SUMB[26][8] ) );
  FA_X1 \mult_22/S2_26_7  ( .A(\mult_22/ab[26][7] ), .B(
        \mult_22/CARRYB[25][7] ), .CI(\mult_22/SUMB[25][8] ), .CO(
        \mult_22/CARRYB[26][7] ), .S(\mult_22/SUMB[26][7] ) );
  FA_X1 \mult_22/S2_26_6  ( .A(\mult_22/ab[26][6] ), .B(
        \mult_22/CARRYB[25][6] ), .CI(\mult_22/SUMB[25][7] ), .CO(
        \mult_22/CARRYB[26][6] ), .S(\mult_22/SUMB[26][6] ) );
  FA_X1 \mult_22/S2_26_5  ( .A(\mult_22/ab[26][5] ), .B(
        \mult_22/CARRYB[25][5] ), .CI(\mult_22/SUMB[25][6] ), .CO(
        \mult_22/CARRYB[26][5] ), .S(\mult_22/SUMB[26][5] ) );
  FA_X1 \mult_22/S2_26_4  ( .A(\mult_22/ab[26][4] ), .B(
        \mult_22/CARRYB[25][4] ), .CI(\mult_22/SUMB[25][5] ), .CO(
        \mult_22/CARRYB[26][4] ), .S(\mult_22/SUMB[26][4] ) );
  FA_X1 \mult_22/S2_26_3  ( .A(\mult_22/ab[26][3] ), .B(
        \mult_22/CARRYB[25][3] ), .CI(\mult_22/SUMB[25][4] ), .CO(
        \mult_22/CARRYB[26][3] ), .S(\mult_22/SUMB[26][3] ) );
  FA_X1 \mult_22/S2_26_2  ( .A(\mult_22/ab[26][2] ), .B(
        \mult_22/CARRYB[25][2] ), .CI(\mult_22/SUMB[25][3] ), .CO(
        \mult_22/CARRYB[26][2] ), .S(\mult_22/SUMB[26][2] ) );
  FA_X1 \mult_22/S2_26_1  ( .A(\mult_22/ab[26][1] ), .B(
        \mult_22/CARRYB[25][1] ), .CI(\mult_22/SUMB[25][2] ), .CO(
        \mult_22/CARRYB[26][1] ), .S(\mult_22/SUMB[26][1] ) );
  FA_X1 \mult_22/S1_26_0  ( .A(\mult_22/ab[26][0] ), .B(
        \mult_22/CARRYB[25][0] ), .CI(\mult_22/SUMB[25][1] ), .CO(
        \mult_22/CARRYB[26][0] ), .S(N154) );
  FA_X1 \mult_22/S3_27_62  ( .A(\mult_22/ab[27][62] ), .B(
        \mult_22/CARRYB[26][62] ), .CI(\mult_22/ab[26][63] ), .CO(
        \mult_22/CARRYB[27][62] ), .S(\mult_22/SUMB[27][62] ) );
  FA_X1 \mult_22/S2_27_61  ( .A(\mult_22/ab[27][61] ), .B(
        \mult_22/CARRYB[26][61] ), .CI(\mult_22/SUMB[26][62] ), .CO(
        \mult_22/CARRYB[27][61] ), .S(\mult_22/SUMB[27][61] ) );
  FA_X1 \mult_22/S2_27_60  ( .A(\mult_22/ab[27][60] ), .B(
        \mult_22/CARRYB[26][60] ), .CI(\mult_22/SUMB[26][61] ), .CO(
        \mult_22/CARRYB[27][60] ), .S(\mult_22/SUMB[27][60] ) );
  FA_X1 \mult_22/S2_27_59  ( .A(\mult_22/ab[27][59] ), .B(
        \mult_22/CARRYB[26][59] ), .CI(\mult_22/SUMB[26][60] ), .CO(
        \mult_22/CARRYB[27][59] ), .S(\mult_22/SUMB[27][59] ) );
  FA_X1 \mult_22/S2_27_58  ( .A(\mult_22/ab[27][58] ), .B(
        \mult_22/CARRYB[26][58] ), .CI(\mult_22/SUMB[26][59] ), .CO(
        \mult_22/CARRYB[27][58] ), .S(\mult_22/SUMB[27][58] ) );
  FA_X1 \mult_22/S2_27_57  ( .A(\mult_22/ab[27][57] ), .B(
        \mult_22/CARRYB[26][57] ), .CI(\mult_22/SUMB[26][58] ), .CO(
        \mult_22/CARRYB[27][57] ), .S(\mult_22/SUMB[27][57] ) );
  FA_X1 \mult_22/S2_27_56  ( .A(\mult_22/ab[27][56] ), .B(
        \mult_22/CARRYB[26][56] ), .CI(\mult_22/SUMB[26][57] ), .CO(
        \mult_22/CARRYB[27][56] ), .S(\mult_22/SUMB[27][56] ) );
  FA_X1 \mult_22/S2_27_55  ( .A(\mult_22/ab[27][55] ), .B(
        \mult_22/CARRYB[26][55] ), .CI(\mult_22/SUMB[26][56] ), .CO(
        \mult_22/CARRYB[27][55] ), .S(\mult_22/SUMB[27][55] ) );
  FA_X1 \mult_22/S2_27_54  ( .A(\mult_22/ab[27][54] ), .B(
        \mult_22/CARRYB[26][54] ), .CI(\mult_22/SUMB[26][55] ), .CO(
        \mult_22/CARRYB[27][54] ), .S(\mult_22/SUMB[27][54] ) );
  FA_X1 \mult_22/S2_27_53  ( .A(\mult_22/ab[27][53] ), .B(
        \mult_22/CARRYB[26][53] ), .CI(\mult_22/SUMB[26][54] ), .CO(
        \mult_22/CARRYB[27][53] ), .S(\mult_22/SUMB[27][53] ) );
  FA_X1 \mult_22/S2_27_52  ( .A(\mult_22/ab[27][52] ), .B(
        \mult_22/CARRYB[26][52] ), .CI(\mult_22/SUMB[26][53] ), .CO(
        \mult_22/CARRYB[27][52] ), .S(\mult_22/SUMB[27][52] ) );
  FA_X1 \mult_22/S2_27_51  ( .A(\mult_22/ab[27][51] ), .B(
        \mult_22/CARRYB[26][51] ), .CI(\mult_22/SUMB[26][52] ), .CO(
        \mult_22/CARRYB[27][51] ), .S(\mult_22/SUMB[27][51] ) );
  FA_X1 \mult_22/S2_27_50  ( .A(\mult_22/ab[27][50] ), .B(
        \mult_22/CARRYB[26][50] ), .CI(\mult_22/SUMB[26][51] ), .CO(
        \mult_22/CARRYB[27][50] ), .S(\mult_22/SUMB[27][50] ) );
  FA_X1 \mult_22/S2_27_49  ( .A(\mult_22/ab[27][49] ), .B(
        \mult_22/CARRYB[26][49] ), .CI(\mult_22/SUMB[26][50] ), .CO(
        \mult_22/CARRYB[27][49] ), .S(\mult_22/SUMB[27][49] ) );
  FA_X1 \mult_22/S2_27_48  ( .A(\mult_22/ab[27][48] ), .B(
        \mult_22/CARRYB[26][48] ), .CI(\mult_22/SUMB[26][49] ), .CO(
        \mult_22/CARRYB[27][48] ), .S(\mult_22/SUMB[27][48] ) );
  FA_X1 \mult_22/S2_27_47  ( .A(\mult_22/ab[27][47] ), .B(
        \mult_22/CARRYB[26][47] ), .CI(\mult_22/SUMB[26][48] ), .CO(
        \mult_22/CARRYB[27][47] ), .S(\mult_22/SUMB[27][47] ) );
  FA_X1 \mult_22/S2_27_46  ( .A(\mult_22/ab[27][46] ), .B(
        \mult_22/CARRYB[26][46] ), .CI(\mult_22/SUMB[26][47] ), .CO(
        \mult_22/CARRYB[27][46] ), .S(\mult_22/SUMB[27][46] ) );
  FA_X1 \mult_22/S2_27_45  ( .A(\mult_22/ab[27][45] ), .B(
        \mult_22/CARRYB[26][45] ), .CI(\mult_22/SUMB[26][46] ), .CO(
        \mult_22/CARRYB[27][45] ), .S(\mult_22/SUMB[27][45] ) );
  FA_X1 \mult_22/S2_27_44  ( .A(\mult_22/ab[27][44] ), .B(
        \mult_22/CARRYB[26][44] ), .CI(\mult_22/SUMB[26][45] ), .CO(
        \mult_22/CARRYB[27][44] ), .S(\mult_22/SUMB[27][44] ) );
  FA_X1 \mult_22/S2_27_43  ( .A(\mult_22/ab[27][43] ), .B(
        \mult_22/CARRYB[26][43] ), .CI(\mult_22/SUMB[26][44] ), .CO(
        \mult_22/CARRYB[27][43] ), .S(\mult_22/SUMB[27][43] ) );
  FA_X1 \mult_22/S2_27_42  ( .A(\mult_22/ab[27][42] ), .B(
        \mult_22/CARRYB[26][42] ), .CI(\mult_22/SUMB[26][43] ), .CO(
        \mult_22/CARRYB[27][42] ), .S(\mult_22/SUMB[27][42] ) );
  FA_X1 \mult_22/S2_27_41  ( .A(\mult_22/ab[27][41] ), .B(
        \mult_22/CARRYB[26][41] ), .CI(\mult_22/SUMB[26][42] ), .CO(
        \mult_22/CARRYB[27][41] ), .S(\mult_22/SUMB[27][41] ) );
  FA_X1 \mult_22/S2_27_40  ( .A(\mult_22/ab[27][40] ), .B(
        \mult_22/CARRYB[26][40] ), .CI(\mult_22/SUMB[26][41] ), .CO(
        \mult_22/CARRYB[27][40] ), .S(\mult_22/SUMB[27][40] ) );
  FA_X1 \mult_22/S2_27_39  ( .A(\mult_22/ab[27][39] ), .B(
        \mult_22/CARRYB[26][39] ), .CI(\mult_22/SUMB[26][40] ), .CO(
        \mult_22/CARRYB[27][39] ), .S(\mult_22/SUMB[27][39] ) );
  FA_X1 \mult_22/S2_27_38  ( .A(\mult_22/CARRYB[26][38] ), .B(
        \mult_22/ab[27][38] ), .CI(\mult_22/SUMB[26][39] ), .CO(
        \mult_22/CARRYB[27][38] ), .S(\mult_22/SUMB[27][38] ) );
  FA_X1 \mult_22/S2_27_37  ( .A(\mult_22/ab[27][37] ), .B(
        \mult_22/CARRYB[26][37] ), .CI(\mult_22/SUMB[26][38] ), .CO(
        \mult_22/CARRYB[27][37] ), .S(\mult_22/SUMB[27][37] ) );
  FA_X1 \mult_22/S2_27_36  ( .A(\mult_22/ab[27][36] ), .B(
        \mult_22/CARRYB[26][36] ), .CI(\mult_22/SUMB[26][37] ), .CO(
        \mult_22/CARRYB[27][36] ), .S(\mult_22/SUMB[27][36] ) );
  FA_X1 \mult_22/S2_27_35  ( .A(\mult_22/ab[27][35] ), .B(
        \mult_22/CARRYB[26][35] ), .CI(\mult_22/SUMB[26][36] ), .CO(
        \mult_22/CARRYB[27][35] ), .S(\mult_22/SUMB[27][35] ) );
  FA_X1 \mult_22/S2_27_34  ( .A(\mult_22/ab[27][34] ), .B(
        \mult_22/SUMB[26][35] ), .CI(\mult_22/CARRYB[26][34] ), .CO(
        \mult_22/CARRYB[27][34] ), .S(\mult_22/SUMB[27][34] ) );
  FA_X1 \mult_22/S2_27_33  ( .A(\mult_22/ab[27][33] ), .B(
        \mult_22/CARRYB[26][33] ), .CI(\mult_22/SUMB[26][34] ), .CO(
        \mult_22/CARRYB[27][33] ), .S(\mult_22/SUMB[27][33] ) );
  FA_X1 \mult_22/S2_27_32  ( .A(\mult_22/ab[27][32] ), .B(
        \mult_22/CARRYB[26][32] ), .CI(\mult_22/SUMB[26][33] ), .CO(
        \mult_22/CARRYB[27][32] ), .S(\mult_22/SUMB[27][32] ) );
  FA_X1 \mult_22/S2_27_31  ( .A(\mult_22/ab[27][31] ), .B(
        \mult_22/CARRYB[26][31] ), .CI(\mult_22/SUMB[26][32] ), .CO(
        \mult_22/CARRYB[27][31] ), .S(\mult_22/SUMB[27][31] ) );
  FA_X1 \mult_22/S2_27_30  ( .A(\mult_22/ab[27][30] ), .B(
        \mult_22/CARRYB[26][30] ), .CI(\mult_22/SUMB[26][31] ), .CO(
        \mult_22/CARRYB[27][30] ), .S(\mult_22/SUMB[27][30] ) );
  FA_X1 \mult_22/S2_27_29  ( .A(\mult_22/ab[27][29] ), .B(
        \mult_22/CARRYB[26][29] ), .CI(\mult_22/SUMB[26][30] ), .CO(
        \mult_22/CARRYB[27][29] ), .S(\mult_22/SUMB[27][29] ) );
  FA_X1 \mult_22/S2_27_28  ( .A(\mult_22/ab[27][28] ), .B(
        \mult_22/CARRYB[26][28] ), .CI(\mult_22/SUMB[26][29] ), .CO(
        \mult_22/CARRYB[27][28] ), .S(\mult_22/SUMB[27][28] ) );
  FA_X1 \mult_22/S2_27_27  ( .A(\mult_22/ab[27][27] ), .B(
        \mult_22/CARRYB[26][27] ), .CI(\mult_22/SUMB[26][28] ), .CO(
        \mult_22/CARRYB[27][27] ), .S(\mult_22/SUMB[27][27] ) );
  FA_X1 \mult_22/S2_27_26  ( .A(\mult_22/ab[27][26] ), .B(
        \mult_22/CARRYB[26][26] ), .CI(\mult_22/SUMB[26][27] ), .CO(
        \mult_22/CARRYB[27][26] ), .S(\mult_22/SUMB[27][26] ) );
  FA_X1 \mult_22/S2_27_25  ( .A(\mult_22/ab[27][25] ), .B(
        \mult_22/CARRYB[26][25] ), .CI(\mult_22/SUMB[26][26] ), .CO(
        \mult_22/CARRYB[27][25] ), .S(\mult_22/SUMB[27][25] ) );
  FA_X1 \mult_22/S2_27_24  ( .A(\mult_22/ab[27][24] ), .B(
        \mult_22/CARRYB[26][24] ), .CI(\mult_22/SUMB[26][25] ), .CO(
        \mult_22/CARRYB[27][24] ), .S(\mult_22/SUMB[27][24] ) );
  FA_X1 \mult_22/S2_27_23  ( .A(\mult_22/ab[27][23] ), .B(
        \mult_22/CARRYB[26][23] ), .CI(\mult_22/SUMB[26][24] ), .CO(
        \mult_22/CARRYB[27][23] ), .S(\mult_22/SUMB[27][23] ) );
  FA_X1 \mult_22/S2_27_22  ( .A(\mult_22/ab[27][22] ), .B(
        \mult_22/CARRYB[26][22] ), .CI(\mult_22/SUMB[26][23] ), .CO(
        \mult_22/CARRYB[27][22] ), .S(\mult_22/SUMB[27][22] ) );
  FA_X1 \mult_22/S2_27_21  ( .A(\mult_22/ab[27][21] ), .B(
        \mult_22/CARRYB[26][21] ), .CI(\mult_22/SUMB[26][22] ), .CO(
        \mult_22/CARRYB[27][21] ), .S(\mult_22/SUMB[27][21] ) );
  FA_X1 \mult_22/S2_27_20  ( .A(\mult_22/ab[27][20] ), .B(
        \mult_22/CARRYB[26][20] ), .CI(\mult_22/SUMB[26][21] ), .CO(
        \mult_22/CARRYB[27][20] ), .S(\mult_22/SUMB[27][20] ) );
  FA_X1 \mult_22/S2_27_19  ( .A(\mult_22/ab[27][19] ), .B(
        \mult_22/CARRYB[26][19] ), .CI(\mult_22/SUMB[26][20] ), .CO(
        \mult_22/CARRYB[27][19] ), .S(\mult_22/SUMB[27][19] ) );
  FA_X1 \mult_22/S2_27_18  ( .A(\mult_22/ab[27][18] ), .B(
        \mult_22/CARRYB[26][18] ), .CI(\mult_22/SUMB[26][19] ), .CO(
        \mult_22/CARRYB[27][18] ), .S(\mult_22/SUMB[27][18] ) );
  FA_X1 \mult_22/S2_27_17  ( .A(\mult_22/ab[27][17] ), .B(
        \mult_22/CARRYB[26][17] ), .CI(\mult_22/SUMB[26][18] ), .CO(
        \mult_22/CARRYB[27][17] ), .S(\mult_22/SUMB[27][17] ) );
  FA_X1 \mult_22/S2_27_16  ( .A(\mult_22/ab[27][16] ), .B(
        \mult_22/CARRYB[26][16] ), .CI(\mult_22/SUMB[26][17] ), .CO(
        \mult_22/CARRYB[27][16] ), .S(\mult_22/SUMB[27][16] ) );
  FA_X1 \mult_22/S2_27_15  ( .A(\mult_22/ab[27][15] ), .B(
        \mult_22/CARRYB[26][15] ), .CI(\mult_22/SUMB[26][16] ), .CO(
        \mult_22/CARRYB[27][15] ), .S(\mult_22/SUMB[27][15] ) );
  FA_X1 \mult_22/S2_27_14  ( .A(\mult_22/ab[27][14] ), .B(
        \mult_22/CARRYB[26][14] ), .CI(\mult_22/SUMB[26][15] ), .CO(
        \mult_22/CARRYB[27][14] ), .S(\mult_22/SUMB[27][14] ) );
  FA_X1 \mult_22/S2_27_13  ( .A(\mult_22/ab[27][13] ), .B(
        \mult_22/CARRYB[26][13] ), .CI(\mult_22/SUMB[26][14] ), .CO(
        \mult_22/CARRYB[27][13] ), .S(\mult_22/SUMB[27][13] ) );
  FA_X1 \mult_22/S2_27_12  ( .A(\mult_22/ab[27][12] ), .B(
        \mult_22/CARRYB[26][12] ), .CI(\mult_22/SUMB[26][13] ), .CO(
        \mult_22/CARRYB[27][12] ), .S(\mult_22/SUMB[27][12] ) );
  FA_X1 \mult_22/S2_27_11  ( .A(\mult_22/ab[27][11] ), .B(
        \mult_22/CARRYB[26][11] ), .CI(\mult_22/SUMB[26][12] ), .CO(
        \mult_22/CARRYB[27][11] ), .S(\mult_22/SUMB[27][11] ) );
  FA_X1 \mult_22/S2_27_10  ( .A(\mult_22/ab[27][10] ), .B(
        \mult_22/CARRYB[26][10] ), .CI(\mult_22/SUMB[26][11] ), .CO(
        \mult_22/CARRYB[27][10] ), .S(\mult_22/SUMB[27][10] ) );
  FA_X1 \mult_22/S2_27_9  ( .A(\mult_22/ab[27][9] ), .B(
        \mult_22/CARRYB[26][9] ), .CI(\mult_22/SUMB[26][10] ), .CO(
        \mult_22/CARRYB[27][9] ), .S(\mult_22/SUMB[27][9] ) );
  FA_X1 \mult_22/S2_27_8  ( .A(\mult_22/ab[27][8] ), .B(
        \mult_22/CARRYB[26][8] ), .CI(\mult_22/SUMB[26][9] ), .CO(
        \mult_22/CARRYB[27][8] ), .S(\mult_22/SUMB[27][8] ) );
  FA_X1 \mult_22/S2_27_7  ( .A(\mult_22/ab[27][7] ), .B(
        \mult_22/CARRYB[26][7] ), .CI(\mult_22/SUMB[26][8] ), .CO(
        \mult_22/CARRYB[27][7] ), .S(\mult_22/SUMB[27][7] ) );
  FA_X1 \mult_22/S2_27_6  ( .A(\mult_22/ab[27][6] ), .B(
        \mult_22/CARRYB[26][6] ), .CI(\mult_22/SUMB[26][7] ), .CO(
        \mult_22/CARRYB[27][6] ), .S(\mult_22/SUMB[27][6] ) );
  FA_X1 \mult_22/S2_27_5  ( .A(\mult_22/ab[27][5] ), .B(
        \mult_22/CARRYB[26][5] ), .CI(\mult_22/SUMB[26][6] ), .CO(
        \mult_22/CARRYB[27][5] ), .S(\mult_22/SUMB[27][5] ) );
  FA_X1 \mult_22/S2_27_4  ( .A(\mult_22/ab[27][4] ), .B(
        \mult_22/CARRYB[26][4] ), .CI(\mult_22/SUMB[26][5] ), .CO(
        \mult_22/CARRYB[27][4] ), .S(\mult_22/SUMB[27][4] ) );
  FA_X1 \mult_22/S2_27_3  ( .A(\mult_22/ab[27][3] ), .B(
        \mult_22/CARRYB[26][3] ), .CI(\mult_22/SUMB[26][4] ), .CO(
        \mult_22/CARRYB[27][3] ), .S(\mult_22/SUMB[27][3] ) );
  FA_X1 \mult_22/S2_27_2  ( .A(\mult_22/ab[27][2] ), .B(
        \mult_22/CARRYB[26][2] ), .CI(\mult_22/SUMB[26][3] ), .CO(
        \mult_22/CARRYB[27][2] ), .S(\mult_22/SUMB[27][2] ) );
  FA_X1 \mult_22/S2_27_1  ( .A(\mult_22/ab[27][1] ), .B(
        \mult_22/CARRYB[26][1] ), .CI(\mult_22/SUMB[26][2] ), .CO(
        \mult_22/CARRYB[27][1] ), .S(\mult_22/SUMB[27][1] ) );
  FA_X1 \mult_22/S1_27_0  ( .A(\mult_22/ab[27][0] ), .B(
        \mult_22/CARRYB[26][0] ), .CI(\mult_22/SUMB[26][1] ), .CO(
        \mult_22/CARRYB[27][0] ), .S(N155) );
  FA_X1 \mult_22/S3_28_62  ( .A(\mult_22/ab[28][62] ), .B(
        \mult_22/CARRYB[27][62] ), .CI(\mult_22/ab[27][63] ), .CO(
        \mult_22/CARRYB[28][62] ), .S(\mult_22/SUMB[28][62] ) );
  FA_X1 \mult_22/S2_28_61  ( .A(\mult_22/ab[28][61] ), .B(
        \mult_22/CARRYB[27][61] ), .CI(\mult_22/SUMB[27][62] ), .CO(
        \mult_22/CARRYB[28][61] ), .S(\mult_22/SUMB[28][61] ) );
  FA_X1 \mult_22/S2_28_60  ( .A(\mult_22/ab[28][60] ), .B(
        \mult_22/CARRYB[27][60] ), .CI(\mult_22/SUMB[27][61] ), .CO(
        \mult_22/CARRYB[28][60] ), .S(\mult_22/SUMB[28][60] ) );
  FA_X1 \mult_22/S2_28_59  ( .A(\mult_22/ab[28][59] ), .B(
        \mult_22/CARRYB[27][59] ), .CI(\mult_22/SUMB[27][60] ), .CO(
        \mult_22/CARRYB[28][59] ), .S(\mult_22/SUMB[28][59] ) );
  FA_X1 \mult_22/S2_28_58  ( .A(\mult_22/ab[28][58] ), .B(
        \mult_22/CARRYB[27][58] ), .CI(\mult_22/SUMB[27][59] ), .CO(
        \mult_22/CARRYB[28][58] ), .S(\mult_22/SUMB[28][58] ) );
  FA_X1 \mult_22/S2_28_57  ( .A(\mult_22/ab[28][57] ), .B(
        \mult_22/CARRYB[27][57] ), .CI(\mult_22/SUMB[27][58] ), .CO(
        \mult_22/CARRYB[28][57] ), .S(\mult_22/SUMB[28][57] ) );
  FA_X1 \mult_22/S2_28_56  ( .A(\mult_22/ab[28][56] ), .B(
        \mult_22/CARRYB[27][56] ), .CI(\mult_22/SUMB[27][57] ), .CO(
        \mult_22/CARRYB[28][56] ), .S(\mult_22/SUMB[28][56] ) );
  FA_X1 \mult_22/S2_28_55  ( .A(\mult_22/ab[28][55] ), .B(
        \mult_22/CARRYB[27][55] ), .CI(\mult_22/SUMB[27][56] ), .CO(
        \mult_22/CARRYB[28][55] ), .S(\mult_22/SUMB[28][55] ) );
  FA_X1 \mult_22/S2_28_54  ( .A(\mult_22/ab[28][54] ), .B(
        \mult_22/CARRYB[27][54] ), .CI(\mult_22/SUMB[27][55] ), .CO(
        \mult_22/CARRYB[28][54] ), .S(\mult_22/SUMB[28][54] ) );
  FA_X1 \mult_22/S2_28_53  ( .A(\mult_22/ab[28][53] ), .B(
        \mult_22/CARRYB[27][53] ), .CI(\mult_22/SUMB[27][54] ), .CO(
        \mult_22/CARRYB[28][53] ), .S(\mult_22/SUMB[28][53] ) );
  FA_X1 \mult_22/S2_28_52  ( .A(\mult_22/ab[28][52] ), .B(
        \mult_22/CARRYB[27][52] ), .CI(\mult_22/SUMB[27][53] ), .CO(
        \mult_22/CARRYB[28][52] ), .S(\mult_22/SUMB[28][52] ) );
  FA_X1 \mult_22/S2_28_51  ( .A(\mult_22/ab[28][51] ), .B(
        \mult_22/CARRYB[27][51] ), .CI(\mult_22/SUMB[27][52] ), .CO(
        \mult_22/CARRYB[28][51] ), .S(\mult_22/SUMB[28][51] ) );
  FA_X1 \mult_22/S2_28_50  ( .A(\mult_22/ab[28][50] ), .B(
        \mult_22/CARRYB[27][50] ), .CI(\mult_22/SUMB[27][51] ), .CO(
        \mult_22/CARRYB[28][50] ), .S(\mult_22/SUMB[28][50] ) );
  FA_X1 \mult_22/S2_28_49  ( .A(\mult_22/ab[28][49] ), .B(
        \mult_22/CARRYB[27][49] ), .CI(\mult_22/SUMB[27][50] ), .CO(
        \mult_22/CARRYB[28][49] ), .S(\mult_22/SUMB[28][49] ) );
  FA_X1 \mult_22/S2_28_48  ( .A(\mult_22/ab[28][48] ), .B(
        \mult_22/CARRYB[27][48] ), .CI(\mult_22/SUMB[27][49] ), .CO(
        \mult_22/CARRYB[28][48] ), .S(\mult_22/SUMB[28][48] ) );
  FA_X1 \mult_22/S2_28_47  ( .A(\mult_22/ab[28][47] ), .B(
        \mult_22/CARRYB[27][47] ), .CI(\mult_22/SUMB[27][48] ), .CO(
        \mult_22/CARRYB[28][47] ), .S(\mult_22/SUMB[28][47] ) );
  FA_X1 \mult_22/S2_28_46  ( .A(\mult_22/ab[28][46] ), .B(
        \mult_22/CARRYB[27][46] ), .CI(\mult_22/SUMB[27][47] ), .CO(
        \mult_22/CARRYB[28][46] ), .S(\mult_22/SUMB[28][46] ) );
  FA_X1 \mult_22/S2_28_45  ( .A(\mult_22/ab[28][45] ), .B(
        \mult_22/CARRYB[27][45] ), .CI(\mult_22/SUMB[27][46] ), .CO(
        \mult_22/CARRYB[28][45] ), .S(\mult_22/SUMB[28][45] ) );
  FA_X1 \mult_22/S2_28_44  ( .A(\mult_22/ab[28][44] ), .B(
        \mult_22/CARRYB[27][44] ), .CI(\mult_22/SUMB[27][45] ), .CO(
        \mult_22/CARRYB[28][44] ), .S(\mult_22/SUMB[28][44] ) );
  FA_X1 \mult_22/S2_28_43  ( .A(\mult_22/ab[28][43] ), .B(
        \mult_22/CARRYB[27][43] ), .CI(\mult_22/SUMB[27][44] ), .CO(
        \mult_22/CARRYB[28][43] ), .S(\mult_22/SUMB[28][43] ) );
  FA_X1 \mult_22/S2_28_42  ( .A(\mult_22/ab[28][42] ), .B(
        \mult_22/CARRYB[27][42] ), .CI(\mult_22/SUMB[27][43] ), .CO(
        \mult_22/CARRYB[28][42] ), .S(\mult_22/SUMB[28][42] ) );
  FA_X1 \mult_22/S2_28_41  ( .A(\mult_22/ab[28][41] ), .B(
        \mult_22/CARRYB[27][41] ), .CI(\mult_22/SUMB[27][42] ), .CO(
        \mult_22/CARRYB[28][41] ), .S(\mult_22/SUMB[28][41] ) );
  FA_X1 \mult_22/S2_28_40  ( .A(\mult_22/ab[28][40] ), .B(
        \mult_22/CARRYB[27][40] ), .CI(\mult_22/SUMB[27][41] ), .CO(
        \mult_22/CARRYB[28][40] ), .S(\mult_22/SUMB[28][40] ) );
  FA_X1 \mult_22/S2_28_39  ( .A(\mult_22/ab[28][39] ), .B(
        \mult_22/CARRYB[27][39] ), .CI(\mult_22/SUMB[27][40] ), .CO(
        \mult_22/CARRYB[28][39] ), .S(\mult_22/SUMB[28][39] ) );
  FA_X1 \mult_22/S2_28_38  ( .A(\mult_22/ab[28][38] ), .B(
        \mult_22/CARRYB[27][38] ), .CI(\mult_22/SUMB[27][39] ), .CO(
        \mult_22/CARRYB[28][38] ), .S(\mult_22/SUMB[28][38] ) );
  FA_X1 \mult_22/S2_28_37  ( .A(\mult_22/ab[28][37] ), .B(
        \mult_22/CARRYB[27][37] ), .CI(\mult_22/SUMB[27][38] ), .CO(
        \mult_22/CARRYB[28][37] ), .S(\mult_22/SUMB[28][37] ) );
  FA_X1 \mult_22/S2_28_36  ( .A(\mult_22/ab[28][36] ), .B(
        \mult_22/CARRYB[27][36] ), .CI(\mult_22/SUMB[27][37] ), .CO(
        \mult_22/CARRYB[28][36] ), .S(\mult_22/SUMB[28][36] ) );
  FA_X1 \mult_22/S2_28_35  ( .A(\mult_22/ab[28][35] ), .B(
        \mult_22/CARRYB[27][35] ), .CI(\mult_22/SUMB[27][36] ), .CO(
        \mult_22/CARRYB[28][35] ), .S(\mult_22/SUMB[28][35] ) );
  FA_X1 \mult_22/S2_28_34  ( .A(\mult_22/ab[28][34] ), .B(
        \mult_22/CARRYB[27][34] ), .CI(\mult_22/SUMB[27][35] ), .CO(
        \mult_22/CARRYB[28][34] ), .S(\mult_22/SUMB[28][34] ) );
  FA_X1 \mult_22/S2_28_33  ( .A(\mult_22/ab[28][33] ), .B(
        \mult_22/CARRYB[27][33] ), .CI(\mult_22/SUMB[27][34] ), .CO(
        \mult_22/CARRYB[28][33] ), .S(\mult_22/SUMB[28][33] ) );
  FA_X1 \mult_22/S2_28_32  ( .A(\mult_22/ab[28][32] ), .B(
        \mult_22/CARRYB[27][32] ), .CI(\mult_22/SUMB[27][33] ), .CO(
        \mult_22/CARRYB[28][32] ), .S(\mult_22/SUMB[28][32] ) );
  FA_X1 \mult_22/S2_28_31  ( .A(\mult_22/ab[28][31] ), .B(
        \mult_22/CARRYB[27][31] ), .CI(\mult_22/SUMB[27][32] ), .CO(
        \mult_22/CARRYB[28][31] ), .S(\mult_22/SUMB[28][31] ) );
  FA_X1 \mult_22/S2_28_29  ( .A(\mult_22/ab[28][29] ), .B(
        \mult_22/CARRYB[27][29] ), .CI(\mult_22/SUMB[27][30] ), .CO(
        \mult_22/CARRYB[28][29] ), .S(\mult_22/SUMB[28][29] ) );
  FA_X1 \mult_22/S2_28_28  ( .A(\mult_22/ab[28][28] ), .B(
        \mult_22/CARRYB[27][28] ), .CI(\mult_22/SUMB[27][29] ), .CO(
        \mult_22/CARRYB[28][28] ), .S(\mult_22/SUMB[28][28] ) );
  FA_X1 \mult_22/S2_28_27  ( .A(\mult_22/ab[28][27] ), .B(
        \mult_22/CARRYB[27][27] ), .CI(\mult_22/SUMB[27][28] ), .CO(
        \mult_22/CARRYB[28][27] ), .S(\mult_22/SUMB[28][27] ) );
  FA_X1 \mult_22/S2_28_26  ( .A(\mult_22/ab[28][26] ), .B(
        \mult_22/CARRYB[27][26] ), .CI(\mult_22/SUMB[27][27] ), .CO(
        \mult_22/CARRYB[28][26] ), .S(\mult_22/SUMB[28][26] ) );
  FA_X1 \mult_22/S2_28_25  ( .A(\mult_22/ab[28][25] ), .B(
        \mult_22/CARRYB[27][25] ), .CI(\mult_22/SUMB[27][26] ), .CO(
        \mult_22/CARRYB[28][25] ), .S(\mult_22/SUMB[28][25] ) );
  FA_X1 \mult_22/S2_28_24  ( .A(\mult_22/ab[28][24] ), .B(
        \mult_22/CARRYB[27][24] ), .CI(\mult_22/SUMB[27][25] ), .CO(
        \mult_22/CARRYB[28][24] ), .S(\mult_22/SUMB[28][24] ) );
  FA_X1 \mult_22/S2_28_23  ( .A(\mult_22/ab[28][23] ), .B(
        \mult_22/CARRYB[27][23] ), .CI(\mult_22/SUMB[27][24] ), .CO(
        \mult_22/CARRYB[28][23] ), .S(\mult_22/SUMB[28][23] ) );
  FA_X1 \mult_22/S2_28_22  ( .A(\mult_22/ab[28][22] ), .B(
        \mult_22/CARRYB[27][22] ), .CI(\mult_22/SUMB[27][23] ), .CO(
        \mult_22/CARRYB[28][22] ), .S(\mult_22/SUMB[28][22] ) );
  FA_X1 \mult_22/S2_28_21  ( .A(\mult_22/ab[28][21] ), .B(
        \mult_22/CARRYB[27][21] ), .CI(\mult_22/SUMB[27][22] ), .CO(
        \mult_22/CARRYB[28][21] ), .S(\mult_22/SUMB[28][21] ) );
  FA_X1 \mult_22/S2_28_20  ( .A(\mult_22/ab[28][20] ), .B(
        \mult_22/CARRYB[27][20] ), .CI(\mult_22/SUMB[27][21] ), .CO(
        \mult_22/CARRYB[28][20] ), .S(\mult_22/SUMB[28][20] ) );
  FA_X1 \mult_22/S2_28_19  ( .A(\mult_22/ab[28][19] ), .B(
        \mult_22/CARRYB[27][19] ), .CI(\mult_22/SUMB[27][20] ), .CO(
        \mult_22/CARRYB[28][19] ), .S(\mult_22/SUMB[28][19] ) );
  FA_X1 \mult_22/S2_28_18  ( .A(\mult_22/ab[28][18] ), .B(
        \mult_22/CARRYB[27][18] ), .CI(\mult_22/SUMB[27][19] ), .CO(
        \mult_22/CARRYB[28][18] ), .S(\mult_22/SUMB[28][18] ) );
  FA_X1 \mult_22/S2_28_17  ( .A(\mult_22/ab[28][17] ), .B(
        \mult_22/CARRYB[27][17] ), .CI(\mult_22/SUMB[27][18] ), .CO(
        \mult_22/CARRYB[28][17] ), .S(\mult_22/SUMB[28][17] ) );
  FA_X1 \mult_22/S2_28_16  ( .A(\mult_22/ab[28][16] ), .B(
        \mult_22/CARRYB[27][16] ), .CI(\mult_22/SUMB[27][17] ), .CO(
        \mult_22/CARRYB[28][16] ), .S(\mult_22/SUMB[28][16] ) );
  FA_X1 \mult_22/S2_28_15  ( .A(\mult_22/ab[28][15] ), .B(
        \mult_22/CARRYB[27][15] ), .CI(\mult_22/SUMB[27][16] ), .CO(
        \mult_22/CARRYB[28][15] ), .S(\mult_22/SUMB[28][15] ) );
  FA_X1 \mult_22/S2_28_14  ( .A(\mult_22/ab[28][14] ), .B(
        \mult_22/CARRYB[27][14] ), .CI(\mult_22/SUMB[27][15] ), .CO(
        \mult_22/CARRYB[28][14] ), .S(\mult_22/SUMB[28][14] ) );
  FA_X1 \mult_22/S2_28_13  ( .A(\mult_22/ab[28][13] ), .B(
        \mult_22/CARRYB[27][13] ), .CI(\mult_22/SUMB[27][14] ), .CO(
        \mult_22/CARRYB[28][13] ), .S(\mult_22/SUMB[28][13] ) );
  FA_X1 \mult_22/S2_28_12  ( .A(\mult_22/ab[28][12] ), .B(
        \mult_22/CARRYB[27][12] ), .CI(\mult_22/SUMB[27][13] ), .CO(
        \mult_22/CARRYB[28][12] ), .S(\mult_22/SUMB[28][12] ) );
  FA_X1 \mult_22/S2_28_11  ( .A(\mult_22/ab[28][11] ), .B(
        \mult_22/CARRYB[27][11] ), .CI(\mult_22/SUMB[27][12] ), .CO(
        \mult_22/CARRYB[28][11] ), .S(\mult_22/SUMB[28][11] ) );
  FA_X1 \mult_22/S2_28_10  ( .A(\mult_22/ab[28][10] ), .B(
        \mult_22/CARRYB[27][10] ), .CI(\mult_22/SUMB[27][11] ), .CO(
        \mult_22/CARRYB[28][10] ), .S(\mult_22/SUMB[28][10] ) );
  FA_X1 \mult_22/S2_28_9  ( .A(\mult_22/ab[28][9] ), .B(
        \mult_22/CARRYB[27][9] ), .CI(\mult_22/SUMB[27][10] ), .CO(
        \mult_22/CARRYB[28][9] ), .S(\mult_22/SUMB[28][9] ) );
  FA_X1 \mult_22/S2_28_8  ( .A(\mult_22/ab[28][8] ), .B(
        \mult_22/CARRYB[27][8] ), .CI(\mult_22/SUMB[27][9] ), .CO(
        \mult_22/CARRYB[28][8] ), .S(\mult_22/SUMB[28][8] ) );
  FA_X1 \mult_22/S2_28_7  ( .A(\mult_22/ab[28][7] ), .B(
        \mult_22/CARRYB[27][7] ), .CI(\mult_22/SUMB[27][8] ), .CO(
        \mult_22/CARRYB[28][7] ), .S(\mult_22/SUMB[28][7] ) );
  FA_X1 \mult_22/S2_28_6  ( .A(\mult_22/ab[28][6] ), .B(
        \mult_22/CARRYB[27][6] ), .CI(\mult_22/SUMB[27][7] ), .CO(
        \mult_22/CARRYB[28][6] ), .S(\mult_22/SUMB[28][6] ) );
  FA_X1 \mult_22/S2_28_5  ( .A(\mult_22/ab[28][5] ), .B(
        \mult_22/CARRYB[27][5] ), .CI(\mult_22/SUMB[27][6] ), .CO(
        \mult_22/CARRYB[28][5] ), .S(\mult_22/SUMB[28][5] ) );
  FA_X1 \mult_22/S2_28_4  ( .A(\mult_22/ab[28][4] ), .B(
        \mult_22/CARRYB[27][4] ), .CI(\mult_22/SUMB[27][5] ), .CO(
        \mult_22/CARRYB[28][4] ), .S(\mult_22/SUMB[28][4] ) );
  FA_X1 \mult_22/S2_28_3  ( .A(\mult_22/ab[28][3] ), .B(
        \mult_22/CARRYB[27][3] ), .CI(\mult_22/SUMB[27][4] ), .CO(
        \mult_22/CARRYB[28][3] ), .S(\mult_22/SUMB[28][3] ) );
  FA_X1 \mult_22/S2_28_2  ( .A(\mult_22/ab[28][2] ), .B(
        \mult_22/CARRYB[27][2] ), .CI(\mult_22/SUMB[27][3] ), .CO(
        \mult_22/CARRYB[28][2] ), .S(\mult_22/SUMB[28][2] ) );
  FA_X1 \mult_22/S2_28_1  ( .A(\mult_22/ab[28][1] ), .B(
        \mult_22/CARRYB[27][1] ), .CI(\mult_22/SUMB[27][2] ), .CO(
        \mult_22/CARRYB[28][1] ), .S(\mult_22/SUMB[28][1] ) );
  FA_X1 \mult_22/S1_28_0  ( .A(\mult_22/ab[28][0] ), .B(
        \mult_22/CARRYB[27][0] ), .CI(\mult_22/SUMB[27][1] ), .CO(
        \mult_22/CARRYB[28][0] ), .S(N156) );
  FA_X1 \mult_22/S3_29_62  ( .A(\mult_22/ab[29][62] ), .B(
        \mult_22/CARRYB[28][62] ), .CI(\mult_22/ab[28][63] ), .CO(
        \mult_22/CARRYB[29][62] ), .S(\mult_22/SUMB[29][62] ) );
  FA_X1 \mult_22/S2_29_61  ( .A(\mult_22/ab[29][61] ), .B(
        \mult_22/CARRYB[28][61] ), .CI(\mult_22/SUMB[28][62] ), .CO(
        \mult_22/CARRYB[29][61] ), .S(\mult_22/SUMB[29][61] ) );
  FA_X1 \mult_22/S2_29_60  ( .A(\mult_22/ab[29][60] ), .B(
        \mult_22/CARRYB[28][60] ), .CI(\mult_22/SUMB[28][61] ), .CO(
        \mult_22/CARRYB[29][60] ), .S(\mult_22/SUMB[29][60] ) );
  FA_X1 \mult_22/S2_29_59  ( .A(\mult_22/ab[29][59] ), .B(
        \mult_22/CARRYB[28][59] ), .CI(\mult_22/SUMB[28][60] ), .CO(
        \mult_22/CARRYB[29][59] ), .S(\mult_22/SUMB[29][59] ) );
  FA_X1 \mult_22/S2_29_58  ( .A(\mult_22/ab[29][58] ), .B(
        \mult_22/CARRYB[28][58] ), .CI(\mult_22/SUMB[28][59] ), .CO(
        \mult_22/CARRYB[29][58] ), .S(\mult_22/SUMB[29][58] ) );
  FA_X1 \mult_22/S2_29_57  ( .A(\mult_22/ab[29][57] ), .B(
        \mult_22/CARRYB[28][57] ), .CI(\mult_22/SUMB[28][58] ), .CO(
        \mult_22/CARRYB[29][57] ), .S(\mult_22/SUMB[29][57] ) );
  FA_X1 \mult_22/S2_29_56  ( .A(\mult_22/ab[29][56] ), .B(
        \mult_22/CARRYB[28][56] ), .CI(\mult_22/SUMB[28][57] ), .CO(
        \mult_22/CARRYB[29][56] ), .S(\mult_22/SUMB[29][56] ) );
  FA_X1 \mult_22/S2_29_55  ( .A(\mult_22/ab[29][55] ), .B(
        \mult_22/CARRYB[28][55] ), .CI(\mult_22/SUMB[28][56] ), .CO(
        \mult_22/CARRYB[29][55] ), .S(\mult_22/SUMB[29][55] ) );
  FA_X1 \mult_22/S2_29_54  ( .A(\mult_22/ab[29][54] ), .B(
        \mult_22/CARRYB[28][54] ), .CI(\mult_22/SUMB[28][55] ), .CO(
        \mult_22/CARRYB[29][54] ), .S(\mult_22/SUMB[29][54] ) );
  FA_X1 \mult_22/S2_29_53  ( .A(\mult_22/ab[29][53] ), .B(
        \mult_22/CARRYB[28][53] ), .CI(\mult_22/SUMB[28][54] ), .CO(
        \mult_22/CARRYB[29][53] ), .S(\mult_22/SUMB[29][53] ) );
  FA_X1 \mult_22/S2_29_52  ( .A(\mult_22/ab[29][52] ), .B(
        \mult_22/CARRYB[28][52] ), .CI(\mult_22/SUMB[28][53] ), .CO(
        \mult_22/CARRYB[29][52] ), .S(\mult_22/SUMB[29][52] ) );
  FA_X1 \mult_22/S2_29_51  ( .A(\mult_22/ab[29][51] ), .B(
        \mult_22/CARRYB[28][51] ), .CI(\mult_22/SUMB[28][52] ), .CO(
        \mult_22/CARRYB[29][51] ), .S(\mult_22/SUMB[29][51] ) );
  FA_X1 \mult_22/S2_29_50  ( .A(\mult_22/ab[29][50] ), .B(
        \mult_22/CARRYB[28][50] ), .CI(\mult_22/SUMB[28][51] ), .CO(
        \mult_22/CARRYB[29][50] ), .S(\mult_22/SUMB[29][50] ) );
  FA_X1 \mult_22/S2_29_49  ( .A(\mult_22/ab[29][49] ), .B(
        \mult_22/CARRYB[28][49] ), .CI(\mult_22/SUMB[28][50] ), .CO(
        \mult_22/CARRYB[29][49] ), .S(\mult_22/SUMB[29][49] ) );
  FA_X1 \mult_22/S2_29_48  ( .A(\mult_22/ab[29][48] ), .B(
        \mult_22/CARRYB[28][48] ), .CI(\mult_22/SUMB[28][49] ), .CO(
        \mult_22/CARRYB[29][48] ), .S(\mult_22/SUMB[29][48] ) );
  FA_X1 \mult_22/S2_29_47  ( .A(\mult_22/ab[29][47] ), .B(
        \mult_22/CARRYB[28][47] ), .CI(\mult_22/SUMB[28][48] ), .CO(
        \mult_22/CARRYB[29][47] ), .S(\mult_22/SUMB[29][47] ) );
  FA_X1 \mult_22/S2_29_46  ( .A(\mult_22/ab[29][46] ), .B(
        \mult_22/CARRYB[28][46] ), .CI(\mult_22/SUMB[28][47] ), .CO(
        \mult_22/CARRYB[29][46] ), .S(\mult_22/SUMB[29][46] ) );
  FA_X1 \mult_22/S2_29_45  ( .A(\mult_22/ab[29][45] ), .B(
        \mult_22/CARRYB[28][45] ), .CI(\mult_22/SUMB[28][46] ), .CO(
        \mult_22/CARRYB[29][45] ), .S(\mult_22/SUMB[29][45] ) );
  FA_X1 \mult_22/S2_29_44  ( .A(\mult_22/ab[29][44] ), .B(
        \mult_22/CARRYB[28][44] ), .CI(\mult_22/SUMB[28][45] ), .CO(
        \mult_22/CARRYB[29][44] ), .S(\mult_22/SUMB[29][44] ) );
  FA_X1 \mult_22/S2_29_43  ( .A(\mult_22/ab[29][43] ), .B(
        \mult_22/CARRYB[28][43] ), .CI(\mult_22/SUMB[28][44] ), .CO(
        \mult_22/CARRYB[29][43] ), .S(\mult_22/SUMB[29][43] ) );
  FA_X1 \mult_22/S2_29_42  ( .A(\mult_22/ab[29][42] ), .B(
        \mult_22/CARRYB[28][42] ), .CI(\mult_22/SUMB[28][43] ), .CO(
        \mult_22/CARRYB[29][42] ), .S(\mult_22/SUMB[29][42] ) );
  FA_X1 \mult_22/S2_29_41  ( .A(\mult_22/ab[29][41] ), .B(
        \mult_22/CARRYB[28][41] ), .CI(\mult_22/SUMB[28][42] ), .CO(
        \mult_22/CARRYB[29][41] ), .S(\mult_22/SUMB[29][41] ) );
  FA_X1 \mult_22/S2_29_40  ( .A(\mult_22/ab[29][40] ), .B(
        \mult_22/CARRYB[28][40] ), .CI(\mult_22/SUMB[28][41] ), .CO(
        \mult_22/CARRYB[29][40] ), .S(\mult_22/SUMB[29][40] ) );
  FA_X1 \mult_22/S2_29_39  ( .A(\mult_22/ab[29][39] ), .B(
        \mult_22/CARRYB[28][39] ), .CI(\mult_22/SUMB[28][40] ), .CO(
        \mult_22/CARRYB[29][39] ), .S(\mult_22/SUMB[29][39] ) );
  FA_X1 \mult_22/S2_29_38  ( .A(\mult_22/ab[29][38] ), .B(
        \mult_22/CARRYB[28][38] ), .CI(\mult_22/SUMB[28][39] ), .CO(
        \mult_22/CARRYB[29][38] ), .S(\mult_22/SUMB[29][38] ) );
  FA_X1 \mult_22/S2_29_37  ( .A(\mult_22/ab[29][37] ), .B(
        \mult_22/CARRYB[28][37] ), .CI(\mult_22/SUMB[28][38] ), .CO(
        \mult_22/CARRYB[29][37] ), .S(\mult_22/SUMB[29][37] ) );
  FA_X1 \mult_22/S2_29_36  ( .A(\mult_22/ab[29][36] ), .B(
        \mult_22/CARRYB[28][36] ), .CI(\mult_22/SUMB[28][37] ), .CO(
        \mult_22/CARRYB[29][36] ), .S(\mult_22/SUMB[29][36] ) );
  FA_X1 \mult_22/S2_29_35  ( .A(\mult_22/ab[29][35] ), .B(
        \mult_22/CARRYB[28][35] ), .CI(\mult_22/SUMB[28][36] ), .CO(
        \mult_22/CARRYB[29][35] ), .S(\mult_22/SUMB[29][35] ) );
  FA_X1 \mult_22/S2_29_34  ( .A(\mult_22/ab[29][34] ), .B(
        \mult_22/CARRYB[28][34] ), .CI(\mult_22/SUMB[28][35] ), .CO(
        \mult_22/CARRYB[29][34] ), .S(\mult_22/SUMB[29][34] ) );
  FA_X1 \mult_22/S2_29_31  ( .A(\mult_22/ab[29][31] ), .B(
        \mult_22/CARRYB[28][31] ), .CI(\mult_22/SUMB[28][32] ), .CO(
        \mult_22/CARRYB[29][31] ), .S(\mult_22/SUMB[29][31] ) );
  FA_X1 \mult_22/S2_29_30  ( .A(\mult_22/ab[29][30] ), .B(
        \mult_22/CARRYB[28][30] ), .CI(\mult_22/SUMB[28][31] ), .CO(
        \mult_22/CARRYB[29][30] ), .S(\mult_22/SUMB[29][30] ) );
  FA_X1 \mult_22/S2_29_29  ( .A(\mult_22/ab[29][29] ), .B(
        \mult_22/CARRYB[28][29] ), .CI(\mult_22/SUMB[28][30] ), .CO(
        \mult_22/CARRYB[29][29] ), .S(\mult_22/SUMB[29][29] ) );
  FA_X1 \mult_22/S2_29_28  ( .A(\mult_22/ab[29][28] ), .B(
        \mult_22/CARRYB[28][28] ), .CI(\mult_22/SUMB[28][29] ), .CO(
        \mult_22/CARRYB[29][28] ), .S(\mult_22/SUMB[29][28] ) );
  FA_X1 \mult_22/S2_29_27  ( .A(\mult_22/ab[29][27] ), .B(
        \mult_22/CARRYB[28][27] ), .CI(\mult_22/SUMB[28][28] ), .CO(
        \mult_22/CARRYB[29][27] ), .S(\mult_22/SUMB[29][27] ) );
  FA_X1 \mult_22/S2_29_26  ( .A(\mult_22/ab[29][26] ), .B(
        \mult_22/CARRYB[28][26] ), .CI(\mult_22/SUMB[28][27] ), .CO(
        \mult_22/CARRYB[29][26] ), .S(\mult_22/SUMB[29][26] ) );
  FA_X1 \mult_22/S2_29_25  ( .A(\mult_22/ab[29][25] ), .B(
        \mult_22/CARRYB[28][25] ), .CI(\mult_22/SUMB[28][26] ), .CO(
        \mult_22/CARRYB[29][25] ), .S(\mult_22/SUMB[29][25] ) );
  FA_X1 \mult_22/S2_29_24  ( .A(\mult_22/ab[29][24] ), .B(
        \mult_22/CARRYB[28][24] ), .CI(\mult_22/SUMB[28][25] ), .CO(
        \mult_22/CARRYB[29][24] ), .S(\mult_22/SUMB[29][24] ) );
  FA_X1 \mult_22/S2_29_23  ( .A(\mult_22/ab[29][23] ), .B(
        \mult_22/CARRYB[28][23] ), .CI(\mult_22/SUMB[28][24] ), .CO(
        \mult_22/CARRYB[29][23] ), .S(\mult_22/SUMB[29][23] ) );
  FA_X1 \mult_22/S2_29_22  ( .A(\mult_22/ab[29][22] ), .B(
        \mult_22/CARRYB[28][22] ), .CI(\mult_22/SUMB[28][23] ), .CO(
        \mult_22/CARRYB[29][22] ), .S(\mult_22/SUMB[29][22] ) );
  FA_X1 \mult_22/S2_29_21  ( .A(\mult_22/ab[29][21] ), .B(
        \mult_22/CARRYB[28][21] ), .CI(\mult_22/SUMB[28][22] ), .CO(
        \mult_22/CARRYB[29][21] ), .S(\mult_22/SUMB[29][21] ) );
  FA_X1 \mult_22/S2_29_20  ( .A(\mult_22/ab[29][20] ), .B(
        \mult_22/CARRYB[28][20] ), .CI(\mult_22/SUMB[28][21] ), .CO(
        \mult_22/CARRYB[29][20] ), .S(\mult_22/SUMB[29][20] ) );
  FA_X1 \mult_22/S2_29_19  ( .A(\mult_22/ab[29][19] ), .B(
        \mult_22/CARRYB[28][19] ), .CI(\mult_22/SUMB[28][20] ), .CO(
        \mult_22/CARRYB[29][19] ), .S(\mult_22/SUMB[29][19] ) );
  FA_X1 \mult_22/S2_29_18  ( .A(\mult_22/ab[29][18] ), .B(
        \mult_22/CARRYB[28][18] ), .CI(\mult_22/SUMB[28][19] ), .CO(
        \mult_22/CARRYB[29][18] ), .S(\mult_22/SUMB[29][18] ) );
  FA_X1 \mult_22/S2_29_17  ( .A(\mult_22/ab[29][17] ), .B(
        \mult_22/CARRYB[28][17] ), .CI(\mult_22/SUMB[28][18] ), .CO(
        \mult_22/CARRYB[29][17] ), .S(\mult_22/SUMB[29][17] ) );
  FA_X1 \mult_22/S2_29_16  ( .A(\mult_22/ab[29][16] ), .B(
        \mult_22/CARRYB[28][16] ), .CI(\mult_22/SUMB[28][17] ), .CO(
        \mult_22/CARRYB[29][16] ), .S(\mult_22/SUMB[29][16] ) );
  FA_X1 \mult_22/S2_29_15  ( .A(\mult_22/ab[29][15] ), .B(
        \mult_22/CARRYB[28][15] ), .CI(\mult_22/SUMB[28][16] ), .CO(
        \mult_22/CARRYB[29][15] ), .S(\mult_22/SUMB[29][15] ) );
  FA_X1 \mult_22/S2_29_14  ( .A(\mult_22/ab[29][14] ), .B(
        \mult_22/CARRYB[28][14] ), .CI(\mult_22/SUMB[28][15] ), .CO(
        \mult_22/CARRYB[29][14] ), .S(\mult_22/SUMB[29][14] ) );
  FA_X1 \mult_22/S2_29_13  ( .A(\mult_22/ab[29][13] ), .B(
        \mult_22/CARRYB[28][13] ), .CI(\mult_22/SUMB[28][14] ), .CO(
        \mult_22/CARRYB[29][13] ), .S(\mult_22/SUMB[29][13] ) );
  FA_X1 \mult_22/S2_29_12  ( .A(\mult_22/ab[29][12] ), .B(
        \mult_22/CARRYB[28][12] ), .CI(\mult_22/SUMB[28][13] ), .CO(
        \mult_22/CARRYB[29][12] ), .S(\mult_22/SUMB[29][12] ) );
  FA_X1 \mult_22/S2_29_11  ( .A(\mult_22/ab[29][11] ), .B(
        \mult_22/CARRYB[28][11] ), .CI(\mult_22/SUMB[28][12] ), .CO(
        \mult_22/CARRYB[29][11] ), .S(\mult_22/SUMB[29][11] ) );
  FA_X1 \mult_22/S2_29_10  ( .A(\mult_22/ab[29][10] ), .B(
        \mult_22/CARRYB[28][10] ), .CI(\mult_22/SUMB[28][11] ), .CO(
        \mult_22/CARRYB[29][10] ), .S(\mult_22/SUMB[29][10] ) );
  FA_X1 \mult_22/S2_29_9  ( .A(\mult_22/ab[29][9] ), .B(
        \mult_22/CARRYB[28][9] ), .CI(\mult_22/SUMB[28][10] ), .CO(
        \mult_22/CARRYB[29][9] ), .S(\mult_22/SUMB[29][9] ) );
  FA_X1 \mult_22/S2_29_8  ( .A(\mult_22/ab[29][8] ), .B(
        \mult_22/CARRYB[28][8] ), .CI(\mult_22/SUMB[28][9] ), .CO(
        \mult_22/CARRYB[29][8] ), .S(\mult_22/SUMB[29][8] ) );
  FA_X1 \mult_22/S2_29_7  ( .A(\mult_22/ab[29][7] ), .B(
        \mult_22/CARRYB[28][7] ), .CI(\mult_22/SUMB[28][8] ), .CO(
        \mult_22/CARRYB[29][7] ), .S(\mult_22/SUMB[29][7] ) );
  FA_X1 \mult_22/S2_29_6  ( .A(\mult_22/ab[29][6] ), .B(
        \mult_22/CARRYB[28][6] ), .CI(\mult_22/SUMB[28][7] ), .CO(
        \mult_22/CARRYB[29][6] ), .S(\mult_22/SUMB[29][6] ) );
  FA_X1 \mult_22/S2_29_5  ( .A(\mult_22/ab[29][5] ), .B(
        \mult_22/CARRYB[28][5] ), .CI(\mult_22/SUMB[28][6] ), .CO(
        \mult_22/CARRYB[29][5] ), .S(\mult_22/SUMB[29][5] ) );
  FA_X1 \mult_22/S2_29_4  ( .A(\mult_22/ab[29][4] ), .B(
        \mult_22/CARRYB[28][4] ), .CI(\mult_22/SUMB[28][5] ), .CO(
        \mult_22/CARRYB[29][4] ), .S(\mult_22/SUMB[29][4] ) );
  FA_X1 \mult_22/S2_29_3  ( .A(\mult_22/ab[29][3] ), .B(
        \mult_22/CARRYB[28][3] ), .CI(\mult_22/SUMB[28][4] ), .CO(
        \mult_22/CARRYB[29][3] ), .S(\mult_22/SUMB[29][3] ) );
  FA_X1 \mult_22/S2_29_2  ( .A(\mult_22/ab[29][2] ), .B(
        \mult_22/CARRYB[28][2] ), .CI(\mult_22/SUMB[28][3] ), .CO(
        \mult_22/CARRYB[29][2] ), .S(\mult_22/SUMB[29][2] ) );
  FA_X1 \mult_22/S2_29_1  ( .A(\mult_22/ab[29][1] ), .B(
        \mult_22/CARRYB[28][1] ), .CI(\mult_22/SUMB[28][2] ), .CO(
        \mult_22/CARRYB[29][1] ), .S(\mult_22/SUMB[29][1] ) );
  FA_X1 \mult_22/S1_29_0  ( .A(\mult_22/ab[29][0] ), .B(
        \mult_22/CARRYB[28][0] ), .CI(\mult_22/SUMB[28][1] ), .CO(
        \mult_22/CARRYB[29][0] ), .S(N157) );
  FA_X1 \mult_22/S3_30_62  ( .A(\mult_22/ab[30][62] ), .B(
        \mult_22/CARRYB[29][62] ), .CI(\mult_22/ab[29][63] ), .CO(
        \mult_22/CARRYB[30][62] ), .S(\mult_22/SUMB[30][62] ) );
  FA_X1 \mult_22/S2_30_61  ( .A(\mult_22/ab[30][61] ), .B(
        \mult_22/CARRYB[29][61] ), .CI(\mult_22/SUMB[29][62] ), .CO(
        \mult_22/CARRYB[30][61] ), .S(\mult_22/SUMB[30][61] ) );
  FA_X1 \mult_22/S2_30_60  ( .A(\mult_22/ab[30][60] ), .B(
        \mult_22/CARRYB[29][60] ), .CI(\mult_22/SUMB[29][61] ), .CO(
        \mult_22/CARRYB[30][60] ), .S(\mult_22/SUMB[30][60] ) );
  FA_X1 \mult_22/S2_30_59  ( .A(\mult_22/ab[30][59] ), .B(
        \mult_22/CARRYB[29][59] ), .CI(\mult_22/SUMB[29][60] ), .CO(
        \mult_22/CARRYB[30][59] ), .S(\mult_22/SUMB[30][59] ) );
  FA_X1 \mult_22/S2_30_58  ( .A(\mult_22/ab[30][58] ), .B(
        \mult_22/CARRYB[29][58] ), .CI(\mult_22/SUMB[29][59] ), .CO(
        \mult_22/CARRYB[30][58] ), .S(\mult_22/SUMB[30][58] ) );
  FA_X1 \mult_22/S2_30_57  ( .A(\mult_22/ab[30][57] ), .B(
        \mult_22/CARRYB[29][57] ), .CI(\mult_22/SUMB[29][58] ), .CO(
        \mult_22/CARRYB[30][57] ), .S(\mult_22/SUMB[30][57] ) );
  FA_X1 \mult_22/S2_30_56  ( .A(\mult_22/ab[30][56] ), .B(
        \mult_22/CARRYB[29][56] ), .CI(\mult_22/SUMB[29][57] ), .CO(
        \mult_22/CARRYB[30][56] ), .S(\mult_22/SUMB[30][56] ) );
  FA_X1 \mult_22/S2_30_55  ( .A(\mult_22/ab[30][55] ), .B(
        \mult_22/CARRYB[29][55] ), .CI(\mult_22/SUMB[29][56] ), .CO(
        \mult_22/CARRYB[30][55] ), .S(\mult_22/SUMB[30][55] ) );
  FA_X1 \mult_22/S2_30_54  ( .A(\mult_22/ab[30][54] ), .B(
        \mult_22/CARRYB[29][54] ), .CI(\mult_22/SUMB[29][55] ), .CO(
        \mult_22/CARRYB[30][54] ), .S(\mult_22/SUMB[30][54] ) );
  FA_X1 \mult_22/S2_30_53  ( .A(\mult_22/ab[30][53] ), .B(
        \mult_22/CARRYB[29][53] ), .CI(\mult_22/SUMB[29][54] ), .CO(
        \mult_22/CARRYB[30][53] ), .S(\mult_22/SUMB[30][53] ) );
  FA_X1 \mult_22/S2_30_52  ( .A(\mult_22/ab[30][52] ), .B(
        \mult_22/CARRYB[29][52] ), .CI(\mult_22/SUMB[29][53] ), .CO(
        \mult_22/CARRYB[30][52] ), .S(\mult_22/SUMB[30][52] ) );
  FA_X1 \mult_22/S2_30_51  ( .A(\mult_22/ab[30][51] ), .B(
        \mult_22/CARRYB[29][51] ), .CI(\mult_22/SUMB[29][52] ), .CO(
        \mult_22/CARRYB[30][51] ), .S(\mult_22/SUMB[30][51] ) );
  FA_X1 \mult_22/S2_30_50  ( .A(\mult_22/ab[30][50] ), .B(
        \mult_22/CARRYB[29][50] ), .CI(\mult_22/SUMB[29][51] ), .CO(
        \mult_22/CARRYB[30][50] ), .S(\mult_22/SUMB[30][50] ) );
  FA_X1 \mult_22/S2_30_49  ( .A(\mult_22/ab[30][49] ), .B(
        \mult_22/CARRYB[29][49] ), .CI(\mult_22/SUMB[29][50] ), .CO(
        \mult_22/CARRYB[30][49] ), .S(\mult_22/SUMB[30][49] ) );
  FA_X1 \mult_22/S2_30_48  ( .A(\mult_22/ab[30][48] ), .B(
        \mult_22/CARRYB[29][48] ), .CI(\mult_22/SUMB[29][49] ), .CO(
        \mult_22/CARRYB[30][48] ), .S(\mult_22/SUMB[30][48] ) );
  FA_X1 \mult_22/S2_30_47  ( .A(\mult_22/ab[30][47] ), .B(
        \mult_22/CARRYB[29][47] ), .CI(\mult_22/SUMB[29][48] ), .CO(
        \mult_22/CARRYB[30][47] ), .S(\mult_22/SUMB[30][47] ) );
  FA_X1 \mult_22/S2_30_46  ( .A(\mult_22/ab[30][46] ), .B(
        \mult_22/CARRYB[29][46] ), .CI(\mult_22/SUMB[29][47] ), .CO(
        \mult_22/CARRYB[30][46] ), .S(\mult_22/SUMB[30][46] ) );
  FA_X1 \mult_22/S2_30_45  ( .A(\mult_22/ab[30][45] ), .B(
        \mult_22/CARRYB[29][45] ), .CI(\mult_22/SUMB[29][46] ), .CO(
        \mult_22/CARRYB[30][45] ), .S(\mult_22/SUMB[30][45] ) );
  FA_X1 \mult_22/S2_30_44  ( .A(\mult_22/ab[30][44] ), .B(
        \mult_22/CARRYB[29][44] ), .CI(\mult_22/SUMB[29][45] ), .CO(
        \mult_22/CARRYB[30][44] ), .S(\mult_22/SUMB[30][44] ) );
  FA_X1 \mult_22/S2_30_43  ( .A(\mult_22/ab[30][43] ), .B(
        \mult_22/CARRYB[29][43] ), .CI(\mult_22/SUMB[29][44] ), .CO(
        \mult_22/CARRYB[30][43] ), .S(\mult_22/SUMB[30][43] ) );
  FA_X1 \mult_22/S2_30_42  ( .A(\mult_22/ab[30][42] ), .B(
        \mult_22/CARRYB[29][42] ), .CI(\mult_22/SUMB[29][43] ), .CO(
        \mult_22/CARRYB[30][42] ), .S(\mult_22/SUMB[30][42] ) );
  FA_X1 \mult_22/S2_30_41  ( .A(\mult_22/ab[30][41] ), .B(
        \mult_22/CARRYB[29][41] ), .CI(\mult_22/SUMB[29][42] ), .CO(
        \mult_22/CARRYB[30][41] ), .S(\mult_22/SUMB[30][41] ) );
  FA_X1 \mult_22/S2_30_40  ( .A(\mult_22/ab[30][40] ), .B(
        \mult_22/CARRYB[29][40] ), .CI(\mult_22/SUMB[29][41] ), .CO(
        \mult_22/CARRYB[30][40] ), .S(\mult_22/SUMB[30][40] ) );
  FA_X1 \mult_22/S2_30_39  ( .A(\mult_22/ab[30][39] ), .B(
        \mult_22/CARRYB[29][39] ), .CI(\mult_22/SUMB[29][40] ), .CO(
        \mult_22/CARRYB[30][39] ), .S(\mult_22/SUMB[30][39] ) );
  FA_X1 \mult_22/S2_30_38  ( .A(\mult_22/ab[30][38] ), .B(
        \mult_22/CARRYB[29][38] ), .CI(\mult_22/SUMB[29][39] ), .CO(
        \mult_22/CARRYB[30][38] ), .S(\mult_22/SUMB[30][38] ) );
  FA_X1 \mult_22/S2_30_37  ( .A(\mult_22/ab[30][37] ), .B(
        \mult_22/CARRYB[29][37] ), .CI(\mult_22/SUMB[29][38] ), .CO(
        \mult_22/CARRYB[30][37] ), .S(\mult_22/SUMB[30][37] ) );
  FA_X1 \mult_22/S2_30_36  ( .A(\mult_22/CARRYB[29][36] ), .B(
        \mult_22/ab[30][36] ), .CI(\mult_22/SUMB[29][37] ), .CO(
        \mult_22/CARRYB[30][36] ), .S(\mult_22/SUMB[30][36] ) );
  FA_X1 \mult_22/S2_30_35  ( .A(\mult_22/ab[30][35] ), .B(
        \mult_22/CARRYB[29][35] ), .CI(\mult_22/SUMB[29][36] ), .CO(
        \mult_22/CARRYB[30][35] ), .S(\mult_22/SUMB[30][35] ) );
  FA_X1 \mult_22/S2_30_34  ( .A(\mult_22/ab[30][34] ), .B(
        \mult_22/CARRYB[29][34] ), .CI(\mult_22/SUMB[29][35] ), .CO(
        \mult_22/CARRYB[30][34] ), .S(\mult_22/SUMB[30][34] ) );
  FA_X1 \mult_22/S2_30_33  ( .A(\mult_22/ab[30][33] ), .B(
        \mult_22/CARRYB[29][33] ), .CI(\mult_22/SUMB[29][34] ), .CO(
        \mult_22/CARRYB[30][33] ), .S(\mult_22/SUMB[30][33] ) );
  FA_X1 \mult_22/S2_30_31  ( .A(\mult_22/ab[30][31] ), .B(
        \mult_22/CARRYB[29][31] ), .CI(\mult_22/SUMB[29][32] ), .CO(
        \mult_22/CARRYB[30][31] ), .S(\mult_22/SUMB[30][31] ) );
  FA_X1 \mult_22/S2_30_30  ( .A(\mult_22/ab[30][30] ), .B(
        \mult_22/CARRYB[29][30] ), .CI(\mult_22/SUMB[29][31] ), .CO(
        \mult_22/CARRYB[30][30] ), .S(\mult_22/SUMB[30][30] ) );
  FA_X1 \mult_22/S2_30_29  ( .A(\mult_22/ab[30][29] ), .B(
        \mult_22/CARRYB[29][29] ), .CI(\mult_22/SUMB[29][30] ), .CO(
        \mult_22/CARRYB[30][29] ), .S(\mult_22/SUMB[30][29] ) );
  FA_X1 \mult_22/S2_30_28  ( .A(\mult_22/ab[30][28] ), .B(
        \mult_22/CARRYB[29][28] ), .CI(\mult_22/SUMB[29][29] ), .CO(
        \mult_22/CARRYB[30][28] ), .S(\mult_22/SUMB[30][28] ) );
  FA_X1 \mult_22/S2_30_27  ( .A(\mult_22/ab[30][27] ), .B(
        \mult_22/CARRYB[29][27] ), .CI(\mult_22/SUMB[29][28] ), .CO(
        \mult_22/CARRYB[30][27] ), .S(\mult_22/SUMB[30][27] ) );
  FA_X1 \mult_22/S2_30_26  ( .A(\mult_22/ab[30][26] ), .B(
        \mult_22/CARRYB[29][26] ), .CI(\mult_22/SUMB[29][27] ), .CO(
        \mult_22/CARRYB[30][26] ), .S(\mult_22/SUMB[30][26] ) );
  FA_X1 \mult_22/S2_30_25  ( .A(\mult_22/ab[30][25] ), .B(
        \mult_22/CARRYB[29][25] ), .CI(\mult_22/SUMB[29][26] ), .CO(
        \mult_22/CARRYB[30][25] ), .S(\mult_22/SUMB[30][25] ) );
  FA_X1 \mult_22/S2_30_24  ( .A(\mult_22/ab[30][24] ), .B(
        \mult_22/CARRYB[29][24] ), .CI(\mult_22/SUMB[29][25] ), .CO(
        \mult_22/CARRYB[30][24] ), .S(\mult_22/SUMB[30][24] ) );
  FA_X1 \mult_22/S2_30_23  ( .A(\mult_22/ab[30][23] ), .B(
        \mult_22/CARRYB[29][23] ), .CI(\mult_22/SUMB[29][24] ), .CO(
        \mult_22/CARRYB[30][23] ), .S(\mult_22/SUMB[30][23] ) );
  FA_X1 \mult_22/S2_30_22  ( .A(\mult_22/ab[30][22] ), .B(
        \mult_22/CARRYB[29][22] ), .CI(\mult_22/SUMB[29][23] ), .CO(
        \mult_22/CARRYB[30][22] ), .S(\mult_22/SUMB[30][22] ) );
  FA_X1 \mult_22/S2_30_21  ( .A(\mult_22/ab[30][21] ), .B(
        \mult_22/CARRYB[29][21] ), .CI(\mult_22/SUMB[29][22] ), .CO(
        \mult_22/CARRYB[30][21] ), .S(\mult_22/SUMB[30][21] ) );
  FA_X1 \mult_22/S2_30_20  ( .A(\mult_22/ab[30][20] ), .B(
        \mult_22/CARRYB[29][20] ), .CI(\mult_22/SUMB[29][21] ), .CO(
        \mult_22/CARRYB[30][20] ), .S(\mult_22/SUMB[30][20] ) );
  FA_X1 \mult_22/S2_30_19  ( .A(\mult_22/ab[30][19] ), .B(
        \mult_22/CARRYB[29][19] ), .CI(\mult_22/SUMB[29][20] ), .CO(
        \mult_22/CARRYB[30][19] ), .S(\mult_22/SUMB[30][19] ) );
  FA_X1 \mult_22/S2_30_18  ( .A(\mult_22/ab[30][18] ), .B(
        \mult_22/CARRYB[29][18] ), .CI(\mult_22/SUMB[29][19] ), .CO(
        \mult_22/CARRYB[30][18] ), .S(\mult_22/SUMB[30][18] ) );
  FA_X1 \mult_22/S2_30_17  ( .A(\mult_22/ab[30][17] ), .B(
        \mult_22/CARRYB[29][17] ), .CI(\mult_22/SUMB[29][18] ), .CO(
        \mult_22/CARRYB[30][17] ), .S(\mult_22/SUMB[30][17] ) );
  FA_X1 \mult_22/S2_30_16  ( .A(\mult_22/ab[30][16] ), .B(
        \mult_22/CARRYB[29][16] ), .CI(\mult_22/SUMB[29][17] ), .CO(
        \mult_22/CARRYB[30][16] ), .S(\mult_22/SUMB[30][16] ) );
  FA_X1 \mult_22/S2_30_15  ( .A(\mult_22/ab[30][15] ), .B(
        \mult_22/CARRYB[29][15] ), .CI(\mult_22/SUMB[29][16] ), .CO(
        \mult_22/CARRYB[30][15] ), .S(\mult_22/SUMB[30][15] ) );
  FA_X1 \mult_22/S2_30_14  ( .A(\mult_22/ab[30][14] ), .B(
        \mult_22/CARRYB[29][14] ), .CI(\mult_22/SUMB[29][15] ), .CO(
        \mult_22/CARRYB[30][14] ), .S(\mult_22/SUMB[30][14] ) );
  FA_X1 \mult_22/S2_30_13  ( .A(\mult_22/ab[30][13] ), .B(
        \mult_22/CARRYB[29][13] ), .CI(\mult_22/SUMB[29][14] ), .CO(
        \mult_22/CARRYB[30][13] ), .S(\mult_22/SUMB[30][13] ) );
  FA_X1 \mult_22/S2_30_12  ( .A(\mult_22/ab[30][12] ), .B(
        \mult_22/CARRYB[29][12] ), .CI(\mult_22/SUMB[29][13] ), .CO(
        \mult_22/CARRYB[30][12] ), .S(\mult_22/SUMB[30][12] ) );
  FA_X1 \mult_22/S2_30_11  ( .A(\mult_22/ab[30][11] ), .B(
        \mult_22/CARRYB[29][11] ), .CI(\mult_22/SUMB[29][12] ), .CO(
        \mult_22/CARRYB[30][11] ), .S(\mult_22/SUMB[30][11] ) );
  FA_X1 \mult_22/S2_30_10  ( .A(\mult_22/ab[30][10] ), .B(
        \mult_22/CARRYB[29][10] ), .CI(\mult_22/SUMB[29][11] ), .CO(
        \mult_22/CARRYB[30][10] ), .S(\mult_22/SUMB[30][10] ) );
  FA_X1 \mult_22/S2_30_9  ( .A(\mult_22/ab[30][9] ), .B(
        \mult_22/CARRYB[29][9] ), .CI(\mult_22/SUMB[29][10] ), .CO(
        \mult_22/CARRYB[30][9] ), .S(\mult_22/SUMB[30][9] ) );
  FA_X1 \mult_22/S2_30_8  ( .A(\mult_22/ab[30][8] ), .B(
        \mult_22/CARRYB[29][8] ), .CI(\mult_22/SUMB[29][9] ), .CO(
        \mult_22/CARRYB[30][8] ), .S(\mult_22/SUMB[30][8] ) );
  FA_X1 \mult_22/S2_30_7  ( .A(\mult_22/ab[30][7] ), .B(
        \mult_22/CARRYB[29][7] ), .CI(\mult_22/SUMB[29][8] ), .CO(
        \mult_22/CARRYB[30][7] ), .S(\mult_22/SUMB[30][7] ) );
  FA_X1 \mult_22/S2_30_6  ( .A(\mult_22/ab[30][6] ), .B(
        \mult_22/CARRYB[29][6] ), .CI(\mult_22/SUMB[29][7] ), .CO(
        \mult_22/CARRYB[30][6] ), .S(\mult_22/SUMB[30][6] ) );
  FA_X1 \mult_22/S2_30_5  ( .A(\mult_22/ab[30][5] ), .B(
        \mult_22/CARRYB[29][5] ), .CI(\mult_22/SUMB[29][6] ), .CO(
        \mult_22/CARRYB[30][5] ), .S(\mult_22/SUMB[30][5] ) );
  FA_X1 \mult_22/S2_30_4  ( .A(\mult_22/ab[30][4] ), .B(
        \mult_22/CARRYB[29][4] ), .CI(\mult_22/SUMB[29][5] ), .CO(
        \mult_22/CARRYB[30][4] ), .S(\mult_22/SUMB[30][4] ) );
  FA_X1 \mult_22/S2_30_3  ( .A(\mult_22/ab[30][3] ), .B(
        \mult_22/CARRYB[29][3] ), .CI(\mult_22/SUMB[29][4] ), .CO(
        \mult_22/CARRYB[30][3] ), .S(\mult_22/SUMB[30][3] ) );
  FA_X1 \mult_22/S2_30_2  ( .A(\mult_22/ab[30][2] ), .B(
        \mult_22/CARRYB[29][2] ), .CI(\mult_22/SUMB[29][3] ), .CO(
        \mult_22/CARRYB[30][2] ), .S(\mult_22/SUMB[30][2] ) );
  FA_X1 \mult_22/S2_30_1  ( .A(\mult_22/ab[30][1] ), .B(
        \mult_22/CARRYB[29][1] ), .CI(\mult_22/SUMB[29][2] ), .CO(
        \mult_22/CARRYB[30][1] ), .S(\mult_22/SUMB[30][1] ) );
  FA_X1 \mult_22/S1_30_0  ( .A(\mult_22/ab[30][0] ), .B(
        \mult_22/CARRYB[29][0] ), .CI(\mult_22/SUMB[29][1] ), .CO(
        \mult_22/CARRYB[30][0] ), .S(N158) );
  FA_X1 \mult_22/S3_31_62  ( .A(\mult_22/ab[31][62] ), .B(
        \mult_22/CARRYB[30][62] ), .CI(\mult_22/ab[30][63] ), .CO(
        \mult_22/CARRYB[31][62] ), .S(\mult_22/SUMB[31][62] ) );
  FA_X1 \mult_22/S2_31_61  ( .A(\mult_22/ab[31][61] ), .B(
        \mult_22/CARRYB[30][61] ), .CI(\mult_22/SUMB[30][62] ), .CO(
        \mult_22/CARRYB[31][61] ), .S(\mult_22/SUMB[31][61] ) );
  FA_X1 \mult_22/S2_31_60  ( .A(\mult_22/ab[31][60] ), .B(
        \mult_22/CARRYB[30][60] ), .CI(\mult_22/SUMB[30][61] ), .CO(
        \mult_22/CARRYB[31][60] ), .S(\mult_22/SUMB[31][60] ) );
  FA_X1 \mult_22/S2_31_59  ( .A(\mult_22/ab[31][59] ), .B(
        \mult_22/CARRYB[30][59] ), .CI(\mult_22/SUMB[30][60] ), .CO(
        \mult_22/CARRYB[31][59] ), .S(\mult_22/SUMB[31][59] ) );
  FA_X1 \mult_22/S2_31_58  ( .A(\mult_22/ab[31][58] ), .B(
        \mult_22/CARRYB[30][58] ), .CI(\mult_22/SUMB[30][59] ), .CO(
        \mult_22/CARRYB[31][58] ), .S(\mult_22/SUMB[31][58] ) );
  FA_X1 \mult_22/S2_31_57  ( .A(\mult_22/ab[31][57] ), .B(
        \mult_22/CARRYB[30][57] ), .CI(\mult_22/SUMB[30][58] ), .CO(
        \mult_22/CARRYB[31][57] ), .S(\mult_22/SUMB[31][57] ) );
  FA_X1 \mult_22/S2_31_56  ( .A(\mult_22/ab[31][56] ), .B(
        \mult_22/CARRYB[30][56] ), .CI(\mult_22/SUMB[30][57] ), .CO(
        \mult_22/CARRYB[31][56] ), .S(\mult_22/SUMB[31][56] ) );
  FA_X1 \mult_22/S2_31_55  ( .A(\mult_22/ab[31][55] ), .B(
        \mult_22/CARRYB[30][55] ), .CI(\mult_22/SUMB[30][56] ), .CO(
        \mult_22/CARRYB[31][55] ), .S(\mult_22/SUMB[31][55] ) );
  FA_X1 \mult_22/S2_31_54  ( .A(\mult_22/ab[31][54] ), .B(
        \mult_22/CARRYB[30][54] ), .CI(\mult_22/SUMB[30][55] ), .CO(
        \mult_22/CARRYB[31][54] ), .S(\mult_22/SUMB[31][54] ) );
  FA_X1 \mult_22/S2_31_53  ( .A(\mult_22/ab[31][53] ), .B(
        \mult_22/CARRYB[30][53] ), .CI(\mult_22/SUMB[30][54] ), .CO(
        \mult_22/CARRYB[31][53] ), .S(\mult_22/SUMB[31][53] ) );
  FA_X1 \mult_22/S2_31_52  ( .A(\mult_22/ab[31][52] ), .B(
        \mult_22/CARRYB[30][52] ), .CI(\mult_22/SUMB[30][53] ), .CO(
        \mult_22/CARRYB[31][52] ), .S(\mult_22/SUMB[31][52] ) );
  FA_X1 \mult_22/S2_31_51  ( .A(\mult_22/ab[31][51] ), .B(
        \mult_22/CARRYB[30][51] ), .CI(\mult_22/SUMB[30][52] ), .CO(
        \mult_22/CARRYB[31][51] ), .S(\mult_22/SUMB[31][51] ) );
  FA_X1 \mult_22/S2_31_50  ( .A(\mult_22/ab[31][50] ), .B(
        \mult_22/CARRYB[30][50] ), .CI(\mult_22/SUMB[30][51] ), .CO(
        \mult_22/CARRYB[31][50] ), .S(\mult_22/SUMB[31][50] ) );
  FA_X1 \mult_22/S2_31_49  ( .A(\mult_22/ab[31][49] ), .B(
        \mult_22/CARRYB[30][49] ), .CI(\mult_22/SUMB[30][50] ), .CO(
        \mult_22/CARRYB[31][49] ), .S(\mult_22/SUMB[31][49] ) );
  FA_X1 \mult_22/S2_31_48  ( .A(\mult_22/ab[31][48] ), .B(
        \mult_22/CARRYB[30][48] ), .CI(\mult_22/SUMB[30][49] ), .CO(
        \mult_22/CARRYB[31][48] ), .S(\mult_22/SUMB[31][48] ) );
  FA_X1 \mult_22/S2_31_47  ( .A(\mult_22/ab[31][47] ), .B(
        \mult_22/CARRYB[30][47] ), .CI(\mult_22/SUMB[30][48] ), .CO(
        \mult_22/CARRYB[31][47] ), .S(\mult_22/SUMB[31][47] ) );
  FA_X1 \mult_22/S2_31_46  ( .A(\mult_22/ab[31][46] ), .B(
        \mult_22/CARRYB[30][46] ), .CI(\mult_22/SUMB[30][47] ), .CO(
        \mult_22/CARRYB[31][46] ), .S(\mult_22/SUMB[31][46] ) );
  FA_X1 \mult_22/S2_31_45  ( .A(\mult_22/ab[31][45] ), .B(
        \mult_22/CARRYB[30][45] ), .CI(\mult_22/SUMB[30][46] ), .CO(
        \mult_22/CARRYB[31][45] ), .S(\mult_22/SUMB[31][45] ) );
  FA_X1 \mult_22/S2_31_44  ( .A(\mult_22/ab[31][44] ), .B(
        \mult_22/CARRYB[30][44] ), .CI(\mult_22/SUMB[30][45] ), .CO(
        \mult_22/CARRYB[31][44] ), .S(\mult_22/SUMB[31][44] ) );
  FA_X1 \mult_22/S2_31_43  ( .A(\mult_22/ab[31][43] ), .B(
        \mult_22/CARRYB[30][43] ), .CI(\mult_22/SUMB[30][44] ), .CO(
        \mult_22/CARRYB[31][43] ), .S(\mult_22/SUMB[31][43] ) );
  FA_X1 \mult_22/S2_31_42  ( .A(\mult_22/ab[31][42] ), .B(
        \mult_22/CARRYB[30][42] ), .CI(\mult_22/SUMB[30][43] ), .CO(
        \mult_22/CARRYB[31][42] ), .S(\mult_22/SUMB[31][42] ) );
  FA_X1 \mult_22/S2_31_41  ( .A(\mult_22/ab[31][41] ), .B(
        \mult_22/CARRYB[30][41] ), .CI(\mult_22/SUMB[30][42] ), .CO(
        \mult_22/CARRYB[31][41] ), .S(\mult_22/SUMB[31][41] ) );
  FA_X1 \mult_22/S2_31_40  ( .A(\mult_22/ab[31][40] ), .B(
        \mult_22/CARRYB[30][40] ), .CI(\mult_22/SUMB[30][41] ), .CO(
        \mult_22/CARRYB[31][40] ), .S(\mult_22/SUMB[31][40] ) );
  FA_X1 \mult_22/S2_31_39  ( .A(\mult_22/ab[31][39] ), .B(
        \mult_22/CARRYB[30][39] ), .CI(\mult_22/SUMB[30][40] ), .CO(
        \mult_22/CARRYB[31][39] ), .S(\mult_22/SUMB[31][39] ) );
  FA_X1 \mult_22/S2_31_38  ( .A(\mult_22/ab[31][38] ), .B(
        \mult_22/CARRYB[30][38] ), .CI(\mult_22/SUMB[30][39] ), .CO(
        \mult_22/CARRYB[31][38] ), .S(\mult_22/SUMB[31][38] ) );
  FA_X1 \mult_22/S2_31_37  ( .A(\mult_22/ab[31][37] ), .B(
        \mult_22/CARRYB[30][37] ), .CI(\mult_22/SUMB[30][38] ), .CO(
        \mult_22/CARRYB[31][37] ), .S(\mult_22/SUMB[31][37] ) );
  FA_X1 \mult_22/S2_31_36  ( .A(\mult_22/ab[31][36] ), .B(
        \mult_22/CARRYB[30][36] ), .CI(\mult_22/SUMB[30][37] ), .CO(
        \mult_22/CARRYB[31][36] ), .S(\mult_22/SUMB[31][36] ) );
  FA_X1 \mult_22/S2_31_35  ( .A(\mult_22/ab[31][35] ), .B(
        \mult_22/CARRYB[30][35] ), .CI(\mult_22/SUMB[30][36] ), .CO(
        \mult_22/CARRYB[31][35] ), .S(\mult_22/SUMB[31][35] ) );
  FA_X1 \mult_22/S2_31_34  ( .A(\mult_22/ab[31][34] ), .B(
        \mult_22/CARRYB[30][34] ), .CI(\mult_22/SUMB[30][35] ), .CO(
        \mult_22/CARRYB[31][34] ), .S(\mult_22/SUMB[31][34] ) );
  FA_X1 \mult_22/S2_31_33  ( .A(\mult_22/ab[31][33] ), .B(
        \mult_22/CARRYB[30][33] ), .CI(\mult_22/SUMB[30][34] ), .CO(
        \mult_22/CARRYB[31][33] ), .S(\mult_22/SUMB[31][33] ) );
  FA_X1 \mult_22/S2_31_32  ( .A(\mult_22/ab[31][32] ), .B(
        \mult_22/CARRYB[30][32] ), .CI(\mult_22/SUMB[30][33] ), .CO(
        \mult_22/CARRYB[31][32] ), .S(\mult_22/SUMB[31][32] ) );
  FA_X1 \mult_22/S2_31_30  ( .A(\mult_22/CARRYB[30][30] ), .B(
        \mult_22/ab[31][30] ), .CI(\mult_22/SUMB[30][31] ), .CO(
        \mult_22/CARRYB[31][30] ), .S(\mult_22/SUMB[31][30] ) );
  FA_X1 \mult_22/S2_31_29  ( .A(\mult_22/ab[31][29] ), .B(
        \mult_22/CARRYB[30][29] ), .CI(\mult_22/SUMB[30][30] ), .CO(
        \mult_22/CARRYB[31][29] ), .S(\mult_22/SUMB[31][29] ) );
  FA_X1 \mult_22/S2_31_28  ( .A(\mult_22/ab[31][28] ), .B(
        \mult_22/CARRYB[30][28] ), .CI(\mult_22/SUMB[30][29] ), .CO(
        \mult_22/CARRYB[31][28] ), .S(\mult_22/SUMB[31][28] ) );
  FA_X1 \mult_22/S2_31_27  ( .A(\mult_22/ab[31][27] ), .B(
        \mult_22/CARRYB[30][27] ), .CI(\mult_22/SUMB[30][28] ), .CO(
        \mult_22/CARRYB[31][27] ), .S(\mult_22/SUMB[31][27] ) );
  FA_X1 \mult_22/S2_31_26  ( .A(\mult_22/ab[31][26] ), .B(
        \mult_22/CARRYB[30][26] ), .CI(\mult_22/SUMB[30][27] ), .CO(
        \mult_22/CARRYB[31][26] ), .S(\mult_22/SUMB[31][26] ) );
  FA_X1 \mult_22/S2_31_25  ( .A(\mult_22/ab[31][25] ), .B(
        \mult_22/CARRYB[30][25] ), .CI(\mult_22/SUMB[30][26] ), .CO(
        \mult_22/CARRYB[31][25] ), .S(\mult_22/SUMB[31][25] ) );
  FA_X1 \mult_22/S2_31_24  ( .A(\mult_22/ab[31][24] ), .B(
        \mult_22/CARRYB[30][24] ), .CI(\mult_22/SUMB[30][25] ), .CO(
        \mult_22/CARRYB[31][24] ), .S(\mult_22/SUMB[31][24] ) );
  FA_X1 \mult_22/S2_31_23  ( .A(\mult_22/ab[31][23] ), .B(
        \mult_22/CARRYB[30][23] ), .CI(\mult_22/SUMB[30][24] ), .CO(
        \mult_22/CARRYB[31][23] ), .S(\mult_22/SUMB[31][23] ) );
  FA_X1 \mult_22/S2_31_22  ( .A(\mult_22/ab[31][22] ), .B(
        \mult_22/CARRYB[30][22] ), .CI(\mult_22/SUMB[30][23] ), .CO(
        \mult_22/CARRYB[31][22] ), .S(\mult_22/SUMB[31][22] ) );
  FA_X1 \mult_22/S2_31_21  ( .A(\mult_22/ab[31][21] ), .B(
        \mult_22/CARRYB[30][21] ), .CI(\mult_22/SUMB[30][22] ), .CO(
        \mult_22/CARRYB[31][21] ), .S(\mult_22/SUMB[31][21] ) );
  FA_X1 \mult_22/S2_31_20  ( .A(\mult_22/ab[31][20] ), .B(
        \mult_22/CARRYB[30][20] ), .CI(\mult_22/SUMB[30][21] ), .CO(
        \mult_22/CARRYB[31][20] ), .S(\mult_22/SUMB[31][20] ) );
  FA_X1 \mult_22/S2_31_19  ( .A(\mult_22/ab[31][19] ), .B(
        \mult_22/CARRYB[30][19] ), .CI(\mult_22/SUMB[30][20] ), .CO(
        \mult_22/CARRYB[31][19] ), .S(\mult_22/SUMB[31][19] ) );
  FA_X1 \mult_22/S2_31_18  ( .A(\mult_22/ab[31][18] ), .B(
        \mult_22/CARRYB[30][18] ), .CI(\mult_22/SUMB[30][19] ), .CO(
        \mult_22/CARRYB[31][18] ), .S(\mult_22/SUMB[31][18] ) );
  FA_X1 \mult_22/S2_31_17  ( .A(\mult_22/ab[31][17] ), .B(
        \mult_22/CARRYB[30][17] ), .CI(\mult_22/SUMB[30][18] ), .CO(
        \mult_22/CARRYB[31][17] ), .S(\mult_22/SUMB[31][17] ) );
  FA_X1 \mult_22/S2_31_16  ( .A(\mult_22/ab[31][16] ), .B(
        \mult_22/CARRYB[30][16] ), .CI(\mult_22/SUMB[30][17] ), .CO(
        \mult_22/CARRYB[31][16] ), .S(\mult_22/SUMB[31][16] ) );
  FA_X1 \mult_22/S2_31_15  ( .A(\mult_22/ab[31][15] ), .B(
        \mult_22/CARRYB[30][15] ), .CI(\mult_22/SUMB[30][16] ), .CO(
        \mult_22/CARRYB[31][15] ), .S(\mult_22/SUMB[31][15] ) );
  FA_X1 \mult_22/S2_31_14  ( .A(\mult_22/ab[31][14] ), .B(
        \mult_22/CARRYB[30][14] ), .CI(\mult_22/SUMB[30][15] ), .CO(
        \mult_22/CARRYB[31][14] ), .S(\mult_22/SUMB[31][14] ) );
  FA_X1 \mult_22/S2_31_13  ( .A(\mult_22/ab[31][13] ), .B(
        \mult_22/CARRYB[30][13] ), .CI(\mult_22/SUMB[30][14] ), .CO(
        \mult_22/CARRYB[31][13] ), .S(\mult_22/SUMB[31][13] ) );
  FA_X1 \mult_22/S2_31_12  ( .A(\mult_22/ab[31][12] ), .B(
        \mult_22/CARRYB[30][12] ), .CI(\mult_22/SUMB[30][13] ), .CO(
        \mult_22/CARRYB[31][12] ), .S(\mult_22/SUMB[31][12] ) );
  FA_X1 \mult_22/S2_31_11  ( .A(\mult_22/ab[31][11] ), .B(
        \mult_22/CARRYB[30][11] ), .CI(\mult_22/SUMB[30][12] ), .CO(
        \mult_22/CARRYB[31][11] ), .S(\mult_22/SUMB[31][11] ) );
  FA_X1 \mult_22/S2_31_10  ( .A(\mult_22/ab[31][10] ), .B(
        \mult_22/CARRYB[30][10] ), .CI(\mult_22/SUMB[30][11] ), .CO(
        \mult_22/CARRYB[31][10] ), .S(\mult_22/SUMB[31][10] ) );
  FA_X1 \mult_22/S2_31_9  ( .A(\mult_22/ab[31][9] ), .B(
        \mult_22/CARRYB[30][9] ), .CI(\mult_22/SUMB[30][10] ), .CO(
        \mult_22/CARRYB[31][9] ), .S(\mult_22/SUMB[31][9] ) );
  FA_X1 \mult_22/S2_31_8  ( .A(\mult_22/ab[31][8] ), .B(
        \mult_22/CARRYB[30][8] ), .CI(\mult_22/SUMB[30][9] ), .CO(
        \mult_22/CARRYB[31][8] ), .S(\mult_22/SUMB[31][8] ) );
  FA_X1 \mult_22/S2_31_7  ( .A(\mult_22/ab[31][7] ), .B(
        \mult_22/CARRYB[30][7] ), .CI(\mult_22/SUMB[30][8] ), .CO(
        \mult_22/CARRYB[31][7] ), .S(\mult_22/SUMB[31][7] ) );
  FA_X1 \mult_22/S2_31_6  ( .A(\mult_22/ab[31][6] ), .B(
        \mult_22/CARRYB[30][6] ), .CI(\mult_22/SUMB[30][7] ), .CO(
        \mult_22/CARRYB[31][6] ), .S(\mult_22/SUMB[31][6] ) );
  FA_X1 \mult_22/S2_31_5  ( .A(\mult_22/ab[31][5] ), .B(
        \mult_22/CARRYB[30][5] ), .CI(\mult_22/SUMB[30][6] ), .CO(
        \mult_22/CARRYB[31][5] ), .S(\mult_22/SUMB[31][5] ) );
  FA_X1 \mult_22/S2_31_4  ( .A(\mult_22/ab[31][4] ), .B(
        \mult_22/CARRYB[30][4] ), .CI(\mult_22/SUMB[30][5] ), .CO(
        \mult_22/CARRYB[31][4] ), .S(\mult_22/SUMB[31][4] ) );
  FA_X1 \mult_22/S2_31_3  ( .A(\mult_22/ab[31][3] ), .B(
        \mult_22/CARRYB[30][3] ), .CI(\mult_22/SUMB[30][4] ), .CO(
        \mult_22/CARRYB[31][3] ), .S(\mult_22/SUMB[31][3] ) );
  FA_X1 \mult_22/S2_31_2  ( .A(\mult_22/ab[31][2] ), .B(
        \mult_22/CARRYB[30][2] ), .CI(\mult_22/SUMB[30][3] ), .CO(
        \mult_22/CARRYB[31][2] ), .S(\mult_22/SUMB[31][2] ) );
  FA_X1 \mult_22/S2_31_1  ( .A(\mult_22/ab[31][1] ), .B(
        \mult_22/CARRYB[30][1] ), .CI(\mult_22/SUMB[30][2] ), .CO(
        \mult_22/CARRYB[31][1] ), .S(\mult_22/SUMB[31][1] ) );
  FA_X1 \mult_22/S1_31_0  ( .A(\mult_22/ab[31][0] ), .B(
        \mult_22/CARRYB[30][0] ), .CI(\mult_22/SUMB[30][1] ), .CO(
        \mult_22/CARRYB[31][0] ), .S(N159) );
  FA_X1 \mult_22/S3_32_62  ( .A(\mult_22/ab[32][62] ), .B(
        \mult_22/CARRYB[31][62] ), .CI(\mult_22/ab[31][63] ), .CO(
        \mult_22/CARRYB[32][62] ), .S(\mult_22/SUMB[32][62] ) );
  FA_X1 \mult_22/S2_32_61  ( .A(\mult_22/ab[32][61] ), .B(
        \mult_22/CARRYB[31][61] ), .CI(\mult_22/SUMB[31][62] ), .CO(
        \mult_22/CARRYB[32][61] ), .S(\mult_22/SUMB[32][61] ) );
  FA_X1 \mult_22/S2_32_60  ( .A(\mult_22/ab[32][60] ), .B(
        \mult_22/CARRYB[31][60] ), .CI(\mult_22/SUMB[31][61] ), .CO(
        \mult_22/CARRYB[32][60] ), .S(\mult_22/SUMB[32][60] ) );
  FA_X1 \mult_22/S2_32_59  ( .A(\mult_22/ab[32][59] ), .B(
        \mult_22/CARRYB[31][59] ), .CI(\mult_22/SUMB[31][60] ), .CO(
        \mult_22/CARRYB[32][59] ), .S(\mult_22/SUMB[32][59] ) );
  FA_X1 \mult_22/S2_32_58  ( .A(\mult_22/ab[32][58] ), .B(
        \mult_22/CARRYB[31][58] ), .CI(\mult_22/SUMB[31][59] ), .CO(
        \mult_22/CARRYB[32][58] ), .S(\mult_22/SUMB[32][58] ) );
  FA_X1 \mult_22/S2_32_57  ( .A(\mult_22/ab[32][57] ), .B(
        \mult_22/CARRYB[31][57] ), .CI(\mult_22/SUMB[31][58] ), .CO(
        \mult_22/CARRYB[32][57] ), .S(\mult_22/SUMB[32][57] ) );
  FA_X1 \mult_22/S2_32_56  ( .A(\mult_22/ab[32][56] ), .B(
        \mult_22/CARRYB[31][56] ), .CI(\mult_22/SUMB[31][57] ), .CO(
        \mult_22/CARRYB[32][56] ), .S(\mult_22/SUMB[32][56] ) );
  FA_X1 \mult_22/S2_32_55  ( .A(\mult_22/ab[32][55] ), .B(
        \mult_22/CARRYB[31][55] ), .CI(\mult_22/SUMB[31][56] ), .CO(
        \mult_22/CARRYB[32][55] ), .S(\mult_22/SUMB[32][55] ) );
  FA_X1 \mult_22/S2_32_54  ( .A(\mult_22/ab[32][54] ), .B(
        \mult_22/CARRYB[31][54] ), .CI(\mult_22/SUMB[31][55] ), .CO(
        \mult_22/CARRYB[32][54] ), .S(\mult_22/SUMB[32][54] ) );
  FA_X1 \mult_22/S2_32_53  ( .A(\mult_22/ab[32][53] ), .B(
        \mult_22/CARRYB[31][53] ), .CI(\mult_22/SUMB[31][54] ), .CO(
        \mult_22/CARRYB[32][53] ), .S(\mult_22/SUMB[32][53] ) );
  FA_X1 \mult_22/S2_32_52  ( .A(\mult_22/ab[32][52] ), .B(
        \mult_22/CARRYB[31][52] ), .CI(\mult_22/SUMB[31][53] ), .CO(
        \mult_22/CARRYB[32][52] ), .S(\mult_22/SUMB[32][52] ) );
  FA_X1 \mult_22/S2_32_51  ( .A(\mult_22/ab[32][51] ), .B(
        \mult_22/CARRYB[31][51] ), .CI(\mult_22/SUMB[31][52] ), .CO(
        \mult_22/CARRYB[32][51] ), .S(\mult_22/SUMB[32][51] ) );
  FA_X1 \mult_22/S2_32_50  ( .A(\mult_22/ab[32][50] ), .B(
        \mult_22/CARRYB[31][50] ), .CI(\mult_22/SUMB[31][51] ), .CO(
        \mult_22/CARRYB[32][50] ), .S(\mult_22/SUMB[32][50] ) );
  FA_X1 \mult_22/S2_32_49  ( .A(\mult_22/ab[32][49] ), .B(
        \mult_22/CARRYB[31][49] ), .CI(\mult_22/SUMB[31][50] ), .CO(
        \mult_22/CARRYB[32][49] ), .S(\mult_22/SUMB[32][49] ) );
  FA_X1 \mult_22/S2_32_48  ( .A(\mult_22/ab[32][48] ), .B(
        \mult_22/CARRYB[31][48] ), .CI(\mult_22/SUMB[31][49] ), .CO(
        \mult_22/CARRYB[32][48] ), .S(\mult_22/SUMB[32][48] ) );
  FA_X1 \mult_22/S2_32_47  ( .A(\mult_22/ab[32][47] ), .B(
        \mult_22/CARRYB[31][47] ), .CI(\mult_22/SUMB[31][48] ), .CO(
        \mult_22/CARRYB[32][47] ), .S(\mult_22/SUMB[32][47] ) );
  FA_X1 \mult_22/S2_32_46  ( .A(\mult_22/ab[32][46] ), .B(
        \mult_22/CARRYB[31][46] ), .CI(\mult_22/SUMB[31][47] ), .CO(
        \mult_22/CARRYB[32][46] ), .S(\mult_22/SUMB[32][46] ) );
  FA_X1 \mult_22/S2_32_45  ( .A(\mult_22/ab[32][45] ), .B(
        \mult_22/CARRYB[31][45] ), .CI(\mult_22/SUMB[31][46] ), .CO(
        \mult_22/CARRYB[32][45] ), .S(\mult_22/SUMB[32][45] ) );
  FA_X1 \mult_22/S2_32_44  ( .A(\mult_22/ab[32][44] ), .B(
        \mult_22/CARRYB[31][44] ), .CI(\mult_22/SUMB[31][45] ), .CO(
        \mult_22/CARRYB[32][44] ), .S(\mult_22/SUMB[32][44] ) );
  FA_X1 \mult_22/S2_32_43  ( .A(\mult_22/ab[32][43] ), .B(
        \mult_22/CARRYB[31][43] ), .CI(\mult_22/SUMB[31][44] ), .CO(
        \mult_22/CARRYB[32][43] ), .S(\mult_22/SUMB[32][43] ) );
  FA_X1 \mult_22/S2_32_42  ( .A(\mult_22/ab[32][42] ), .B(
        \mult_22/CARRYB[31][42] ), .CI(\mult_22/SUMB[31][43] ), .CO(
        \mult_22/CARRYB[32][42] ), .S(\mult_22/SUMB[32][42] ) );
  FA_X1 \mult_22/S2_32_41  ( .A(\mult_22/ab[32][41] ), .B(
        \mult_22/CARRYB[31][41] ), .CI(\mult_22/SUMB[31][42] ), .CO(
        \mult_22/CARRYB[32][41] ), .S(\mult_22/SUMB[32][41] ) );
  FA_X1 \mult_22/S2_32_40  ( .A(\mult_22/ab[32][40] ), .B(
        \mult_22/CARRYB[31][40] ), .CI(\mult_22/SUMB[31][41] ), .CO(
        \mult_22/CARRYB[32][40] ), .S(\mult_22/SUMB[32][40] ) );
  FA_X1 \mult_22/S2_32_39  ( .A(\mult_22/ab[32][39] ), .B(
        \mult_22/CARRYB[31][39] ), .CI(\mult_22/SUMB[31][40] ), .CO(
        \mult_22/CARRYB[32][39] ), .S(\mult_22/SUMB[32][39] ) );
  FA_X1 \mult_22/S2_32_38  ( .A(\mult_22/ab[32][38] ), .B(
        \mult_22/CARRYB[31][38] ), .CI(\mult_22/SUMB[31][39] ), .CO(
        \mult_22/CARRYB[32][38] ), .S(\mult_22/SUMB[32][38] ) );
  FA_X1 \mult_22/S2_32_37  ( .A(\mult_22/ab[32][37] ), .B(
        \mult_22/CARRYB[31][37] ), .CI(\mult_22/SUMB[31][38] ), .CO(
        \mult_22/CARRYB[32][37] ), .S(\mult_22/SUMB[32][37] ) );
  FA_X1 \mult_22/S2_32_36  ( .A(\mult_22/ab[32][36] ), .B(
        \mult_22/CARRYB[31][36] ), .CI(\mult_22/SUMB[31][37] ), .CO(
        \mult_22/CARRYB[32][36] ), .S(\mult_22/SUMB[32][36] ) );
  FA_X1 \mult_22/S2_32_35  ( .A(\mult_22/ab[32][35] ), .B(
        \mult_22/CARRYB[31][35] ), .CI(\mult_22/SUMB[31][36] ), .CO(
        \mult_22/CARRYB[32][35] ), .S(\mult_22/SUMB[32][35] ) );
  FA_X1 \mult_22/S2_32_34  ( .A(\mult_22/CARRYB[31][34] ), .B(
        \mult_22/ab[32][34] ), .CI(\mult_22/SUMB[31][35] ), .CO(
        \mult_22/CARRYB[32][34] ), .S(\mult_22/SUMB[32][34] ) );
  FA_X1 \mult_22/S2_32_33  ( .A(\mult_22/ab[32][33] ), .B(
        \mult_22/CARRYB[31][33] ), .CI(\mult_22/SUMB[31][34] ), .CO(
        \mult_22/CARRYB[32][33] ), .S(\mult_22/SUMB[32][33] ) );
  FA_X1 \mult_22/S2_32_32  ( .A(\mult_22/ab[32][32] ), .B(
        \mult_22/CARRYB[31][32] ), .CI(\mult_22/SUMB[31][33] ), .CO(
        \mult_22/CARRYB[32][32] ), .S(\mult_22/SUMB[32][32] ) );
  FA_X1 \mult_22/S2_32_31  ( .A(\mult_22/ab[32][31] ), .B(
        \mult_22/CARRYB[31][31] ), .CI(\mult_22/SUMB[31][32] ), .CO(
        \mult_22/CARRYB[32][31] ), .S(\mult_22/SUMB[32][31] ) );
  FA_X1 \mult_22/S2_32_30  ( .A(\mult_22/ab[32][30] ), .B(
        \mult_22/CARRYB[31][30] ), .CI(\mult_22/SUMB[31][31] ), .CO(
        \mult_22/CARRYB[32][30] ), .S(\mult_22/SUMB[32][30] ) );
  FA_X1 \mult_22/S2_32_28  ( .A(\mult_22/ab[32][28] ), .B(
        \mult_22/CARRYB[31][28] ), .CI(\mult_22/SUMB[31][29] ), .CO(
        \mult_22/CARRYB[32][28] ), .S(\mult_22/SUMB[32][28] ) );
  FA_X1 \mult_22/S2_32_27  ( .A(\mult_22/ab[32][27] ), .B(
        \mult_22/CARRYB[31][27] ), .CI(\mult_22/SUMB[31][28] ), .CO(
        \mult_22/CARRYB[32][27] ), .S(\mult_22/SUMB[32][27] ) );
  FA_X1 \mult_22/S2_32_26  ( .A(\mult_22/ab[32][26] ), .B(
        \mult_22/CARRYB[31][26] ), .CI(\mult_22/SUMB[31][27] ), .CO(
        \mult_22/CARRYB[32][26] ), .S(\mult_22/SUMB[32][26] ) );
  FA_X1 \mult_22/S2_32_25  ( .A(\mult_22/ab[32][25] ), .B(
        \mult_22/CARRYB[31][25] ), .CI(\mult_22/SUMB[31][26] ), .CO(
        \mult_22/CARRYB[32][25] ), .S(\mult_22/SUMB[32][25] ) );
  FA_X1 \mult_22/S2_32_24  ( .A(\mult_22/ab[32][24] ), .B(
        \mult_22/CARRYB[31][24] ), .CI(\mult_22/SUMB[31][25] ), .CO(
        \mult_22/CARRYB[32][24] ), .S(\mult_22/SUMB[32][24] ) );
  FA_X1 \mult_22/S2_32_23  ( .A(\mult_22/ab[32][23] ), .B(
        \mult_22/CARRYB[31][23] ), .CI(\mult_22/SUMB[31][24] ), .CO(
        \mult_22/CARRYB[32][23] ), .S(\mult_22/SUMB[32][23] ) );
  FA_X1 \mult_22/S2_32_22  ( .A(\mult_22/ab[32][22] ), .B(
        \mult_22/CARRYB[31][22] ), .CI(\mult_22/SUMB[31][23] ), .CO(
        \mult_22/CARRYB[32][22] ), .S(\mult_22/SUMB[32][22] ) );
  FA_X1 \mult_22/S2_32_21  ( .A(\mult_22/ab[32][21] ), .B(
        \mult_22/CARRYB[31][21] ), .CI(\mult_22/SUMB[31][22] ), .CO(
        \mult_22/CARRYB[32][21] ), .S(\mult_22/SUMB[32][21] ) );
  FA_X1 \mult_22/S2_32_20  ( .A(\mult_22/ab[32][20] ), .B(
        \mult_22/CARRYB[31][20] ), .CI(\mult_22/SUMB[31][21] ), .CO(
        \mult_22/CARRYB[32][20] ), .S(\mult_22/SUMB[32][20] ) );
  FA_X1 \mult_22/S2_32_19  ( .A(\mult_22/ab[32][19] ), .B(
        \mult_22/CARRYB[31][19] ), .CI(\mult_22/SUMB[31][20] ), .CO(
        \mult_22/CARRYB[32][19] ), .S(\mult_22/SUMB[32][19] ) );
  FA_X1 \mult_22/S2_32_18  ( .A(\mult_22/ab[32][18] ), .B(
        \mult_22/CARRYB[31][18] ), .CI(\mult_22/SUMB[31][19] ), .CO(
        \mult_22/CARRYB[32][18] ), .S(\mult_22/SUMB[32][18] ) );
  FA_X1 \mult_22/S2_32_17  ( .A(\mult_22/ab[32][17] ), .B(
        \mult_22/CARRYB[31][17] ), .CI(\mult_22/SUMB[31][18] ), .CO(
        \mult_22/CARRYB[32][17] ), .S(\mult_22/SUMB[32][17] ) );
  FA_X1 \mult_22/S2_32_16  ( .A(\mult_22/ab[32][16] ), .B(
        \mult_22/CARRYB[31][16] ), .CI(\mult_22/SUMB[31][17] ), .CO(
        \mult_22/CARRYB[32][16] ), .S(\mult_22/SUMB[32][16] ) );
  FA_X1 \mult_22/S2_32_15  ( .A(\mult_22/ab[32][15] ), .B(
        \mult_22/CARRYB[31][15] ), .CI(\mult_22/SUMB[31][16] ), .CO(
        \mult_22/CARRYB[32][15] ), .S(\mult_22/SUMB[32][15] ) );
  FA_X1 \mult_22/S2_32_14  ( .A(\mult_22/ab[32][14] ), .B(
        \mult_22/CARRYB[31][14] ), .CI(\mult_22/SUMB[31][15] ), .CO(
        \mult_22/CARRYB[32][14] ), .S(\mult_22/SUMB[32][14] ) );
  FA_X1 \mult_22/S2_32_13  ( .A(\mult_22/ab[32][13] ), .B(
        \mult_22/CARRYB[31][13] ), .CI(\mult_22/SUMB[31][14] ), .CO(
        \mult_22/CARRYB[32][13] ), .S(\mult_22/SUMB[32][13] ) );
  FA_X1 \mult_22/S2_32_12  ( .A(\mult_22/ab[32][12] ), .B(
        \mult_22/CARRYB[31][12] ), .CI(\mult_22/SUMB[31][13] ), .CO(
        \mult_22/CARRYB[32][12] ), .S(\mult_22/SUMB[32][12] ) );
  FA_X1 \mult_22/S2_32_11  ( .A(\mult_22/ab[32][11] ), .B(
        \mult_22/CARRYB[31][11] ), .CI(\mult_22/SUMB[31][12] ), .CO(
        \mult_22/CARRYB[32][11] ), .S(\mult_22/SUMB[32][11] ) );
  FA_X1 \mult_22/S2_32_10  ( .A(\mult_22/ab[32][10] ), .B(
        \mult_22/CARRYB[31][10] ), .CI(\mult_22/SUMB[31][11] ), .CO(
        \mult_22/CARRYB[32][10] ), .S(\mult_22/SUMB[32][10] ) );
  FA_X1 \mult_22/S2_32_9  ( .A(\mult_22/ab[32][9] ), .B(
        \mult_22/CARRYB[31][9] ), .CI(\mult_22/SUMB[31][10] ), .CO(
        \mult_22/CARRYB[32][9] ), .S(\mult_22/SUMB[32][9] ) );
  FA_X1 \mult_22/S2_32_8  ( .A(\mult_22/ab[32][8] ), .B(
        \mult_22/CARRYB[31][8] ), .CI(\mult_22/SUMB[31][9] ), .CO(
        \mult_22/CARRYB[32][8] ), .S(\mult_22/SUMB[32][8] ) );
  FA_X1 \mult_22/S2_32_7  ( .A(\mult_22/ab[32][7] ), .B(
        \mult_22/CARRYB[31][7] ), .CI(\mult_22/SUMB[31][8] ), .CO(
        \mult_22/CARRYB[32][7] ), .S(\mult_22/SUMB[32][7] ) );
  FA_X1 \mult_22/S2_32_6  ( .A(\mult_22/ab[32][6] ), .B(
        \mult_22/CARRYB[31][6] ), .CI(\mult_22/SUMB[31][7] ), .CO(
        \mult_22/CARRYB[32][6] ), .S(\mult_22/SUMB[32][6] ) );
  FA_X1 \mult_22/S2_32_5  ( .A(\mult_22/ab[32][5] ), .B(
        \mult_22/CARRYB[31][5] ), .CI(\mult_22/SUMB[31][6] ), .CO(
        \mult_22/CARRYB[32][5] ), .S(\mult_22/SUMB[32][5] ) );
  FA_X1 \mult_22/S2_32_4  ( .A(\mult_22/ab[32][4] ), .B(
        \mult_22/CARRYB[31][4] ), .CI(\mult_22/SUMB[31][5] ), .CO(
        \mult_22/CARRYB[32][4] ), .S(\mult_22/SUMB[32][4] ) );
  FA_X1 \mult_22/S2_32_3  ( .A(\mult_22/ab[32][3] ), .B(
        \mult_22/CARRYB[31][3] ), .CI(\mult_22/SUMB[31][4] ), .CO(
        \mult_22/CARRYB[32][3] ), .S(\mult_22/SUMB[32][3] ) );
  FA_X1 \mult_22/S2_32_2  ( .A(\mult_22/ab[32][2] ), .B(
        \mult_22/CARRYB[31][2] ), .CI(\mult_22/SUMB[31][3] ), .CO(
        \mult_22/CARRYB[32][2] ), .S(\mult_22/SUMB[32][2] ) );
  FA_X1 \mult_22/S2_32_1  ( .A(\mult_22/ab[32][1] ), .B(
        \mult_22/CARRYB[31][1] ), .CI(\mult_22/SUMB[31][2] ), .CO(
        \mult_22/CARRYB[32][1] ), .S(\mult_22/SUMB[32][1] ) );
  FA_X1 \mult_22/S1_32_0  ( .A(\mult_22/ab[32][0] ), .B(
        \mult_22/CARRYB[31][0] ), .CI(\mult_22/SUMB[31][1] ), .CO(
        \mult_22/CARRYB[32][0] ), .S(N160) );
  FA_X1 \mult_22/S3_33_62  ( .A(\mult_22/ab[33][62] ), .B(
        \mult_22/CARRYB[32][62] ), .CI(\mult_22/ab[32][63] ), .CO(
        \mult_22/CARRYB[33][62] ), .S(\mult_22/SUMB[33][62] ) );
  FA_X1 \mult_22/S2_33_61  ( .A(\mult_22/ab[33][61] ), .B(
        \mult_22/CARRYB[32][61] ), .CI(\mult_22/SUMB[32][62] ), .CO(
        \mult_22/CARRYB[33][61] ), .S(\mult_22/SUMB[33][61] ) );
  FA_X1 \mult_22/S2_33_60  ( .A(\mult_22/ab[33][60] ), .B(
        \mult_22/CARRYB[32][60] ), .CI(\mult_22/SUMB[32][61] ), .CO(
        \mult_22/CARRYB[33][60] ), .S(\mult_22/SUMB[33][60] ) );
  FA_X1 \mult_22/S2_33_59  ( .A(\mult_22/ab[33][59] ), .B(
        \mult_22/CARRYB[32][59] ), .CI(\mult_22/SUMB[32][60] ), .CO(
        \mult_22/CARRYB[33][59] ), .S(\mult_22/SUMB[33][59] ) );
  FA_X1 \mult_22/S2_33_58  ( .A(\mult_22/ab[33][58] ), .B(
        \mult_22/CARRYB[32][58] ), .CI(\mult_22/SUMB[32][59] ), .CO(
        \mult_22/CARRYB[33][58] ), .S(\mult_22/SUMB[33][58] ) );
  FA_X1 \mult_22/S2_33_57  ( .A(\mult_22/ab[33][57] ), .B(
        \mult_22/CARRYB[32][57] ), .CI(\mult_22/SUMB[32][58] ), .CO(
        \mult_22/CARRYB[33][57] ), .S(\mult_22/SUMB[33][57] ) );
  FA_X1 \mult_22/S2_33_56  ( .A(\mult_22/ab[33][56] ), .B(
        \mult_22/CARRYB[32][56] ), .CI(\mult_22/SUMB[32][57] ), .CO(
        \mult_22/CARRYB[33][56] ), .S(\mult_22/SUMB[33][56] ) );
  FA_X1 \mult_22/S2_33_55  ( .A(\mult_22/ab[33][55] ), .B(
        \mult_22/CARRYB[32][55] ), .CI(\mult_22/SUMB[32][56] ), .CO(
        \mult_22/CARRYB[33][55] ), .S(\mult_22/SUMB[33][55] ) );
  FA_X1 \mult_22/S2_33_54  ( .A(\mult_22/ab[33][54] ), .B(
        \mult_22/CARRYB[32][54] ), .CI(\mult_22/SUMB[32][55] ), .CO(
        \mult_22/CARRYB[33][54] ), .S(\mult_22/SUMB[33][54] ) );
  FA_X1 \mult_22/S2_33_53  ( .A(\mult_22/ab[33][53] ), .B(
        \mult_22/CARRYB[32][53] ), .CI(\mult_22/SUMB[32][54] ), .CO(
        \mult_22/CARRYB[33][53] ), .S(\mult_22/SUMB[33][53] ) );
  FA_X1 \mult_22/S2_33_52  ( .A(\mult_22/ab[33][52] ), .B(
        \mult_22/CARRYB[32][52] ), .CI(\mult_22/SUMB[32][53] ), .CO(
        \mult_22/CARRYB[33][52] ), .S(\mult_22/SUMB[33][52] ) );
  FA_X1 \mult_22/S2_33_51  ( .A(\mult_22/ab[33][51] ), .B(
        \mult_22/CARRYB[32][51] ), .CI(\mult_22/SUMB[32][52] ), .CO(
        \mult_22/CARRYB[33][51] ), .S(\mult_22/SUMB[33][51] ) );
  FA_X1 \mult_22/S2_33_50  ( .A(\mult_22/ab[33][50] ), .B(
        \mult_22/CARRYB[32][50] ), .CI(\mult_22/SUMB[32][51] ), .CO(
        \mult_22/CARRYB[33][50] ), .S(\mult_22/SUMB[33][50] ) );
  FA_X1 \mult_22/S2_33_49  ( .A(\mult_22/ab[33][49] ), .B(
        \mult_22/CARRYB[32][49] ), .CI(\mult_22/SUMB[32][50] ), .CO(
        \mult_22/CARRYB[33][49] ), .S(\mult_22/SUMB[33][49] ) );
  FA_X1 \mult_22/S2_33_48  ( .A(\mult_22/ab[33][48] ), .B(
        \mult_22/CARRYB[32][48] ), .CI(\mult_22/SUMB[32][49] ), .CO(
        \mult_22/CARRYB[33][48] ), .S(\mult_22/SUMB[33][48] ) );
  FA_X1 \mult_22/S2_33_47  ( .A(\mult_22/ab[33][47] ), .B(
        \mult_22/CARRYB[32][47] ), .CI(\mult_22/SUMB[32][48] ), .CO(
        \mult_22/CARRYB[33][47] ), .S(\mult_22/SUMB[33][47] ) );
  FA_X1 \mult_22/S2_33_46  ( .A(\mult_22/ab[33][46] ), .B(
        \mult_22/CARRYB[32][46] ), .CI(\mult_22/SUMB[32][47] ), .CO(
        \mult_22/CARRYB[33][46] ), .S(\mult_22/SUMB[33][46] ) );
  FA_X1 \mult_22/S2_33_45  ( .A(\mult_22/ab[33][45] ), .B(
        \mult_22/CARRYB[32][45] ), .CI(\mult_22/SUMB[32][46] ), .CO(
        \mult_22/CARRYB[33][45] ), .S(\mult_22/SUMB[33][45] ) );
  FA_X1 \mult_22/S2_33_44  ( .A(\mult_22/ab[33][44] ), .B(
        \mult_22/CARRYB[32][44] ), .CI(\mult_22/SUMB[32][45] ), .CO(
        \mult_22/CARRYB[33][44] ), .S(\mult_22/SUMB[33][44] ) );
  FA_X1 \mult_22/S2_33_43  ( .A(\mult_22/ab[33][43] ), .B(
        \mult_22/CARRYB[32][43] ), .CI(\mult_22/SUMB[32][44] ), .CO(
        \mult_22/CARRYB[33][43] ), .S(\mult_22/SUMB[33][43] ) );
  FA_X1 \mult_22/S2_33_42  ( .A(\mult_22/ab[33][42] ), .B(
        \mult_22/CARRYB[32][42] ), .CI(\mult_22/SUMB[32][43] ), .CO(
        \mult_22/CARRYB[33][42] ), .S(\mult_22/SUMB[33][42] ) );
  FA_X1 \mult_22/S2_33_41  ( .A(\mult_22/ab[33][41] ), .B(
        \mult_22/CARRYB[32][41] ), .CI(\mult_22/SUMB[32][42] ), .CO(
        \mult_22/CARRYB[33][41] ), .S(\mult_22/SUMB[33][41] ) );
  FA_X1 \mult_22/S2_33_40  ( .A(\mult_22/ab[33][40] ), .B(
        \mult_22/CARRYB[32][40] ), .CI(\mult_22/SUMB[32][41] ), .CO(
        \mult_22/CARRYB[33][40] ), .S(\mult_22/SUMB[33][40] ) );
  FA_X1 \mult_22/S2_33_39  ( .A(\mult_22/ab[33][39] ), .B(
        \mult_22/CARRYB[32][39] ), .CI(\mult_22/SUMB[32][40] ), .CO(
        \mult_22/CARRYB[33][39] ), .S(\mult_22/SUMB[33][39] ) );
  FA_X1 \mult_22/S2_33_38  ( .A(\mult_22/ab[33][38] ), .B(
        \mult_22/CARRYB[32][38] ), .CI(\mult_22/SUMB[32][39] ), .CO(
        \mult_22/CARRYB[33][38] ), .S(\mult_22/SUMB[33][38] ) );
  FA_X1 \mult_22/S2_33_37  ( .A(\mult_22/ab[33][37] ), .B(
        \mult_22/CARRYB[32][37] ), .CI(\mult_22/SUMB[32][38] ), .CO(
        \mult_22/CARRYB[33][37] ), .S(\mult_22/SUMB[33][37] ) );
  FA_X1 \mult_22/S2_33_36  ( .A(\mult_22/ab[33][36] ), .B(
        \mult_22/CARRYB[32][36] ), .CI(\mult_22/SUMB[32][37] ), .CO(
        \mult_22/CARRYB[33][36] ), .S(\mult_22/SUMB[33][36] ) );
  FA_X1 \mult_22/S2_33_35  ( .A(\mult_22/ab[33][35] ), .B(
        \mult_22/CARRYB[32][35] ), .CI(\mult_22/SUMB[32][36] ), .CO(
        \mult_22/CARRYB[33][35] ), .S(\mult_22/SUMB[33][35] ) );
  FA_X1 \mult_22/S2_33_34  ( .A(\mult_22/ab[33][34] ), .B(
        \mult_22/CARRYB[32][34] ), .CI(\mult_22/SUMB[32][35] ), .CO(
        \mult_22/CARRYB[33][34] ), .S(\mult_22/SUMB[33][34] ) );
  FA_X1 \mult_22/S2_33_33  ( .A(\mult_22/ab[33][33] ), .B(
        \mult_22/CARRYB[32][33] ), .CI(\mult_22/SUMB[32][34] ), .CO(
        \mult_22/CARRYB[33][33] ), .S(\mult_22/SUMB[33][33] ) );
  FA_X1 \mult_22/S2_33_32  ( .A(\mult_22/ab[33][32] ), .B(
        \mult_22/CARRYB[32][32] ), .CI(\mult_22/SUMB[32][33] ), .CO(
        \mult_22/CARRYB[33][32] ), .S(\mult_22/SUMB[33][32] ) );
  FA_X1 \mult_22/S2_33_31  ( .A(\mult_22/ab[33][31] ), .B(
        \mult_22/CARRYB[32][31] ), .CI(\mult_22/SUMB[32][32] ), .CO(
        \mult_22/CARRYB[33][31] ), .S(\mult_22/SUMB[33][31] ) );
  FA_X1 \mult_22/S2_33_30  ( .A(\mult_22/ab[33][30] ), .B(
        \mult_22/CARRYB[32][30] ), .CI(\mult_22/SUMB[32][31] ), .CO(
        \mult_22/CARRYB[33][30] ), .S(\mult_22/SUMB[33][30] ) );
  FA_X1 \mult_22/S2_33_29  ( .A(\mult_22/ab[33][29] ), .B(
        \mult_22/CARRYB[32][29] ), .CI(\mult_22/SUMB[32][30] ), .CO(
        \mult_22/CARRYB[33][29] ), .S(\mult_22/SUMB[33][29] ) );
  FA_X1 \mult_22/S2_33_27  ( .A(\mult_22/ab[33][27] ), .B(
        \mult_22/CARRYB[32][27] ), .CI(\mult_22/SUMB[32][28] ), .CO(
        \mult_22/CARRYB[33][27] ), .S(\mult_22/SUMB[33][27] ) );
  FA_X1 \mult_22/S2_33_26  ( .A(\mult_22/ab[33][26] ), .B(
        \mult_22/CARRYB[32][26] ), .CI(\mult_22/SUMB[32][27] ), .CO(
        \mult_22/CARRYB[33][26] ), .S(\mult_22/SUMB[33][26] ) );
  FA_X1 \mult_22/S2_33_25  ( .A(\mult_22/ab[33][25] ), .B(
        \mult_22/CARRYB[32][25] ), .CI(\mult_22/SUMB[32][26] ), .CO(
        \mult_22/CARRYB[33][25] ), .S(\mult_22/SUMB[33][25] ) );
  FA_X1 \mult_22/S2_33_24  ( .A(\mult_22/ab[33][24] ), .B(
        \mult_22/CARRYB[32][24] ), .CI(\mult_22/SUMB[32][25] ), .CO(
        \mult_22/CARRYB[33][24] ), .S(\mult_22/SUMB[33][24] ) );
  FA_X1 \mult_22/S2_33_23  ( .A(\mult_22/ab[33][23] ), .B(
        \mult_22/CARRYB[32][23] ), .CI(\mult_22/SUMB[32][24] ), .CO(
        \mult_22/CARRYB[33][23] ), .S(\mult_22/SUMB[33][23] ) );
  FA_X1 \mult_22/S2_33_22  ( .A(\mult_22/ab[33][22] ), .B(
        \mult_22/CARRYB[32][22] ), .CI(\mult_22/SUMB[32][23] ), .CO(
        \mult_22/CARRYB[33][22] ), .S(\mult_22/SUMB[33][22] ) );
  FA_X1 \mult_22/S2_33_21  ( .A(\mult_22/ab[33][21] ), .B(
        \mult_22/CARRYB[32][21] ), .CI(\mult_22/SUMB[32][22] ), .CO(
        \mult_22/CARRYB[33][21] ), .S(\mult_22/SUMB[33][21] ) );
  FA_X1 \mult_22/S2_33_20  ( .A(\mult_22/ab[33][20] ), .B(
        \mult_22/CARRYB[32][20] ), .CI(\mult_22/SUMB[32][21] ), .CO(
        \mult_22/CARRYB[33][20] ), .S(\mult_22/SUMB[33][20] ) );
  FA_X1 \mult_22/S2_33_19  ( .A(\mult_22/ab[33][19] ), .B(
        \mult_22/CARRYB[32][19] ), .CI(\mult_22/SUMB[32][20] ), .CO(
        \mult_22/CARRYB[33][19] ), .S(\mult_22/SUMB[33][19] ) );
  FA_X1 \mult_22/S2_33_18  ( .A(\mult_22/ab[33][18] ), .B(
        \mult_22/CARRYB[32][18] ), .CI(\mult_22/SUMB[32][19] ), .CO(
        \mult_22/CARRYB[33][18] ), .S(\mult_22/SUMB[33][18] ) );
  FA_X1 \mult_22/S2_33_17  ( .A(\mult_22/ab[33][17] ), .B(
        \mult_22/CARRYB[32][17] ), .CI(\mult_22/SUMB[32][18] ), .CO(
        \mult_22/CARRYB[33][17] ), .S(\mult_22/SUMB[33][17] ) );
  FA_X1 \mult_22/S2_33_16  ( .A(\mult_22/ab[33][16] ), .B(
        \mult_22/CARRYB[32][16] ), .CI(\mult_22/SUMB[32][17] ), .CO(
        \mult_22/CARRYB[33][16] ), .S(\mult_22/SUMB[33][16] ) );
  FA_X1 \mult_22/S2_33_15  ( .A(\mult_22/ab[33][15] ), .B(
        \mult_22/CARRYB[32][15] ), .CI(\mult_22/SUMB[32][16] ), .CO(
        \mult_22/CARRYB[33][15] ), .S(\mult_22/SUMB[33][15] ) );
  FA_X1 \mult_22/S2_33_14  ( .A(\mult_22/ab[33][14] ), .B(
        \mult_22/CARRYB[32][14] ), .CI(\mult_22/SUMB[32][15] ), .CO(
        \mult_22/CARRYB[33][14] ), .S(\mult_22/SUMB[33][14] ) );
  FA_X1 \mult_22/S2_33_13  ( .A(\mult_22/ab[33][13] ), .B(
        \mult_22/CARRYB[32][13] ), .CI(\mult_22/SUMB[32][14] ), .CO(
        \mult_22/CARRYB[33][13] ), .S(\mult_22/SUMB[33][13] ) );
  FA_X1 \mult_22/S2_33_12  ( .A(\mult_22/ab[33][12] ), .B(
        \mult_22/CARRYB[32][12] ), .CI(\mult_22/SUMB[32][13] ), .CO(
        \mult_22/CARRYB[33][12] ), .S(\mult_22/SUMB[33][12] ) );
  FA_X1 \mult_22/S2_33_11  ( .A(\mult_22/ab[33][11] ), .B(
        \mult_22/CARRYB[32][11] ), .CI(\mult_22/SUMB[32][12] ), .CO(
        \mult_22/CARRYB[33][11] ), .S(\mult_22/SUMB[33][11] ) );
  FA_X1 \mult_22/S2_33_10  ( .A(\mult_22/ab[33][10] ), .B(
        \mult_22/CARRYB[32][10] ), .CI(\mult_22/SUMB[32][11] ), .CO(
        \mult_22/CARRYB[33][10] ), .S(\mult_22/SUMB[33][10] ) );
  FA_X1 \mult_22/S2_33_9  ( .A(\mult_22/ab[33][9] ), .B(
        \mult_22/CARRYB[32][9] ), .CI(\mult_22/SUMB[32][10] ), .CO(
        \mult_22/CARRYB[33][9] ), .S(\mult_22/SUMB[33][9] ) );
  FA_X1 \mult_22/S2_33_8  ( .A(\mult_22/ab[33][8] ), .B(
        \mult_22/CARRYB[32][8] ), .CI(\mult_22/SUMB[32][9] ), .CO(
        \mult_22/CARRYB[33][8] ), .S(\mult_22/SUMB[33][8] ) );
  FA_X1 \mult_22/S2_33_7  ( .A(\mult_22/ab[33][7] ), .B(
        \mult_22/CARRYB[32][7] ), .CI(\mult_22/SUMB[32][8] ), .CO(
        \mult_22/CARRYB[33][7] ), .S(\mult_22/SUMB[33][7] ) );
  FA_X1 \mult_22/S2_33_6  ( .A(\mult_22/ab[33][6] ), .B(
        \mult_22/CARRYB[32][6] ), .CI(\mult_22/SUMB[32][7] ), .CO(
        \mult_22/CARRYB[33][6] ), .S(\mult_22/SUMB[33][6] ) );
  FA_X1 \mult_22/S2_33_5  ( .A(\mult_22/ab[33][5] ), .B(
        \mult_22/CARRYB[32][5] ), .CI(\mult_22/SUMB[32][6] ), .CO(
        \mult_22/CARRYB[33][5] ), .S(\mult_22/SUMB[33][5] ) );
  FA_X1 \mult_22/S2_33_4  ( .A(\mult_22/ab[33][4] ), .B(
        \mult_22/CARRYB[32][4] ), .CI(\mult_22/SUMB[32][5] ), .CO(
        \mult_22/CARRYB[33][4] ), .S(\mult_22/SUMB[33][4] ) );
  FA_X1 \mult_22/S2_33_3  ( .A(\mult_22/ab[33][3] ), .B(
        \mult_22/CARRYB[32][3] ), .CI(\mult_22/SUMB[32][4] ), .CO(
        \mult_22/CARRYB[33][3] ), .S(\mult_22/SUMB[33][3] ) );
  FA_X1 \mult_22/S2_33_2  ( .A(\mult_22/ab[33][2] ), .B(
        \mult_22/CARRYB[32][2] ), .CI(\mult_22/SUMB[32][3] ), .CO(
        \mult_22/CARRYB[33][2] ), .S(\mult_22/SUMB[33][2] ) );
  FA_X1 \mult_22/S2_33_1  ( .A(\mult_22/ab[33][1] ), .B(
        \mult_22/CARRYB[32][1] ), .CI(\mult_22/SUMB[32][2] ), .CO(
        \mult_22/CARRYB[33][1] ), .S(\mult_22/SUMB[33][1] ) );
  FA_X1 \mult_22/S1_33_0  ( .A(\mult_22/ab[33][0] ), .B(
        \mult_22/CARRYB[32][0] ), .CI(\mult_22/SUMB[32][1] ), .CO(
        \mult_22/CARRYB[33][0] ), .S(N161) );
  FA_X1 \mult_22/S3_34_62  ( .A(\mult_22/ab[34][62] ), .B(
        \mult_22/CARRYB[33][62] ), .CI(\mult_22/ab[33][63] ), .CO(
        \mult_22/CARRYB[34][62] ), .S(\mult_22/SUMB[34][62] ) );
  FA_X1 \mult_22/S2_34_61  ( .A(\mult_22/ab[34][61] ), .B(
        \mult_22/CARRYB[33][61] ), .CI(\mult_22/SUMB[33][62] ), .CO(
        \mult_22/CARRYB[34][61] ), .S(\mult_22/SUMB[34][61] ) );
  FA_X1 \mult_22/S2_34_60  ( .A(\mult_22/ab[34][60] ), .B(
        \mult_22/CARRYB[33][60] ), .CI(\mult_22/SUMB[33][61] ), .CO(
        \mult_22/CARRYB[34][60] ), .S(\mult_22/SUMB[34][60] ) );
  FA_X1 \mult_22/S2_34_59  ( .A(\mult_22/ab[34][59] ), .B(
        \mult_22/CARRYB[33][59] ), .CI(\mult_22/SUMB[33][60] ), .CO(
        \mult_22/CARRYB[34][59] ), .S(\mult_22/SUMB[34][59] ) );
  FA_X1 \mult_22/S2_34_58  ( .A(\mult_22/ab[34][58] ), .B(
        \mult_22/CARRYB[33][58] ), .CI(\mult_22/SUMB[33][59] ), .CO(
        \mult_22/CARRYB[34][58] ), .S(\mult_22/SUMB[34][58] ) );
  FA_X1 \mult_22/S2_34_57  ( .A(\mult_22/ab[34][57] ), .B(
        \mult_22/CARRYB[33][57] ), .CI(\mult_22/SUMB[33][58] ), .CO(
        \mult_22/CARRYB[34][57] ), .S(\mult_22/SUMB[34][57] ) );
  FA_X1 \mult_22/S2_34_56  ( .A(\mult_22/ab[34][56] ), .B(
        \mult_22/CARRYB[33][56] ), .CI(\mult_22/SUMB[33][57] ), .CO(
        \mult_22/CARRYB[34][56] ), .S(\mult_22/SUMB[34][56] ) );
  FA_X1 \mult_22/S2_34_55  ( .A(\mult_22/ab[34][55] ), .B(
        \mult_22/CARRYB[33][55] ), .CI(\mult_22/SUMB[33][56] ), .CO(
        \mult_22/CARRYB[34][55] ), .S(\mult_22/SUMB[34][55] ) );
  FA_X1 \mult_22/S2_34_54  ( .A(\mult_22/ab[34][54] ), .B(
        \mult_22/CARRYB[33][54] ), .CI(\mult_22/SUMB[33][55] ), .CO(
        \mult_22/CARRYB[34][54] ), .S(\mult_22/SUMB[34][54] ) );
  FA_X1 \mult_22/S2_34_53  ( .A(\mult_22/ab[34][53] ), .B(
        \mult_22/CARRYB[33][53] ), .CI(\mult_22/SUMB[33][54] ), .CO(
        \mult_22/CARRYB[34][53] ), .S(\mult_22/SUMB[34][53] ) );
  FA_X1 \mult_22/S2_34_52  ( .A(\mult_22/ab[34][52] ), .B(
        \mult_22/CARRYB[33][52] ), .CI(\mult_22/SUMB[33][53] ), .CO(
        \mult_22/CARRYB[34][52] ), .S(\mult_22/SUMB[34][52] ) );
  FA_X1 \mult_22/S2_34_51  ( .A(\mult_22/ab[34][51] ), .B(
        \mult_22/CARRYB[33][51] ), .CI(\mult_22/SUMB[33][52] ), .CO(
        \mult_22/CARRYB[34][51] ), .S(\mult_22/SUMB[34][51] ) );
  FA_X1 \mult_22/S2_34_50  ( .A(\mult_22/ab[34][50] ), .B(
        \mult_22/CARRYB[33][50] ), .CI(\mult_22/SUMB[33][51] ), .CO(
        \mult_22/CARRYB[34][50] ), .S(\mult_22/SUMB[34][50] ) );
  FA_X1 \mult_22/S2_34_49  ( .A(\mult_22/ab[34][49] ), .B(
        \mult_22/CARRYB[33][49] ), .CI(\mult_22/SUMB[33][50] ), .CO(
        \mult_22/CARRYB[34][49] ), .S(\mult_22/SUMB[34][49] ) );
  FA_X1 \mult_22/S2_34_48  ( .A(\mult_22/ab[34][48] ), .B(
        \mult_22/CARRYB[33][48] ), .CI(\mult_22/SUMB[33][49] ), .CO(
        \mult_22/CARRYB[34][48] ), .S(\mult_22/SUMB[34][48] ) );
  FA_X1 \mult_22/S2_34_47  ( .A(\mult_22/ab[34][47] ), .B(
        \mult_22/CARRYB[33][47] ), .CI(\mult_22/SUMB[33][48] ), .CO(
        \mult_22/CARRYB[34][47] ), .S(\mult_22/SUMB[34][47] ) );
  FA_X1 \mult_22/S2_34_46  ( .A(\mult_22/ab[34][46] ), .B(
        \mult_22/CARRYB[33][46] ), .CI(\mult_22/SUMB[33][47] ), .CO(
        \mult_22/CARRYB[34][46] ), .S(\mult_22/SUMB[34][46] ) );
  FA_X1 \mult_22/S2_34_45  ( .A(\mult_22/ab[34][45] ), .B(
        \mult_22/CARRYB[33][45] ), .CI(\mult_22/SUMB[33][46] ), .CO(
        \mult_22/CARRYB[34][45] ), .S(\mult_22/SUMB[34][45] ) );
  FA_X1 \mult_22/S2_34_44  ( .A(\mult_22/ab[34][44] ), .B(
        \mult_22/CARRYB[33][44] ), .CI(\mult_22/SUMB[33][45] ), .CO(
        \mult_22/CARRYB[34][44] ), .S(\mult_22/SUMB[34][44] ) );
  FA_X1 \mult_22/S2_34_43  ( .A(\mult_22/ab[34][43] ), .B(
        \mult_22/CARRYB[33][43] ), .CI(\mult_22/SUMB[33][44] ), .CO(
        \mult_22/CARRYB[34][43] ), .S(\mult_22/SUMB[34][43] ) );
  FA_X1 \mult_22/S2_34_42  ( .A(\mult_22/ab[34][42] ), .B(
        \mult_22/CARRYB[33][42] ), .CI(\mult_22/SUMB[33][43] ), .CO(
        \mult_22/CARRYB[34][42] ), .S(\mult_22/SUMB[34][42] ) );
  FA_X1 \mult_22/S2_34_41  ( .A(\mult_22/ab[34][41] ), .B(
        \mult_22/CARRYB[33][41] ), .CI(\mult_22/SUMB[33][42] ), .CO(
        \mult_22/CARRYB[34][41] ), .S(\mult_22/SUMB[34][41] ) );
  FA_X1 \mult_22/S2_34_40  ( .A(\mult_22/ab[34][40] ), .B(
        \mult_22/CARRYB[33][40] ), .CI(\mult_22/SUMB[33][41] ), .CO(
        \mult_22/CARRYB[34][40] ), .S(\mult_22/SUMB[34][40] ) );
  FA_X1 \mult_22/S2_34_39  ( .A(\mult_22/ab[34][39] ), .B(
        \mult_22/CARRYB[33][39] ), .CI(\mult_22/SUMB[33][40] ), .CO(
        \mult_22/CARRYB[34][39] ), .S(\mult_22/SUMB[34][39] ) );
  FA_X1 \mult_22/S2_34_38  ( .A(\mult_22/ab[34][38] ), .B(
        \mult_22/CARRYB[33][38] ), .CI(\mult_22/SUMB[33][39] ), .CO(
        \mult_22/CARRYB[34][38] ), .S(\mult_22/SUMB[34][38] ) );
  FA_X1 \mult_22/S2_34_37  ( .A(\mult_22/ab[34][37] ), .B(
        \mult_22/CARRYB[33][37] ), .CI(\mult_22/SUMB[33][38] ), .CO(
        \mult_22/CARRYB[34][37] ), .S(\mult_22/SUMB[34][37] ) );
  FA_X1 \mult_22/S2_34_36  ( .A(\mult_22/ab[34][36] ), .B(
        \mult_22/CARRYB[33][36] ), .CI(\mult_22/SUMB[33][37] ), .CO(
        \mult_22/CARRYB[34][36] ), .S(\mult_22/SUMB[34][36] ) );
  FA_X1 \mult_22/S2_34_35  ( .A(\mult_22/ab[34][35] ), .B(
        \mult_22/CARRYB[33][35] ), .CI(\mult_22/SUMB[33][36] ), .CO(
        \mult_22/CARRYB[34][35] ), .S(\mult_22/SUMB[34][35] ) );
  FA_X1 \mult_22/S2_34_34  ( .A(\mult_22/ab[34][34] ), .B(
        \mult_22/CARRYB[33][34] ), .CI(\mult_22/SUMB[33][35] ), .CO(
        \mult_22/CARRYB[34][34] ), .S(\mult_22/SUMB[34][34] ) );
  FA_X1 \mult_22/S2_34_33  ( .A(\mult_22/ab[34][33] ), .B(
        \mult_22/CARRYB[33][33] ), .CI(\mult_22/SUMB[33][34] ), .CO(
        \mult_22/CARRYB[34][33] ), .S(\mult_22/SUMB[34][33] ) );
  FA_X1 \mult_22/S2_34_32  ( .A(\mult_22/CARRYB[33][32] ), .B(
        \mult_22/ab[34][32] ), .CI(\mult_22/SUMB[33][33] ), .CO(
        \mult_22/CARRYB[34][32] ), .S(\mult_22/SUMB[34][32] ) );
  FA_X1 \mult_22/S2_34_31  ( .A(\mult_22/ab[34][31] ), .B(
        \mult_22/CARRYB[33][31] ), .CI(\mult_22/SUMB[33][32] ), .CO(
        \mult_22/CARRYB[34][31] ), .S(\mult_22/SUMB[34][31] ) );
  FA_X1 \mult_22/S2_34_30  ( .A(\mult_22/ab[34][30] ), .B(
        \mult_22/CARRYB[33][30] ), .CI(\mult_22/SUMB[33][31] ), .CO(
        \mult_22/CARRYB[34][30] ), .S(\mult_22/SUMB[34][30] ) );
  FA_X1 \mult_22/S2_34_28  ( .A(\mult_22/ab[34][28] ), .B(
        \mult_22/CARRYB[33][28] ), .CI(\mult_22/SUMB[33][29] ), .CO(
        \mult_22/CARRYB[34][28] ), .S(\mult_22/SUMB[34][28] ) );
  FA_X1 \mult_22/S2_34_27  ( .A(\mult_22/ab[34][27] ), .B(
        \mult_22/CARRYB[33][27] ), .CI(\mult_22/SUMB[33][28] ), .CO(
        \mult_22/CARRYB[34][27] ), .S(\mult_22/SUMB[34][27] ) );
  FA_X1 \mult_22/S2_34_26  ( .A(\mult_22/ab[34][26] ), .B(
        \mult_22/CARRYB[33][26] ), .CI(\mult_22/SUMB[33][27] ), .CO(
        \mult_22/CARRYB[34][26] ), .S(\mult_22/SUMB[34][26] ) );
  FA_X1 \mult_22/S2_34_25  ( .A(\mult_22/ab[34][25] ), .B(
        \mult_22/CARRYB[33][25] ), .CI(\mult_22/SUMB[33][26] ), .CO(
        \mult_22/CARRYB[34][25] ), .S(\mult_22/SUMB[34][25] ) );
  FA_X1 \mult_22/S2_34_24  ( .A(\mult_22/ab[34][24] ), .B(
        \mult_22/CARRYB[33][24] ), .CI(\mult_22/SUMB[33][25] ), .CO(
        \mult_22/CARRYB[34][24] ), .S(\mult_22/SUMB[34][24] ) );
  FA_X1 \mult_22/S2_34_23  ( .A(\mult_22/ab[34][23] ), .B(
        \mult_22/CARRYB[33][23] ), .CI(\mult_22/SUMB[33][24] ), .CO(
        \mult_22/CARRYB[34][23] ), .S(\mult_22/SUMB[34][23] ) );
  FA_X1 \mult_22/S2_34_22  ( .A(\mult_22/ab[34][22] ), .B(
        \mult_22/CARRYB[33][22] ), .CI(\mult_22/SUMB[33][23] ), .CO(
        \mult_22/CARRYB[34][22] ), .S(\mult_22/SUMB[34][22] ) );
  FA_X1 \mult_22/S2_34_21  ( .A(\mult_22/ab[34][21] ), .B(
        \mult_22/CARRYB[33][21] ), .CI(\mult_22/SUMB[33][22] ), .CO(
        \mult_22/CARRYB[34][21] ), .S(\mult_22/SUMB[34][21] ) );
  FA_X1 \mult_22/S2_34_20  ( .A(\mult_22/ab[34][20] ), .B(
        \mult_22/CARRYB[33][20] ), .CI(\mult_22/SUMB[33][21] ), .CO(
        \mult_22/CARRYB[34][20] ), .S(\mult_22/SUMB[34][20] ) );
  FA_X1 \mult_22/S2_34_19  ( .A(\mult_22/ab[34][19] ), .B(
        \mult_22/CARRYB[33][19] ), .CI(\mult_22/SUMB[33][20] ), .CO(
        \mult_22/CARRYB[34][19] ), .S(\mult_22/SUMB[34][19] ) );
  FA_X1 \mult_22/S2_34_18  ( .A(\mult_22/ab[34][18] ), .B(
        \mult_22/CARRYB[33][18] ), .CI(\mult_22/SUMB[33][19] ), .CO(
        \mult_22/CARRYB[34][18] ), .S(\mult_22/SUMB[34][18] ) );
  FA_X1 \mult_22/S2_34_17  ( .A(\mult_22/ab[34][17] ), .B(
        \mult_22/CARRYB[33][17] ), .CI(\mult_22/SUMB[33][18] ), .CO(
        \mult_22/CARRYB[34][17] ), .S(\mult_22/SUMB[34][17] ) );
  FA_X1 \mult_22/S2_34_16  ( .A(\mult_22/ab[34][16] ), .B(
        \mult_22/CARRYB[33][16] ), .CI(\mult_22/SUMB[33][17] ), .CO(
        \mult_22/CARRYB[34][16] ), .S(\mult_22/SUMB[34][16] ) );
  FA_X1 \mult_22/S2_34_15  ( .A(\mult_22/ab[34][15] ), .B(
        \mult_22/CARRYB[33][15] ), .CI(\mult_22/SUMB[33][16] ), .CO(
        \mult_22/CARRYB[34][15] ), .S(\mult_22/SUMB[34][15] ) );
  FA_X1 \mult_22/S2_34_14  ( .A(\mult_22/ab[34][14] ), .B(
        \mult_22/CARRYB[33][14] ), .CI(\mult_22/SUMB[33][15] ), .CO(
        \mult_22/CARRYB[34][14] ), .S(\mult_22/SUMB[34][14] ) );
  FA_X1 \mult_22/S2_34_13  ( .A(\mult_22/ab[34][13] ), .B(
        \mult_22/CARRYB[33][13] ), .CI(\mult_22/SUMB[33][14] ), .CO(
        \mult_22/CARRYB[34][13] ), .S(\mult_22/SUMB[34][13] ) );
  FA_X1 \mult_22/S2_34_12  ( .A(\mult_22/ab[34][12] ), .B(
        \mult_22/CARRYB[33][12] ), .CI(\mult_22/SUMB[33][13] ), .CO(
        \mult_22/CARRYB[34][12] ), .S(\mult_22/SUMB[34][12] ) );
  FA_X1 \mult_22/S2_34_11  ( .A(\mult_22/ab[34][11] ), .B(
        \mult_22/CARRYB[33][11] ), .CI(\mult_22/SUMB[33][12] ), .CO(
        \mult_22/CARRYB[34][11] ), .S(\mult_22/SUMB[34][11] ) );
  FA_X1 \mult_22/S2_34_10  ( .A(\mult_22/ab[34][10] ), .B(
        \mult_22/CARRYB[33][10] ), .CI(\mult_22/SUMB[33][11] ), .CO(
        \mult_22/CARRYB[34][10] ), .S(\mult_22/SUMB[34][10] ) );
  FA_X1 \mult_22/S2_34_9  ( .A(\mult_22/ab[34][9] ), .B(
        \mult_22/CARRYB[33][9] ), .CI(\mult_22/SUMB[33][10] ), .CO(
        \mult_22/CARRYB[34][9] ), .S(\mult_22/SUMB[34][9] ) );
  FA_X1 \mult_22/S2_34_8  ( .A(\mult_22/ab[34][8] ), .B(
        \mult_22/CARRYB[33][8] ), .CI(\mult_22/SUMB[33][9] ), .CO(
        \mult_22/CARRYB[34][8] ), .S(\mult_22/SUMB[34][8] ) );
  FA_X1 \mult_22/S2_34_7  ( .A(\mult_22/ab[34][7] ), .B(
        \mult_22/CARRYB[33][7] ), .CI(\mult_22/SUMB[33][8] ), .CO(
        \mult_22/CARRYB[34][7] ), .S(\mult_22/SUMB[34][7] ) );
  FA_X1 \mult_22/S2_34_6  ( .A(\mult_22/ab[34][6] ), .B(
        \mult_22/CARRYB[33][6] ), .CI(\mult_22/SUMB[33][7] ), .CO(
        \mult_22/CARRYB[34][6] ), .S(\mult_22/SUMB[34][6] ) );
  FA_X1 \mult_22/S2_34_5  ( .A(\mult_22/ab[34][5] ), .B(
        \mult_22/CARRYB[33][5] ), .CI(\mult_22/SUMB[33][6] ), .CO(
        \mult_22/CARRYB[34][5] ), .S(\mult_22/SUMB[34][5] ) );
  FA_X1 \mult_22/S2_34_4  ( .A(\mult_22/ab[34][4] ), .B(
        \mult_22/CARRYB[33][4] ), .CI(\mult_22/SUMB[33][5] ), .CO(
        \mult_22/CARRYB[34][4] ), .S(\mult_22/SUMB[34][4] ) );
  FA_X1 \mult_22/S2_34_3  ( .A(\mult_22/ab[34][3] ), .B(
        \mult_22/CARRYB[33][3] ), .CI(\mult_22/SUMB[33][4] ), .CO(
        \mult_22/CARRYB[34][3] ), .S(\mult_22/SUMB[34][3] ) );
  FA_X1 \mult_22/S2_34_2  ( .A(\mult_22/ab[34][2] ), .B(
        \mult_22/CARRYB[33][2] ), .CI(\mult_22/SUMB[33][3] ), .CO(
        \mult_22/CARRYB[34][2] ), .S(\mult_22/SUMB[34][2] ) );
  FA_X1 \mult_22/S2_34_1  ( .A(\mult_22/ab[34][1] ), .B(
        \mult_22/CARRYB[33][1] ), .CI(\mult_22/SUMB[33][2] ), .CO(
        \mult_22/CARRYB[34][1] ), .S(\mult_22/SUMB[34][1] ) );
  FA_X1 \mult_22/S1_34_0  ( .A(\mult_22/ab[34][0] ), .B(
        \mult_22/CARRYB[33][0] ), .CI(\mult_22/SUMB[33][1] ), .CO(
        \mult_22/CARRYB[34][0] ), .S(N162) );
  FA_X1 \mult_22/S3_35_62  ( .A(\mult_22/ab[35][62] ), .B(
        \mult_22/CARRYB[34][62] ), .CI(\mult_22/ab[34][63] ), .CO(
        \mult_22/CARRYB[35][62] ), .S(\mult_22/SUMB[35][62] ) );
  FA_X1 \mult_22/S2_35_61  ( .A(\mult_22/ab[35][61] ), .B(
        \mult_22/CARRYB[34][61] ), .CI(\mult_22/SUMB[34][62] ), .CO(
        \mult_22/CARRYB[35][61] ), .S(\mult_22/SUMB[35][61] ) );
  FA_X1 \mult_22/S2_35_60  ( .A(\mult_22/ab[35][60] ), .B(
        \mult_22/CARRYB[34][60] ), .CI(\mult_22/SUMB[34][61] ), .CO(
        \mult_22/CARRYB[35][60] ), .S(\mult_22/SUMB[35][60] ) );
  FA_X1 \mult_22/S2_35_59  ( .A(\mult_22/ab[35][59] ), .B(
        \mult_22/CARRYB[34][59] ), .CI(\mult_22/SUMB[34][60] ), .CO(
        \mult_22/CARRYB[35][59] ), .S(\mult_22/SUMB[35][59] ) );
  FA_X1 \mult_22/S2_35_58  ( .A(\mult_22/ab[35][58] ), .B(
        \mult_22/CARRYB[34][58] ), .CI(\mult_22/SUMB[34][59] ), .CO(
        \mult_22/CARRYB[35][58] ), .S(\mult_22/SUMB[35][58] ) );
  FA_X1 \mult_22/S2_35_57  ( .A(\mult_22/ab[35][57] ), .B(
        \mult_22/CARRYB[34][57] ), .CI(\mult_22/SUMB[34][58] ), .CO(
        \mult_22/CARRYB[35][57] ), .S(\mult_22/SUMB[35][57] ) );
  FA_X1 \mult_22/S2_35_56  ( .A(\mult_22/ab[35][56] ), .B(
        \mult_22/CARRYB[34][56] ), .CI(\mult_22/SUMB[34][57] ), .CO(
        \mult_22/CARRYB[35][56] ), .S(\mult_22/SUMB[35][56] ) );
  FA_X1 \mult_22/S2_35_55  ( .A(\mult_22/ab[35][55] ), .B(
        \mult_22/CARRYB[34][55] ), .CI(\mult_22/SUMB[34][56] ), .CO(
        \mult_22/CARRYB[35][55] ), .S(\mult_22/SUMB[35][55] ) );
  FA_X1 \mult_22/S2_35_54  ( .A(\mult_22/ab[35][54] ), .B(
        \mult_22/CARRYB[34][54] ), .CI(\mult_22/SUMB[34][55] ), .CO(
        \mult_22/CARRYB[35][54] ), .S(\mult_22/SUMB[35][54] ) );
  FA_X1 \mult_22/S2_35_53  ( .A(\mult_22/ab[35][53] ), .B(
        \mult_22/CARRYB[34][53] ), .CI(\mult_22/SUMB[34][54] ), .CO(
        \mult_22/CARRYB[35][53] ), .S(\mult_22/SUMB[35][53] ) );
  FA_X1 \mult_22/S2_35_52  ( .A(\mult_22/ab[35][52] ), .B(
        \mult_22/CARRYB[34][52] ), .CI(\mult_22/SUMB[34][53] ), .CO(
        \mult_22/CARRYB[35][52] ), .S(\mult_22/SUMB[35][52] ) );
  FA_X1 \mult_22/S2_35_51  ( .A(\mult_22/ab[35][51] ), .B(
        \mult_22/CARRYB[34][51] ), .CI(\mult_22/SUMB[34][52] ), .CO(
        \mult_22/CARRYB[35][51] ), .S(\mult_22/SUMB[35][51] ) );
  FA_X1 \mult_22/S2_35_50  ( .A(\mult_22/ab[35][50] ), .B(
        \mult_22/CARRYB[34][50] ), .CI(\mult_22/SUMB[34][51] ), .CO(
        \mult_22/CARRYB[35][50] ), .S(\mult_22/SUMB[35][50] ) );
  FA_X1 \mult_22/S2_35_49  ( .A(\mult_22/ab[35][49] ), .B(
        \mult_22/CARRYB[34][49] ), .CI(\mult_22/SUMB[34][50] ), .CO(
        \mult_22/CARRYB[35][49] ), .S(\mult_22/SUMB[35][49] ) );
  FA_X1 \mult_22/S2_35_48  ( .A(\mult_22/ab[35][48] ), .B(
        \mult_22/CARRYB[34][48] ), .CI(\mult_22/SUMB[34][49] ), .CO(
        \mult_22/CARRYB[35][48] ), .S(\mult_22/SUMB[35][48] ) );
  FA_X1 \mult_22/S2_35_47  ( .A(\mult_22/ab[35][47] ), .B(
        \mult_22/CARRYB[34][47] ), .CI(\mult_22/SUMB[34][48] ), .CO(
        \mult_22/CARRYB[35][47] ), .S(\mult_22/SUMB[35][47] ) );
  FA_X1 \mult_22/S2_35_46  ( .A(\mult_22/ab[35][46] ), .B(
        \mult_22/CARRYB[34][46] ), .CI(\mult_22/SUMB[34][47] ), .CO(
        \mult_22/CARRYB[35][46] ), .S(\mult_22/SUMB[35][46] ) );
  FA_X1 \mult_22/S2_35_45  ( .A(\mult_22/ab[35][45] ), .B(
        \mult_22/CARRYB[34][45] ), .CI(\mult_22/SUMB[34][46] ), .CO(
        \mult_22/CARRYB[35][45] ), .S(\mult_22/SUMB[35][45] ) );
  FA_X1 \mult_22/S2_35_44  ( .A(\mult_22/ab[35][44] ), .B(
        \mult_22/CARRYB[34][44] ), .CI(\mult_22/SUMB[34][45] ), .CO(
        \mult_22/CARRYB[35][44] ), .S(\mult_22/SUMB[35][44] ) );
  FA_X1 \mult_22/S2_35_43  ( .A(\mult_22/ab[35][43] ), .B(
        \mult_22/CARRYB[34][43] ), .CI(\mult_22/SUMB[34][44] ), .CO(
        \mult_22/CARRYB[35][43] ), .S(\mult_22/SUMB[35][43] ) );
  FA_X1 \mult_22/S2_35_42  ( .A(\mult_22/ab[35][42] ), .B(
        \mult_22/CARRYB[34][42] ), .CI(\mult_22/SUMB[34][43] ), .CO(
        \mult_22/CARRYB[35][42] ), .S(\mult_22/SUMB[35][42] ) );
  FA_X1 \mult_22/S2_35_41  ( .A(\mult_22/ab[35][41] ), .B(
        \mult_22/CARRYB[34][41] ), .CI(\mult_22/SUMB[34][42] ), .CO(
        \mult_22/CARRYB[35][41] ), .S(\mult_22/SUMB[35][41] ) );
  FA_X1 \mult_22/S2_35_40  ( .A(\mult_22/ab[35][40] ), .B(
        \mult_22/CARRYB[34][40] ), .CI(\mult_22/SUMB[34][41] ), .CO(
        \mult_22/CARRYB[35][40] ), .S(\mult_22/SUMB[35][40] ) );
  FA_X1 \mult_22/S2_35_39  ( .A(\mult_22/ab[35][39] ), .B(
        \mult_22/CARRYB[34][39] ), .CI(\mult_22/SUMB[34][40] ), .CO(
        \mult_22/CARRYB[35][39] ), .S(\mult_22/SUMB[35][39] ) );
  FA_X1 \mult_22/S2_35_38  ( .A(\mult_22/ab[35][38] ), .B(
        \mult_22/CARRYB[34][38] ), .CI(\mult_22/SUMB[34][39] ), .CO(
        \mult_22/CARRYB[35][38] ), .S(\mult_22/SUMB[35][38] ) );
  FA_X1 \mult_22/S2_35_37  ( .A(\mult_22/ab[35][37] ), .B(
        \mult_22/CARRYB[34][37] ), .CI(\mult_22/SUMB[34][38] ), .CO(
        \mult_22/CARRYB[35][37] ), .S(\mult_22/SUMB[35][37] ) );
  FA_X1 \mult_22/S2_35_36  ( .A(\mult_22/ab[35][36] ), .B(
        \mult_22/CARRYB[34][36] ), .CI(\mult_22/SUMB[34][37] ), .CO(
        \mult_22/CARRYB[35][36] ), .S(\mult_22/SUMB[35][36] ) );
  FA_X1 \mult_22/S2_35_35  ( .A(\mult_22/ab[35][35] ), .B(
        \mult_22/CARRYB[34][35] ), .CI(\mult_22/SUMB[34][36] ), .CO(
        \mult_22/CARRYB[35][35] ), .S(\mult_22/SUMB[35][35] ) );
  FA_X1 \mult_22/S2_35_34  ( .A(\mult_22/ab[35][34] ), .B(
        \mult_22/CARRYB[34][34] ), .CI(\mult_22/SUMB[34][35] ), .CO(
        \mult_22/CARRYB[35][34] ), .S(\mult_22/SUMB[35][34] ) );
  FA_X1 \mult_22/S2_35_33  ( .A(\mult_22/ab[35][33] ), .B(
        \mult_22/CARRYB[34][33] ), .CI(\mult_22/SUMB[34][34] ), .CO(
        \mult_22/CARRYB[35][33] ), .S(\mult_22/SUMB[35][33] ) );
  FA_X1 \mult_22/S2_35_32  ( .A(\mult_22/ab[35][32] ), .B(
        \mult_22/CARRYB[34][32] ), .CI(\mult_22/SUMB[34][33] ), .CO(
        \mult_22/CARRYB[35][32] ), .S(\mult_22/SUMB[35][32] ) );
  FA_X1 \mult_22/S2_35_31  ( .A(\mult_22/ab[35][31] ), .B(
        \mult_22/CARRYB[34][31] ), .CI(\mult_22/SUMB[34][32] ), .CO(
        \mult_22/CARRYB[35][31] ), .S(\mult_22/SUMB[35][31] ) );
  FA_X1 \mult_22/S2_35_30  ( .A(\mult_22/ab[35][30] ), .B(
        \mult_22/CARRYB[34][30] ), .CI(\mult_22/SUMB[34][31] ), .CO(
        \mult_22/CARRYB[35][30] ), .S(\mult_22/SUMB[35][30] ) );
  FA_X1 \mult_22/S2_35_29  ( .A(\mult_22/ab[35][29] ), .B(
        \mult_22/CARRYB[34][29] ), .CI(\mult_22/SUMB[34][30] ), .CO(
        \mult_22/CARRYB[35][29] ), .S(\mult_22/SUMB[35][29] ) );
  FA_X1 \mult_22/S2_35_28  ( .A(\mult_22/ab[35][28] ), .B(
        \mult_22/CARRYB[34][28] ), .CI(\mult_22/SUMB[34][29] ), .CO(
        \mult_22/CARRYB[35][28] ), .S(\mult_22/SUMB[35][28] ) );
  FA_X1 \mult_22/S2_35_27  ( .A(\mult_22/ab[35][27] ), .B(
        \mult_22/CARRYB[34][27] ), .CI(\mult_22/SUMB[34][28] ), .CO(
        \mult_22/CARRYB[35][27] ), .S(\mult_22/SUMB[35][27] ) );
  FA_X1 \mult_22/S2_35_26  ( .A(\mult_22/ab[35][26] ), .B(
        \mult_22/CARRYB[34][26] ), .CI(\mult_22/SUMB[34][27] ), .CO(
        \mult_22/CARRYB[35][26] ), .S(\mult_22/SUMB[35][26] ) );
  FA_X1 \mult_22/S2_35_25  ( .A(\mult_22/ab[35][25] ), .B(
        \mult_22/CARRYB[34][25] ), .CI(\mult_22/SUMB[34][26] ), .CO(
        \mult_22/CARRYB[35][25] ), .S(\mult_22/SUMB[35][25] ) );
  FA_X1 \mult_22/S2_35_24  ( .A(\mult_22/ab[35][24] ), .B(
        \mult_22/CARRYB[34][24] ), .CI(\mult_22/SUMB[34][25] ), .CO(
        \mult_22/CARRYB[35][24] ), .S(\mult_22/SUMB[35][24] ) );
  FA_X1 \mult_22/S2_35_23  ( .A(\mult_22/ab[35][23] ), .B(
        \mult_22/CARRYB[34][23] ), .CI(\mult_22/SUMB[34][24] ), .CO(
        \mult_22/CARRYB[35][23] ), .S(\mult_22/SUMB[35][23] ) );
  FA_X1 \mult_22/S2_35_22  ( .A(\mult_22/ab[35][22] ), .B(
        \mult_22/CARRYB[34][22] ), .CI(\mult_22/SUMB[34][23] ), .CO(
        \mult_22/CARRYB[35][22] ), .S(\mult_22/SUMB[35][22] ) );
  FA_X1 \mult_22/S2_35_21  ( .A(\mult_22/ab[35][21] ), .B(
        \mult_22/CARRYB[34][21] ), .CI(\mult_22/SUMB[34][22] ), .CO(
        \mult_22/CARRYB[35][21] ), .S(\mult_22/SUMB[35][21] ) );
  FA_X1 \mult_22/S2_35_20  ( .A(\mult_22/ab[35][20] ), .B(
        \mult_22/CARRYB[34][20] ), .CI(\mult_22/SUMB[34][21] ), .CO(
        \mult_22/CARRYB[35][20] ), .S(\mult_22/SUMB[35][20] ) );
  FA_X1 \mult_22/S2_35_19  ( .A(\mult_22/ab[35][19] ), .B(
        \mult_22/CARRYB[34][19] ), .CI(\mult_22/SUMB[34][20] ), .CO(
        \mult_22/CARRYB[35][19] ), .S(\mult_22/SUMB[35][19] ) );
  FA_X1 \mult_22/S2_35_18  ( .A(\mult_22/ab[35][18] ), .B(
        \mult_22/CARRYB[34][18] ), .CI(\mult_22/SUMB[34][19] ), .CO(
        \mult_22/CARRYB[35][18] ), .S(\mult_22/SUMB[35][18] ) );
  FA_X1 \mult_22/S2_35_17  ( .A(\mult_22/ab[35][17] ), .B(
        \mult_22/CARRYB[34][17] ), .CI(\mult_22/SUMB[34][18] ), .CO(
        \mult_22/CARRYB[35][17] ), .S(\mult_22/SUMB[35][17] ) );
  FA_X1 \mult_22/S2_35_16  ( .A(\mult_22/ab[35][16] ), .B(
        \mult_22/CARRYB[34][16] ), .CI(\mult_22/SUMB[34][17] ), .CO(
        \mult_22/CARRYB[35][16] ), .S(\mult_22/SUMB[35][16] ) );
  FA_X1 \mult_22/S2_35_15  ( .A(\mult_22/ab[35][15] ), .B(
        \mult_22/CARRYB[34][15] ), .CI(\mult_22/SUMB[34][16] ), .CO(
        \mult_22/CARRYB[35][15] ), .S(\mult_22/SUMB[35][15] ) );
  FA_X1 \mult_22/S2_35_14  ( .A(\mult_22/ab[35][14] ), .B(
        \mult_22/CARRYB[34][14] ), .CI(\mult_22/SUMB[34][15] ), .CO(
        \mult_22/CARRYB[35][14] ), .S(\mult_22/SUMB[35][14] ) );
  FA_X1 \mult_22/S2_35_13  ( .A(\mult_22/ab[35][13] ), .B(
        \mult_22/CARRYB[34][13] ), .CI(\mult_22/SUMB[34][14] ), .CO(
        \mult_22/CARRYB[35][13] ), .S(\mult_22/SUMB[35][13] ) );
  FA_X1 \mult_22/S2_35_12  ( .A(\mult_22/ab[35][12] ), .B(
        \mult_22/CARRYB[34][12] ), .CI(\mult_22/SUMB[34][13] ), .CO(
        \mult_22/CARRYB[35][12] ), .S(\mult_22/SUMB[35][12] ) );
  FA_X1 \mult_22/S2_35_11  ( .A(\mult_22/ab[35][11] ), .B(
        \mult_22/CARRYB[34][11] ), .CI(\mult_22/SUMB[34][12] ), .CO(
        \mult_22/CARRYB[35][11] ), .S(\mult_22/SUMB[35][11] ) );
  FA_X1 \mult_22/S2_35_10  ( .A(\mult_22/ab[35][10] ), .B(
        \mult_22/CARRYB[34][10] ), .CI(\mult_22/SUMB[34][11] ), .CO(
        \mult_22/CARRYB[35][10] ), .S(\mult_22/SUMB[35][10] ) );
  FA_X1 \mult_22/S2_35_9  ( .A(\mult_22/ab[35][9] ), .B(
        \mult_22/CARRYB[34][9] ), .CI(\mult_22/SUMB[34][10] ), .CO(
        \mult_22/CARRYB[35][9] ), .S(\mult_22/SUMB[35][9] ) );
  FA_X1 \mult_22/S2_35_8  ( .A(\mult_22/ab[35][8] ), .B(
        \mult_22/CARRYB[34][8] ), .CI(\mult_22/SUMB[34][9] ), .CO(
        \mult_22/CARRYB[35][8] ), .S(\mult_22/SUMB[35][8] ) );
  FA_X1 \mult_22/S2_35_7  ( .A(\mult_22/ab[35][7] ), .B(
        \mult_22/CARRYB[34][7] ), .CI(\mult_22/SUMB[34][8] ), .CO(
        \mult_22/CARRYB[35][7] ), .S(\mult_22/SUMB[35][7] ) );
  FA_X1 \mult_22/S2_35_6  ( .A(\mult_22/ab[35][6] ), .B(
        \mult_22/CARRYB[34][6] ), .CI(\mult_22/SUMB[34][7] ), .CO(
        \mult_22/CARRYB[35][6] ), .S(\mult_22/SUMB[35][6] ) );
  FA_X1 \mult_22/S2_35_5  ( .A(\mult_22/ab[35][5] ), .B(
        \mult_22/CARRYB[34][5] ), .CI(\mult_22/SUMB[34][6] ), .CO(
        \mult_22/CARRYB[35][5] ), .S(\mult_22/SUMB[35][5] ) );
  FA_X1 \mult_22/S2_35_4  ( .A(\mult_22/ab[35][4] ), .B(
        \mult_22/CARRYB[34][4] ), .CI(\mult_22/SUMB[34][5] ), .CO(
        \mult_22/CARRYB[35][4] ), .S(\mult_22/SUMB[35][4] ) );
  FA_X1 \mult_22/S2_35_3  ( .A(\mult_22/ab[35][3] ), .B(
        \mult_22/CARRYB[34][3] ), .CI(\mult_22/SUMB[34][4] ), .CO(
        \mult_22/CARRYB[35][3] ), .S(\mult_22/SUMB[35][3] ) );
  FA_X1 \mult_22/S2_35_2  ( .A(\mult_22/ab[35][2] ), .B(
        \mult_22/CARRYB[34][2] ), .CI(\mult_22/SUMB[34][3] ), .CO(
        \mult_22/CARRYB[35][2] ), .S(\mult_22/SUMB[35][2] ) );
  FA_X1 \mult_22/S2_35_1  ( .A(\mult_22/ab[35][1] ), .B(
        \mult_22/CARRYB[34][1] ), .CI(\mult_22/SUMB[34][2] ), .CO(
        \mult_22/CARRYB[35][1] ), .S(\mult_22/SUMB[35][1] ) );
  FA_X1 \mult_22/S1_35_0  ( .A(\mult_22/ab[35][0] ), .B(
        \mult_22/CARRYB[34][0] ), .CI(\mult_22/SUMB[34][1] ), .CO(
        \mult_22/CARRYB[35][0] ), .S(N163) );
  FA_X1 \mult_22/S3_36_62  ( .A(\mult_22/ab[36][62] ), .B(
        \mult_22/CARRYB[35][62] ), .CI(\mult_22/ab[35][63] ), .CO(
        \mult_22/CARRYB[36][62] ), .S(\mult_22/SUMB[36][62] ) );
  FA_X1 \mult_22/S2_36_61  ( .A(\mult_22/ab[36][61] ), .B(
        \mult_22/CARRYB[35][61] ), .CI(\mult_22/SUMB[35][62] ), .CO(
        \mult_22/CARRYB[36][61] ), .S(\mult_22/SUMB[36][61] ) );
  FA_X1 \mult_22/S2_36_60  ( .A(\mult_22/ab[36][60] ), .B(
        \mult_22/CARRYB[35][60] ), .CI(\mult_22/SUMB[35][61] ), .CO(
        \mult_22/CARRYB[36][60] ), .S(\mult_22/SUMB[36][60] ) );
  FA_X1 \mult_22/S2_36_59  ( .A(\mult_22/ab[36][59] ), .B(
        \mult_22/CARRYB[35][59] ), .CI(\mult_22/SUMB[35][60] ), .CO(
        \mult_22/CARRYB[36][59] ), .S(\mult_22/SUMB[36][59] ) );
  FA_X1 \mult_22/S2_36_58  ( .A(\mult_22/ab[36][58] ), .B(
        \mult_22/CARRYB[35][58] ), .CI(\mult_22/SUMB[35][59] ), .CO(
        \mult_22/CARRYB[36][58] ), .S(\mult_22/SUMB[36][58] ) );
  FA_X1 \mult_22/S2_36_57  ( .A(\mult_22/ab[36][57] ), .B(
        \mult_22/CARRYB[35][57] ), .CI(\mult_22/SUMB[35][58] ), .CO(
        \mult_22/CARRYB[36][57] ), .S(\mult_22/SUMB[36][57] ) );
  FA_X1 \mult_22/S2_36_56  ( .A(\mult_22/ab[36][56] ), .B(
        \mult_22/CARRYB[35][56] ), .CI(\mult_22/SUMB[35][57] ), .CO(
        \mult_22/CARRYB[36][56] ), .S(\mult_22/SUMB[36][56] ) );
  FA_X1 \mult_22/S2_36_55  ( .A(\mult_22/ab[36][55] ), .B(
        \mult_22/CARRYB[35][55] ), .CI(\mult_22/SUMB[35][56] ), .CO(
        \mult_22/CARRYB[36][55] ), .S(\mult_22/SUMB[36][55] ) );
  FA_X1 \mult_22/S2_36_54  ( .A(\mult_22/ab[36][54] ), .B(
        \mult_22/CARRYB[35][54] ), .CI(\mult_22/SUMB[35][55] ), .CO(
        \mult_22/CARRYB[36][54] ), .S(\mult_22/SUMB[36][54] ) );
  FA_X1 \mult_22/S2_36_53  ( .A(\mult_22/ab[36][53] ), .B(
        \mult_22/CARRYB[35][53] ), .CI(\mult_22/SUMB[35][54] ), .CO(
        \mult_22/CARRYB[36][53] ), .S(\mult_22/SUMB[36][53] ) );
  FA_X1 \mult_22/S2_36_52  ( .A(\mult_22/ab[36][52] ), .B(
        \mult_22/CARRYB[35][52] ), .CI(\mult_22/SUMB[35][53] ), .CO(
        \mult_22/CARRYB[36][52] ), .S(\mult_22/SUMB[36][52] ) );
  FA_X1 \mult_22/S2_36_51  ( .A(\mult_22/ab[36][51] ), .B(
        \mult_22/CARRYB[35][51] ), .CI(\mult_22/SUMB[35][52] ), .CO(
        \mult_22/CARRYB[36][51] ), .S(\mult_22/SUMB[36][51] ) );
  FA_X1 \mult_22/S2_36_50  ( .A(\mult_22/ab[36][50] ), .B(
        \mult_22/CARRYB[35][50] ), .CI(\mult_22/SUMB[35][51] ), .CO(
        \mult_22/CARRYB[36][50] ), .S(\mult_22/SUMB[36][50] ) );
  FA_X1 \mult_22/S2_36_49  ( .A(\mult_22/ab[36][49] ), .B(
        \mult_22/CARRYB[35][49] ), .CI(\mult_22/SUMB[35][50] ), .CO(
        \mult_22/CARRYB[36][49] ), .S(\mult_22/SUMB[36][49] ) );
  FA_X1 \mult_22/S2_36_48  ( .A(\mult_22/ab[36][48] ), .B(
        \mult_22/CARRYB[35][48] ), .CI(\mult_22/SUMB[35][49] ), .CO(
        \mult_22/CARRYB[36][48] ), .S(\mult_22/SUMB[36][48] ) );
  FA_X1 \mult_22/S2_36_47  ( .A(\mult_22/ab[36][47] ), .B(
        \mult_22/CARRYB[35][47] ), .CI(\mult_22/SUMB[35][48] ), .CO(
        \mult_22/CARRYB[36][47] ), .S(\mult_22/SUMB[36][47] ) );
  FA_X1 \mult_22/S2_36_46  ( .A(\mult_22/ab[36][46] ), .B(
        \mult_22/CARRYB[35][46] ), .CI(\mult_22/SUMB[35][47] ), .CO(
        \mult_22/CARRYB[36][46] ), .S(\mult_22/SUMB[36][46] ) );
  FA_X1 \mult_22/S2_36_45  ( .A(\mult_22/ab[36][45] ), .B(
        \mult_22/CARRYB[35][45] ), .CI(\mult_22/SUMB[35][46] ), .CO(
        \mult_22/CARRYB[36][45] ), .S(\mult_22/SUMB[36][45] ) );
  FA_X1 \mult_22/S2_36_44  ( .A(\mult_22/ab[36][44] ), .B(
        \mult_22/CARRYB[35][44] ), .CI(\mult_22/SUMB[35][45] ), .CO(
        \mult_22/CARRYB[36][44] ), .S(\mult_22/SUMB[36][44] ) );
  FA_X1 \mult_22/S2_36_43  ( .A(\mult_22/ab[36][43] ), .B(
        \mult_22/CARRYB[35][43] ), .CI(\mult_22/SUMB[35][44] ), .CO(
        \mult_22/CARRYB[36][43] ), .S(\mult_22/SUMB[36][43] ) );
  FA_X1 \mult_22/S2_36_42  ( .A(\mult_22/ab[36][42] ), .B(
        \mult_22/CARRYB[35][42] ), .CI(\mult_22/SUMB[35][43] ), .CO(
        \mult_22/CARRYB[36][42] ), .S(\mult_22/SUMB[36][42] ) );
  FA_X1 \mult_22/S2_36_41  ( .A(\mult_22/ab[36][41] ), .B(
        \mult_22/CARRYB[35][41] ), .CI(\mult_22/SUMB[35][42] ), .CO(
        \mult_22/CARRYB[36][41] ), .S(\mult_22/SUMB[36][41] ) );
  FA_X1 \mult_22/S2_36_40  ( .A(\mult_22/ab[36][40] ), .B(
        \mult_22/CARRYB[35][40] ), .CI(\mult_22/SUMB[35][41] ), .CO(
        \mult_22/CARRYB[36][40] ), .S(\mult_22/SUMB[36][40] ) );
  FA_X1 \mult_22/S2_36_39  ( .A(\mult_22/ab[36][39] ), .B(
        \mult_22/CARRYB[35][39] ), .CI(\mult_22/SUMB[35][40] ), .CO(
        \mult_22/CARRYB[36][39] ), .S(\mult_22/SUMB[36][39] ) );
  FA_X1 \mult_22/S2_36_38  ( .A(\mult_22/ab[36][38] ), .B(
        \mult_22/CARRYB[35][38] ), .CI(\mult_22/SUMB[35][39] ), .CO(
        \mult_22/CARRYB[36][38] ), .S(\mult_22/SUMB[36][38] ) );
  FA_X1 \mult_22/S2_36_37  ( .A(\mult_22/ab[36][37] ), .B(
        \mult_22/CARRYB[35][37] ), .CI(\mult_22/SUMB[35][38] ), .CO(
        \mult_22/CARRYB[36][37] ), .S(\mult_22/SUMB[36][37] ) );
  FA_X1 \mult_22/S2_36_36  ( .A(\mult_22/ab[36][36] ), .B(
        \mult_22/CARRYB[35][36] ), .CI(\mult_22/SUMB[35][37] ), .CO(
        \mult_22/CARRYB[36][36] ), .S(\mult_22/SUMB[36][36] ) );
  FA_X1 \mult_22/S2_36_35  ( .A(\mult_22/ab[36][35] ), .B(
        \mult_22/CARRYB[35][35] ), .CI(\mult_22/SUMB[35][36] ), .CO(
        \mult_22/CARRYB[36][35] ), .S(\mult_22/SUMB[36][35] ) );
  FA_X1 \mult_22/S2_36_34  ( .A(\mult_22/ab[36][34] ), .B(
        \mult_22/CARRYB[35][34] ), .CI(\mult_22/SUMB[35][35] ), .CO(
        \mult_22/CARRYB[36][34] ), .S(\mult_22/SUMB[36][34] ) );
  FA_X1 \mult_22/S2_36_33  ( .A(\mult_22/ab[36][33] ), .B(
        \mult_22/CARRYB[35][33] ), .CI(\mult_22/SUMB[35][34] ), .CO(
        \mult_22/CARRYB[36][33] ), .S(\mult_22/SUMB[36][33] ) );
  FA_X1 \mult_22/S2_36_32  ( .A(\mult_22/ab[36][32] ), .B(
        \mult_22/CARRYB[35][32] ), .CI(\mult_22/SUMB[35][33] ), .CO(
        \mult_22/CARRYB[36][32] ), .S(\mult_22/SUMB[36][32] ) );
  FA_X1 \mult_22/S2_36_31  ( .A(\mult_22/ab[36][31] ), .B(
        \mult_22/CARRYB[35][31] ), .CI(\mult_22/SUMB[35][32] ), .CO(
        \mult_22/CARRYB[36][31] ), .S(\mult_22/SUMB[36][31] ) );
  FA_X1 \mult_22/S2_36_30  ( .A(\mult_22/CARRYB[35][30] ), .B(
        \mult_22/ab[36][30] ), .CI(\mult_22/SUMB[35][31] ), .CO(
        \mult_22/CARRYB[36][30] ), .S(\mult_22/SUMB[36][30] ) );
  FA_X1 \mult_22/S2_36_29  ( .A(\mult_22/ab[36][29] ), .B(
        \mult_22/CARRYB[35][29] ), .CI(\mult_22/SUMB[35][30] ), .CO(
        \mult_22/CARRYB[36][29] ), .S(\mult_22/SUMB[36][29] ) );
  FA_X1 \mult_22/S2_36_28  ( .A(\mult_22/ab[36][28] ), .B(
        \mult_22/CARRYB[35][28] ), .CI(\mult_22/SUMB[35][29] ), .CO(
        \mult_22/CARRYB[36][28] ), .S(\mult_22/SUMB[36][28] ) );
  FA_X1 \mult_22/S2_36_27  ( .A(\mult_22/ab[36][27] ), .B(
        \mult_22/CARRYB[35][27] ), .CI(\mult_22/SUMB[35][28] ), .CO(
        \mult_22/CARRYB[36][27] ), .S(\mult_22/SUMB[36][27] ) );
  FA_X1 \mult_22/S2_36_26  ( .A(\mult_22/ab[36][26] ), .B(
        \mult_22/CARRYB[35][26] ), .CI(\mult_22/SUMB[35][27] ), .CO(
        \mult_22/CARRYB[36][26] ), .S(\mult_22/SUMB[36][26] ) );
  FA_X1 \mult_22/S2_36_25  ( .A(\mult_22/ab[36][25] ), .B(
        \mult_22/CARRYB[35][25] ), .CI(\mult_22/SUMB[35][26] ), .CO(
        \mult_22/CARRYB[36][25] ), .S(\mult_22/SUMB[36][25] ) );
  FA_X1 \mult_22/S2_36_24  ( .A(\mult_22/ab[36][24] ), .B(
        \mult_22/CARRYB[35][24] ), .CI(\mult_22/SUMB[35][25] ), .CO(
        \mult_22/CARRYB[36][24] ), .S(\mult_22/SUMB[36][24] ) );
  FA_X1 \mult_22/S2_36_23  ( .A(\mult_22/ab[36][23] ), .B(
        \mult_22/CARRYB[35][23] ), .CI(\mult_22/SUMB[35][24] ), .CO(
        \mult_22/CARRYB[36][23] ), .S(\mult_22/SUMB[36][23] ) );
  FA_X1 \mult_22/S2_36_22  ( .A(\mult_22/ab[36][22] ), .B(
        \mult_22/CARRYB[35][22] ), .CI(\mult_22/SUMB[35][23] ), .CO(
        \mult_22/CARRYB[36][22] ), .S(\mult_22/SUMB[36][22] ) );
  FA_X1 \mult_22/S2_36_21  ( .A(\mult_22/ab[36][21] ), .B(
        \mult_22/CARRYB[35][21] ), .CI(\mult_22/SUMB[35][22] ), .CO(
        \mult_22/CARRYB[36][21] ), .S(\mult_22/SUMB[36][21] ) );
  FA_X1 \mult_22/S2_36_20  ( .A(\mult_22/ab[36][20] ), .B(
        \mult_22/CARRYB[35][20] ), .CI(\mult_22/SUMB[35][21] ), .CO(
        \mult_22/CARRYB[36][20] ), .S(\mult_22/SUMB[36][20] ) );
  FA_X1 \mult_22/S2_36_19  ( .A(\mult_22/ab[36][19] ), .B(
        \mult_22/CARRYB[35][19] ), .CI(\mult_22/SUMB[35][20] ), .CO(
        \mult_22/CARRYB[36][19] ), .S(\mult_22/SUMB[36][19] ) );
  FA_X1 \mult_22/S2_36_18  ( .A(\mult_22/ab[36][18] ), .B(
        \mult_22/CARRYB[35][18] ), .CI(\mult_22/SUMB[35][19] ), .CO(
        \mult_22/CARRYB[36][18] ), .S(\mult_22/SUMB[36][18] ) );
  FA_X1 \mult_22/S2_36_17  ( .A(\mult_22/ab[36][17] ), .B(
        \mult_22/CARRYB[35][17] ), .CI(\mult_22/SUMB[35][18] ), .CO(
        \mult_22/CARRYB[36][17] ), .S(\mult_22/SUMB[36][17] ) );
  FA_X1 \mult_22/S2_36_16  ( .A(\mult_22/ab[36][16] ), .B(
        \mult_22/CARRYB[35][16] ), .CI(\mult_22/SUMB[35][17] ), .CO(
        \mult_22/CARRYB[36][16] ), .S(\mult_22/SUMB[36][16] ) );
  FA_X1 \mult_22/S2_36_15  ( .A(\mult_22/ab[36][15] ), .B(
        \mult_22/CARRYB[35][15] ), .CI(\mult_22/SUMB[35][16] ), .CO(
        \mult_22/CARRYB[36][15] ), .S(\mult_22/SUMB[36][15] ) );
  FA_X1 \mult_22/S2_36_14  ( .A(\mult_22/ab[36][14] ), .B(
        \mult_22/CARRYB[35][14] ), .CI(\mult_22/SUMB[35][15] ), .CO(
        \mult_22/CARRYB[36][14] ), .S(\mult_22/SUMB[36][14] ) );
  FA_X1 \mult_22/S2_36_13  ( .A(\mult_22/ab[36][13] ), .B(
        \mult_22/CARRYB[35][13] ), .CI(\mult_22/SUMB[35][14] ), .CO(
        \mult_22/CARRYB[36][13] ), .S(\mult_22/SUMB[36][13] ) );
  FA_X1 \mult_22/S2_36_12  ( .A(\mult_22/ab[36][12] ), .B(
        \mult_22/CARRYB[35][12] ), .CI(\mult_22/SUMB[35][13] ), .CO(
        \mult_22/CARRYB[36][12] ), .S(\mult_22/SUMB[36][12] ) );
  FA_X1 \mult_22/S2_36_11  ( .A(\mult_22/ab[36][11] ), .B(
        \mult_22/CARRYB[35][11] ), .CI(\mult_22/SUMB[35][12] ), .CO(
        \mult_22/CARRYB[36][11] ), .S(\mult_22/SUMB[36][11] ) );
  FA_X1 \mult_22/S2_36_10  ( .A(\mult_22/ab[36][10] ), .B(
        \mult_22/CARRYB[35][10] ), .CI(\mult_22/SUMB[35][11] ), .CO(
        \mult_22/CARRYB[36][10] ), .S(\mult_22/SUMB[36][10] ) );
  FA_X1 \mult_22/S2_36_9  ( .A(\mult_22/ab[36][9] ), .B(
        \mult_22/CARRYB[35][9] ), .CI(\mult_22/SUMB[35][10] ), .CO(
        \mult_22/CARRYB[36][9] ), .S(\mult_22/SUMB[36][9] ) );
  FA_X1 \mult_22/S2_36_8  ( .A(\mult_22/ab[36][8] ), .B(
        \mult_22/CARRYB[35][8] ), .CI(\mult_22/SUMB[35][9] ), .CO(
        \mult_22/CARRYB[36][8] ), .S(\mult_22/SUMB[36][8] ) );
  FA_X1 \mult_22/S2_36_7  ( .A(\mult_22/ab[36][7] ), .B(
        \mult_22/CARRYB[35][7] ), .CI(\mult_22/SUMB[35][8] ), .CO(
        \mult_22/CARRYB[36][7] ), .S(\mult_22/SUMB[36][7] ) );
  FA_X1 \mult_22/S2_36_6  ( .A(\mult_22/ab[36][6] ), .B(
        \mult_22/CARRYB[35][6] ), .CI(\mult_22/SUMB[35][7] ), .CO(
        \mult_22/CARRYB[36][6] ), .S(\mult_22/SUMB[36][6] ) );
  FA_X1 \mult_22/S2_36_5  ( .A(\mult_22/ab[36][5] ), .B(
        \mult_22/CARRYB[35][5] ), .CI(\mult_22/SUMB[35][6] ), .CO(
        \mult_22/CARRYB[36][5] ), .S(\mult_22/SUMB[36][5] ) );
  FA_X1 \mult_22/S2_36_4  ( .A(\mult_22/ab[36][4] ), .B(
        \mult_22/CARRYB[35][4] ), .CI(\mult_22/SUMB[35][5] ), .CO(
        \mult_22/CARRYB[36][4] ), .S(\mult_22/SUMB[36][4] ) );
  FA_X1 \mult_22/S2_36_3  ( .A(\mult_22/ab[36][3] ), .B(
        \mult_22/CARRYB[35][3] ), .CI(\mult_22/SUMB[35][4] ), .CO(
        \mult_22/CARRYB[36][3] ), .S(\mult_22/SUMB[36][3] ) );
  FA_X1 \mult_22/S2_36_2  ( .A(\mult_22/ab[36][2] ), .B(
        \mult_22/CARRYB[35][2] ), .CI(\mult_22/SUMB[35][3] ), .CO(
        \mult_22/CARRYB[36][2] ), .S(\mult_22/SUMB[36][2] ) );
  FA_X1 \mult_22/S2_36_1  ( .A(\mult_22/ab[36][1] ), .B(
        \mult_22/CARRYB[35][1] ), .CI(\mult_22/SUMB[35][2] ), .CO(
        \mult_22/CARRYB[36][1] ), .S(\mult_22/SUMB[36][1] ) );
  FA_X1 \mult_22/S1_36_0  ( .A(\mult_22/ab[36][0] ), .B(
        \mult_22/CARRYB[35][0] ), .CI(\mult_22/SUMB[35][1] ), .CO(
        \mult_22/CARRYB[36][0] ), .S(N164) );
  FA_X1 \mult_22/S3_37_62  ( .A(\mult_22/ab[37][62] ), .B(
        \mult_22/CARRYB[36][62] ), .CI(\mult_22/ab[36][63] ), .CO(
        \mult_22/CARRYB[37][62] ), .S(\mult_22/SUMB[37][62] ) );
  FA_X1 \mult_22/S2_37_61  ( .A(\mult_22/ab[37][61] ), .B(
        \mult_22/CARRYB[36][61] ), .CI(\mult_22/SUMB[36][62] ), .CO(
        \mult_22/CARRYB[37][61] ), .S(\mult_22/SUMB[37][61] ) );
  FA_X1 \mult_22/S2_37_60  ( .A(\mult_22/ab[37][60] ), .B(
        \mult_22/CARRYB[36][60] ), .CI(\mult_22/SUMB[36][61] ), .CO(
        \mult_22/CARRYB[37][60] ), .S(\mult_22/SUMB[37][60] ) );
  FA_X1 \mult_22/S2_37_59  ( .A(\mult_22/ab[37][59] ), .B(
        \mult_22/CARRYB[36][59] ), .CI(\mult_22/SUMB[36][60] ), .CO(
        \mult_22/CARRYB[37][59] ), .S(\mult_22/SUMB[37][59] ) );
  FA_X1 \mult_22/S2_37_58  ( .A(\mult_22/ab[37][58] ), .B(
        \mult_22/CARRYB[36][58] ), .CI(\mult_22/SUMB[36][59] ), .CO(
        \mult_22/CARRYB[37][58] ), .S(\mult_22/SUMB[37][58] ) );
  FA_X1 \mult_22/S2_37_57  ( .A(\mult_22/ab[37][57] ), .B(
        \mult_22/CARRYB[36][57] ), .CI(\mult_22/SUMB[36][58] ), .CO(
        \mult_22/CARRYB[37][57] ), .S(\mult_22/SUMB[37][57] ) );
  FA_X1 \mult_22/S2_37_56  ( .A(\mult_22/ab[37][56] ), .B(
        \mult_22/CARRYB[36][56] ), .CI(\mult_22/SUMB[36][57] ), .CO(
        \mult_22/CARRYB[37][56] ), .S(\mult_22/SUMB[37][56] ) );
  FA_X1 \mult_22/S2_37_55  ( .A(\mult_22/ab[37][55] ), .B(
        \mult_22/CARRYB[36][55] ), .CI(\mult_22/SUMB[36][56] ), .CO(
        \mult_22/CARRYB[37][55] ), .S(\mult_22/SUMB[37][55] ) );
  FA_X1 \mult_22/S2_37_54  ( .A(\mult_22/ab[37][54] ), .B(
        \mult_22/CARRYB[36][54] ), .CI(\mult_22/SUMB[36][55] ), .CO(
        \mult_22/CARRYB[37][54] ), .S(\mult_22/SUMB[37][54] ) );
  FA_X1 \mult_22/S2_37_53  ( .A(\mult_22/ab[37][53] ), .B(
        \mult_22/CARRYB[36][53] ), .CI(\mult_22/SUMB[36][54] ), .CO(
        \mult_22/CARRYB[37][53] ), .S(\mult_22/SUMB[37][53] ) );
  FA_X1 \mult_22/S2_37_52  ( .A(\mult_22/ab[37][52] ), .B(
        \mult_22/CARRYB[36][52] ), .CI(\mult_22/SUMB[36][53] ), .CO(
        \mult_22/CARRYB[37][52] ), .S(\mult_22/SUMB[37][52] ) );
  FA_X1 \mult_22/S2_37_51  ( .A(\mult_22/ab[37][51] ), .B(
        \mult_22/CARRYB[36][51] ), .CI(\mult_22/SUMB[36][52] ), .CO(
        \mult_22/CARRYB[37][51] ), .S(\mult_22/SUMB[37][51] ) );
  FA_X1 \mult_22/S2_37_50  ( .A(\mult_22/ab[37][50] ), .B(
        \mult_22/CARRYB[36][50] ), .CI(\mult_22/SUMB[36][51] ), .CO(
        \mult_22/CARRYB[37][50] ), .S(\mult_22/SUMB[37][50] ) );
  FA_X1 \mult_22/S2_37_49  ( .A(\mult_22/ab[37][49] ), .B(
        \mult_22/CARRYB[36][49] ), .CI(\mult_22/SUMB[36][50] ), .CO(
        \mult_22/CARRYB[37][49] ), .S(\mult_22/SUMB[37][49] ) );
  FA_X1 \mult_22/S2_37_48  ( .A(\mult_22/ab[37][48] ), .B(
        \mult_22/CARRYB[36][48] ), .CI(\mult_22/SUMB[36][49] ), .CO(
        \mult_22/CARRYB[37][48] ), .S(\mult_22/SUMB[37][48] ) );
  FA_X1 \mult_22/S2_37_47  ( .A(\mult_22/ab[37][47] ), .B(
        \mult_22/CARRYB[36][47] ), .CI(\mult_22/SUMB[36][48] ), .CO(
        \mult_22/CARRYB[37][47] ), .S(\mult_22/SUMB[37][47] ) );
  FA_X1 \mult_22/S2_37_46  ( .A(\mult_22/ab[37][46] ), .B(
        \mult_22/CARRYB[36][46] ), .CI(\mult_22/SUMB[36][47] ), .CO(
        \mult_22/CARRYB[37][46] ), .S(\mult_22/SUMB[37][46] ) );
  FA_X1 \mult_22/S2_37_45  ( .A(\mult_22/ab[37][45] ), .B(
        \mult_22/CARRYB[36][45] ), .CI(\mult_22/SUMB[36][46] ), .CO(
        \mult_22/CARRYB[37][45] ), .S(\mult_22/SUMB[37][45] ) );
  FA_X1 \mult_22/S2_37_44  ( .A(\mult_22/ab[37][44] ), .B(
        \mult_22/CARRYB[36][44] ), .CI(\mult_22/SUMB[36][45] ), .CO(
        \mult_22/CARRYB[37][44] ), .S(\mult_22/SUMB[37][44] ) );
  FA_X1 \mult_22/S2_37_43  ( .A(\mult_22/ab[37][43] ), .B(
        \mult_22/CARRYB[36][43] ), .CI(\mult_22/SUMB[36][44] ), .CO(
        \mult_22/CARRYB[37][43] ), .S(\mult_22/SUMB[37][43] ) );
  FA_X1 \mult_22/S2_37_42  ( .A(\mult_22/ab[37][42] ), .B(
        \mult_22/CARRYB[36][42] ), .CI(\mult_22/SUMB[36][43] ), .CO(
        \mult_22/CARRYB[37][42] ), .S(\mult_22/SUMB[37][42] ) );
  FA_X1 \mult_22/S2_37_41  ( .A(\mult_22/ab[37][41] ), .B(
        \mult_22/CARRYB[36][41] ), .CI(\mult_22/SUMB[36][42] ), .CO(
        \mult_22/CARRYB[37][41] ), .S(\mult_22/SUMB[37][41] ) );
  FA_X1 \mult_22/S2_37_40  ( .A(\mult_22/ab[37][40] ), .B(
        \mult_22/CARRYB[36][40] ), .CI(\mult_22/SUMB[36][41] ), .CO(
        \mult_22/CARRYB[37][40] ), .S(\mult_22/SUMB[37][40] ) );
  FA_X1 \mult_22/S2_37_39  ( .A(\mult_22/ab[37][39] ), .B(
        \mult_22/CARRYB[36][39] ), .CI(\mult_22/SUMB[36][40] ), .CO(
        \mult_22/CARRYB[37][39] ), .S(\mult_22/SUMB[37][39] ) );
  FA_X1 \mult_22/S2_37_38  ( .A(\mult_22/ab[37][38] ), .B(
        \mult_22/CARRYB[36][38] ), .CI(\mult_22/SUMB[36][39] ), .CO(
        \mult_22/CARRYB[37][38] ), .S(\mult_22/SUMB[37][38] ) );
  FA_X1 \mult_22/S2_37_37  ( .A(\mult_22/ab[37][37] ), .B(
        \mult_22/CARRYB[36][37] ), .CI(\mult_22/SUMB[36][38] ), .CO(
        \mult_22/CARRYB[37][37] ), .S(\mult_22/SUMB[37][37] ) );
  FA_X1 \mult_22/S2_37_36  ( .A(\mult_22/ab[37][36] ), .B(
        \mult_22/CARRYB[36][36] ), .CI(\mult_22/SUMB[36][37] ), .CO(
        \mult_22/CARRYB[37][36] ), .S(\mult_22/SUMB[37][36] ) );
  FA_X1 \mult_22/S2_37_35  ( .A(\mult_22/ab[37][35] ), .B(
        \mult_22/CARRYB[36][35] ), .CI(\mult_22/SUMB[36][36] ), .CO(
        \mult_22/CARRYB[37][35] ), .S(\mult_22/SUMB[37][35] ) );
  FA_X1 \mult_22/S2_37_34  ( .A(\mult_22/ab[37][34] ), .B(
        \mult_22/CARRYB[36][34] ), .CI(\mult_22/SUMB[36][35] ), .CO(
        \mult_22/CARRYB[37][34] ), .S(\mult_22/SUMB[37][34] ) );
  FA_X1 \mult_22/S2_37_33  ( .A(\mult_22/ab[37][33] ), .B(
        \mult_22/CARRYB[36][33] ), .CI(\mult_22/SUMB[36][34] ), .CO(
        \mult_22/CARRYB[37][33] ), .S(\mult_22/SUMB[37][33] ) );
  FA_X1 \mult_22/S2_37_32  ( .A(\mult_22/ab[37][32] ), .B(
        \mult_22/CARRYB[36][32] ), .CI(\mult_22/SUMB[36][33] ), .CO(
        \mult_22/CARRYB[37][32] ), .S(\mult_22/SUMB[37][32] ) );
  FA_X1 \mult_22/S2_37_31  ( .A(\mult_22/ab[37][31] ), .B(
        \mult_22/CARRYB[36][31] ), .CI(\mult_22/SUMB[36][32] ), .CO(
        \mult_22/CARRYB[37][31] ), .S(\mult_22/SUMB[37][31] ) );
  FA_X1 \mult_22/S2_37_30  ( .A(\mult_22/ab[37][30] ), .B(
        \mult_22/CARRYB[36][30] ), .CI(\mult_22/SUMB[36][31] ), .CO(
        \mult_22/CARRYB[37][30] ), .S(\mult_22/SUMB[37][30] ) );
  FA_X1 \mult_22/S2_37_29  ( .A(\mult_22/ab[37][29] ), .B(
        \mult_22/CARRYB[36][29] ), .CI(\mult_22/SUMB[36][30] ), .CO(
        \mult_22/CARRYB[37][29] ), .S(\mult_22/SUMB[37][29] ) );
  FA_X1 \mult_22/S2_37_28  ( .A(\mult_22/ab[37][28] ), .B(
        \mult_22/CARRYB[36][28] ), .CI(\mult_22/SUMB[36][29] ), .CO(
        \mult_22/CARRYB[37][28] ), .S(\mult_22/SUMB[37][28] ) );
  FA_X1 \mult_22/S2_37_27  ( .A(\mult_22/CARRYB[36][27] ), .B(
        \mult_22/ab[37][27] ), .CI(\mult_22/SUMB[36][28] ), .CO(
        \mult_22/CARRYB[37][27] ), .S(\mult_22/SUMB[37][27] ) );
  FA_X1 \mult_22/S2_37_26  ( .A(\mult_22/ab[37][26] ), .B(
        \mult_22/CARRYB[36][26] ), .CI(\mult_22/SUMB[36][27] ), .CO(
        \mult_22/CARRYB[37][26] ), .S(\mult_22/SUMB[37][26] ) );
  FA_X1 \mult_22/S2_37_25  ( .A(\mult_22/ab[37][25] ), .B(
        \mult_22/CARRYB[36][25] ), .CI(\mult_22/SUMB[36][26] ), .CO(
        \mult_22/CARRYB[37][25] ), .S(\mult_22/SUMB[37][25] ) );
  FA_X1 \mult_22/S2_37_24  ( .A(\mult_22/ab[37][24] ), .B(
        \mult_22/CARRYB[36][24] ), .CI(\mult_22/SUMB[36][25] ), .CO(
        \mult_22/CARRYB[37][24] ), .S(\mult_22/SUMB[37][24] ) );
  FA_X1 \mult_22/S2_37_23  ( .A(\mult_22/ab[37][23] ), .B(
        \mult_22/CARRYB[36][23] ), .CI(\mult_22/SUMB[36][24] ), .CO(
        \mult_22/CARRYB[37][23] ), .S(\mult_22/SUMB[37][23] ) );
  FA_X1 \mult_22/S2_37_22  ( .A(\mult_22/ab[37][22] ), .B(
        \mult_22/CARRYB[36][22] ), .CI(\mult_22/SUMB[36][23] ), .CO(
        \mult_22/CARRYB[37][22] ), .S(\mult_22/SUMB[37][22] ) );
  FA_X1 \mult_22/S2_37_21  ( .A(\mult_22/ab[37][21] ), .B(
        \mult_22/CARRYB[36][21] ), .CI(\mult_22/SUMB[36][22] ), .CO(
        \mult_22/CARRYB[37][21] ), .S(\mult_22/SUMB[37][21] ) );
  FA_X1 \mult_22/S2_37_20  ( .A(\mult_22/ab[37][20] ), .B(
        \mult_22/CARRYB[36][20] ), .CI(\mult_22/SUMB[36][21] ), .CO(
        \mult_22/CARRYB[37][20] ), .S(\mult_22/SUMB[37][20] ) );
  FA_X1 \mult_22/S2_37_19  ( .A(\mult_22/ab[37][19] ), .B(
        \mult_22/CARRYB[36][19] ), .CI(\mult_22/SUMB[36][20] ), .CO(
        \mult_22/CARRYB[37][19] ), .S(\mult_22/SUMB[37][19] ) );
  FA_X1 \mult_22/S2_37_18  ( .A(\mult_22/ab[37][18] ), .B(
        \mult_22/CARRYB[36][18] ), .CI(\mult_22/SUMB[36][19] ), .CO(
        \mult_22/CARRYB[37][18] ), .S(\mult_22/SUMB[37][18] ) );
  FA_X1 \mult_22/S2_37_17  ( .A(\mult_22/ab[37][17] ), .B(
        \mult_22/CARRYB[36][17] ), .CI(\mult_22/SUMB[36][18] ), .CO(
        \mult_22/CARRYB[37][17] ), .S(\mult_22/SUMB[37][17] ) );
  FA_X1 \mult_22/S2_37_16  ( .A(\mult_22/ab[37][16] ), .B(
        \mult_22/CARRYB[36][16] ), .CI(\mult_22/SUMB[36][17] ), .CO(
        \mult_22/CARRYB[37][16] ), .S(\mult_22/SUMB[37][16] ) );
  FA_X1 \mult_22/S2_37_15  ( .A(\mult_22/ab[37][15] ), .B(
        \mult_22/CARRYB[36][15] ), .CI(\mult_22/SUMB[36][16] ), .CO(
        \mult_22/CARRYB[37][15] ), .S(\mult_22/SUMB[37][15] ) );
  FA_X1 \mult_22/S2_37_14  ( .A(\mult_22/ab[37][14] ), .B(
        \mult_22/CARRYB[36][14] ), .CI(\mult_22/SUMB[36][15] ), .CO(
        \mult_22/CARRYB[37][14] ), .S(\mult_22/SUMB[37][14] ) );
  FA_X1 \mult_22/S2_37_13  ( .A(\mult_22/ab[37][13] ), .B(
        \mult_22/CARRYB[36][13] ), .CI(\mult_22/SUMB[36][14] ), .CO(
        \mult_22/CARRYB[37][13] ), .S(\mult_22/SUMB[37][13] ) );
  FA_X1 \mult_22/S2_37_12  ( .A(\mult_22/ab[37][12] ), .B(
        \mult_22/CARRYB[36][12] ), .CI(\mult_22/SUMB[36][13] ), .CO(
        \mult_22/CARRYB[37][12] ), .S(\mult_22/SUMB[37][12] ) );
  FA_X1 \mult_22/S2_37_11  ( .A(\mult_22/ab[37][11] ), .B(
        \mult_22/CARRYB[36][11] ), .CI(\mult_22/SUMB[36][12] ), .CO(
        \mult_22/CARRYB[37][11] ), .S(\mult_22/SUMB[37][11] ) );
  FA_X1 \mult_22/S2_37_10  ( .A(\mult_22/ab[37][10] ), .B(
        \mult_22/CARRYB[36][10] ), .CI(\mult_22/SUMB[36][11] ), .CO(
        \mult_22/CARRYB[37][10] ), .S(\mult_22/SUMB[37][10] ) );
  FA_X1 \mult_22/S2_37_9  ( .A(\mult_22/ab[37][9] ), .B(
        \mult_22/CARRYB[36][9] ), .CI(\mult_22/SUMB[36][10] ), .CO(
        \mult_22/CARRYB[37][9] ), .S(\mult_22/SUMB[37][9] ) );
  FA_X1 \mult_22/S2_37_8  ( .A(\mult_22/ab[37][8] ), .B(
        \mult_22/CARRYB[36][8] ), .CI(\mult_22/SUMB[36][9] ), .CO(
        \mult_22/CARRYB[37][8] ), .S(\mult_22/SUMB[37][8] ) );
  FA_X1 \mult_22/S2_37_7  ( .A(\mult_22/ab[37][7] ), .B(
        \mult_22/CARRYB[36][7] ), .CI(\mult_22/SUMB[36][8] ), .CO(
        \mult_22/CARRYB[37][7] ), .S(\mult_22/SUMB[37][7] ) );
  FA_X1 \mult_22/S2_37_6  ( .A(\mult_22/ab[37][6] ), .B(
        \mult_22/CARRYB[36][6] ), .CI(\mult_22/SUMB[36][7] ), .CO(
        \mult_22/CARRYB[37][6] ), .S(\mult_22/SUMB[37][6] ) );
  FA_X1 \mult_22/S2_37_5  ( .A(\mult_22/ab[37][5] ), .B(
        \mult_22/CARRYB[36][5] ), .CI(\mult_22/SUMB[36][6] ), .CO(
        \mult_22/CARRYB[37][5] ), .S(\mult_22/SUMB[37][5] ) );
  FA_X1 \mult_22/S2_37_4  ( .A(\mult_22/ab[37][4] ), .B(
        \mult_22/CARRYB[36][4] ), .CI(\mult_22/SUMB[36][5] ), .CO(
        \mult_22/CARRYB[37][4] ), .S(\mult_22/SUMB[37][4] ) );
  FA_X1 \mult_22/S2_37_3  ( .A(\mult_22/ab[37][3] ), .B(
        \mult_22/CARRYB[36][3] ), .CI(\mult_22/SUMB[36][4] ), .CO(
        \mult_22/CARRYB[37][3] ), .S(\mult_22/SUMB[37][3] ) );
  FA_X1 \mult_22/S2_37_2  ( .A(\mult_22/ab[37][2] ), .B(
        \mult_22/CARRYB[36][2] ), .CI(\mult_22/SUMB[36][3] ), .CO(
        \mult_22/CARRYB[37][2] ), .S(\mult_22/SUMB[37][2] ) );
  FA_X1 \mult_22/S2_37_1  ( .A(\mult_22/ab[37][1] ), .B(
        \mult_22/CARRYB[36][1] ), .CI(\mult_22/SUMB[36][2] ), .CO(
        \mult_22/CARRYB[37][1] ), .S(\mult_22/SUMB[37][1] ) );
  FA_X1 \mult_22/S1_37_0  ( .A(\mult_22/ab[37][0] ), .B(
        \mult_22/CARRYB[36][0] ), .CI(\mult_22/SUMB[36][1] ), .CO(
        \mult_22/CARRYB[37][0] ), .S(N165) );
  FA_X1 \mult_22/S3_38_62  ( .A(\mult_22/ab[38][62] ), .B(
        \mult_22/CARRYB[37][62] ), .CI(\mult_22/ab[37][63] ), .CO(
        \mult_22/CARRYB[38][62] ), .S(\mult_22/SUMB[38][62] ) );
  FA_X1 \mult_22/S2_38_61  ( .A(\mult_22/ab[38][61] ), .B(
        \mult_22/CARRYB[37][61] ), .CI(\mult_22/SUMB[37][62] ), .CO(
        \mult_22/CARRYB[38][61] ), .S(\mult_22/SUMB[38][61] ) );
  FA_X1 \mult_22/S2_38_60  ( .A(\mult_22/ab[38][60] ), .B(
        \mult_22/CARRYB[37][60] ), .CI(\mult_22/SUMB[37][61] ), .CO(
        \mult_22/CARRYB[38][60] ), .S(\mult_22/SUMB[38][60] ) );
  FA_X1 \mult_22/S2_38_59  ( .A(\mult_22/ab[38][59] ), .B(
        \mult_22/CARRYB[37][59] ), .CI(\mult_22/SUMB[37][60] ), .CO(
        \mult_22/CARRYB[38][59] ), .S(\mult_22/SUMB[38][59] ) );
  FA_X1 \mult_22/S2_38_58  ( .A(\mult_22/ab[38][58] ), .B(
        \mult_22/CARRYB[37][58] ), .CI(\mult_22/SUMB[37][59] ), .CO(
        \mult_22/CARRYB[38][58] ), .S(\mult_22/SUMB[38][58] ) );
  FA_X1 \mult_22/S2_38_57  ( .A(\mult_22/ab[38][57] ), .B(
        \mult_22/CARRYB[37][57] ), .CI(\mult_22/SUMB[37][58] ), .CO(
        \mult_22/CARRYB[38][57] ), .S(\mult_22/SUMB[38][57] ) );
  FA_X1 \mult_22/S2_38_56  ( .A(\mult_22/ab[38][56] ), .B(
        \mult_22/CARRYB[37][56] ), .CI(\mult_22/SUMB[37][57] ), .CO(
        \mult_22/CARRYB[38][56] ), .S(\mult_22/SUMB[38][56] ) );
  FA_X1 \mult_22/S2_38_55  ( .A(\mult_22/ab[38][55] ), .B(
        \mult_22/CARRYB[37][55] ), .CI(\mult_22/SUMB[37][56] ), .CO(
        \mult_22/CARRYB[38][55] ), .S(\mult_22/SUMB[38][55] ) );
  FA_X1 \mult_22/S2_38_54  ( .A(\mult_22/ab[38][54] ), .B(
        \mult_22/CARRYB[37][54] ), .CI(\mult_22/SUMB[37][55] ), .CO(
        \mult_22/CARRYB[38][54] ), .S(\mult_22/SUMB[38][54] ) );
  FA_X1 \mult_22/S2_38_53  ( .A(\mult_22/ab[38][53] ), .B(
        \mult_22/CARRYB[37][53] ), .CI(\mult_22/SUMB[37][54] ), .CO(
        \mult_22/CARRYB[38][53] ), .S(\mult_22/SUMB[38][53] ) );
  FA_X1 \mult_22/S2_38_52  ( .A(\mult_22/ab[38][52] ), .B(
        \mult_22/CARRYB[37][52] ), .CI(\mult_22/SUMB[37][53] ), .CO(
        \mult_22/CARRYB[38][52] ), .S(\mult_22/SUMB[38][52] ) );
  FA_X1 \mult_22/S2_38_51  ( .A(\mult_22/ab[38][51] ), .B(
        \mult_22/CARRYB[37][51] ), .CI(\mult_22/SUMB[37][52] ), .CO(
        \mult_22/CARRYB[38][51] ), .S(\mult_22/SUMB[38][51] ) );
  FA_X1 \mult_22/S2_38_50  ( .A(\mult_22/ab[38][50] ), .B(
        \mult_22/CARRYB[37][50] ), .CI(\mult_22/SUMB[37][51] ), .CO(
        \mult_22/CARRYB[38][50] ), .S(\mult_22/SUMB[38][50] ) );
  FA_X1 \mult_22/S2_38_49  ( .A(\mult_22/ab[38][49] ), .B(
        \mult_22/CARRYB[37][49] ), .CI(\mult_22/SUMB[37][50] ), .CO(
        \mult_22/CARRYB[38][49] ), .S(\mult_22/SUMB[38][49] ) );
  FA_X1 \mult_22/S2_38_48  ( .A(\mult_22/ab[38][48] ), .B(
        \mult_22/CARRYB[37][48] ), .CI(\mult_22/SUMB[37][49] ), .CO(
        \mult_22/CARRYB[38][48] ), .S(\mult_22/SUMB[38][48] ) );
  FA_X1 \mult_22/S2_38_47  ( .A(\mult_22/ab[38][47] ), .B(
        \mult_22/CARRYB[37][47] ), .CI(\mult_22/SUMB[37][48] ), .CO(
        \mult_22/CARRYB[38][47] ), .S(\mult_22/SUMB[38][47] ) );
  FA_X1 \mult_22/S2_38_46  ( .A(\mult_22/ab[38][46] ), .B(
        \mult_22/CARRYB[37][46] ), .CI(\mult_22/SUMB[37][47] ), .CO(
        \mult_22/CARRYB[38][46] ), .S(\mult_22/SUMB[38][46] ) );
  FA_X1 \mult_22/S2_38_45  ( .A(\mult_22/ab[38][45] ), .B(
        \mult_22/CARRYB[37][45] ), .CI(\mult_22/SUMB[37][46] ), .CO(
        \mult_22/CARRYB[38][45] ), .S(\mult_22/SUMB[38][45] ) );
  FA_X1 \mult_22/S2_38_44  ( .A(\mult_22/ab[38][44] ), .B(
        \mult_22/CARRYB[37][44] ), .CI(\mult_22/SUMB[37][45] ), .CO(
        \mult_22/CARRYB[38][44] ), .S(\mult_22/SUMB[38][44] ) );
  FA_X1 \mult_22/S2_38_43  ( .A(\mult_22/ab[38][43] ), .B(
        \mult_22/CARRYB[37][43] ), .CI(\mult_22/SUMB[37][44] ), .CO(
        \mult_22/CARRYB[38][43] ), .S(\mult_22/SUMB[38][43] ) );
  FA_X1 \mult_22/S2_38_42  ( .A(\mult_22/ab[38][42] ), .B(
        \mult_22/CARRYB[37][42] ), .CI(\mult_22/SUMB[37][43] ), .CO(
        \mult_22/CARRYB[38][42] ), .S(\mult_22/SUMB[38][42] ) );
  FA_X1 \mult_22/S2_38_41  ( .A(\mult_22/ab[38][41] ), .B(
        \mult_22/CARRYB[37][41] ), .CI(\mult_22/SUMB[37][42] ), .CO(
        \mult_22/CARRYB[38][41] ), .S(\mult_22/SUMB[38][41] ) );
  FA_X1 \mult_22/S2_38_40  ( .A(\mult_22/ab[38][40] ), .B(
        \mult_22/CARRYB[37][40] ), .CI(\mult_22/SUMB[37][41] ), .CO(
        \mult_22/CARRYB[38][40] ), .S(\mult_22/SUMB[38][40] ) );
  FA_X1 \mult_22/S2_38_39  ( .A(\mult_22/ab[38][39] ), .B(
        \mult_22/CARRYB[37][39] ), .CI(\mult_22/SUMB[37][40] ), .CO(
        \mult_22/CARRYB[38][39] ), .S(\mult_22/SUMB[38][39] ) );
  FA_X1 \mult_22/S2_38_38  ( .A(\mult_22/ab[38][38] ), .B(
        \mult_22/CARRYB[37][38] ), .CI(\mult_22/SUMB[37][39] ), .CO(
        \mult_22/CARRYB[38][38] ), .S(\mult_22/SUMB[38][38] ) );
  FA_X1 \mult_22/S2_38_37  ( .A(\mult_22/ab[38][37] ), .B(
        \mult_22/CARRYB[37][37] ), .CI(\mult_22/SUMB[37][38] ), .CO(
        \mult_22/CARRYB[38][37] ), .S(\mult_22/SUMB[38][37] ) );
  FA_X1 \mult_22/S2_38_36  ( .A(\mult_22/ab[38][36] ), .B(
        \mult_22/CARRYB[37][36] ), .CI(\mult_22/SUMB[37][37] ), .CO(
        \mult_22/CARRYB[38][36] ), .S(\mult_22/SUMB[38][36] ) );
  FA_X1 \mult_22/S2_38_35  ( .A(\mult_22/ab[38][35] ), .B(
        \mult_22/CARRYB[37][35] ), .CI(\mult_22/SUMB[37][36] ), .CO(
        \mult_22/CARRYB[38][35] ), .S(\mult_22/SUMB[38][35] ) );
  FA_X1 \mult_22/S2_38_34  ( .A(\mult_22/ab[38][34] ), .B(
        \mult_22/CARRYB[37][34] ), .CI(\mult_22/SUMB[37][35] ), .CO(
        \mult_22/CARRYB[38][34] ), .S(\mult_22/SUMB[38][34] ) );
  FA_X1 \mult_22/S2_38_33  ( .A(\mult_22/ab[38][33] ), .B(
        \mult_22/CARRYB[37][33] ), .CI(\mult_22/SUMB[37][34] ), .CO(
        \mult_22/CARRYB[38][33] ), .S(\mult_22/SUMB[38][33] ) );
  FA_X1 \mult_22/S2_38_32  ( .A(\mult_22/ab[38][32] ), .B(
        \mult_22/CARRYB[37][32] ), .CI(\mult_22/SUMB[37][33] ), .CO(
        \mult_22/CARRYB[38][32] ), .S(\mult_22/SUMB[38][32] ) );
  FA_X1 \mult_22/S2_38_31  ( .A(\mult_22/ab[38][31] ), .B(
        \mult_22/CARRYB[37][31] ), .CI(\mult_22/SUMB[37][32] ), .CO(
        \mult_22/CARRYB[38][31] ), .S(\mult_22/SUMB[38][31] ) );
  FA_X1 \mult_22/S2_38_30  ( .A(\mult_22/ab[38][30] ), .B(
        \mult_22/CARRYB[37][30] ), .CI(\mult_22/SUMB[37][31] ), .CO(
        \mult_22/CARRYB[38][30] ), .S(\mult_22/SUMB[38][30] ) );
  FA_X1 \mult_22/S2_38_29  ( .A(\mult_22/ab[38][29] ), .B(
        \mult_22/CARRYB[37][29] ), .CI(\mult_22/SUMB[37][30] ), .CO(
        \mult_22/CARRYB[38][29] ), .S(\mult_22/SUMB[38][29] ) );
  FA_X1 \mult_22/S2_38_28  ( .A(\mult_22/CARRYB[37][28] ), .B(
        \mult_22/ab[38][28] ), .CI(\mult_22/SUMB[37][29] ), .CO(
        \mult_22/CARRYB[38][28] ), .S(\mult_22/SUMB[38][28] ) );
  FA_X1 \mult_22/S2_38_27  ( .A(\mult_22/ab[38][27] ), .B(
        \mult_22/CARRYB[37][27] ), .CI(\mult_22/SUMB[37][28] ), .CO(
        \mult_22/CARRYB[38][27] ), .S(\mult_22/SUMB[38][27] ) );
  FA_X1 \mult_22/S2_38_26  ( .A(\mult_22/ab[38][26] ), .B(
        \mult_22/CARRYB[37][26] ), .CI(\mult_22/SUMB[37][27] ), .CO(
        \mult_22/CARRYB[38][26] ), .S(\mult_22/SUMB[38][26] ) );
  FA_X1 \mult_22/S2_38_25  ( .A(\mult_22/ab[38][25] ), .B(
        \mult_22/CARRYB[37][25] ), .CI(\mult_22/SUMB[37][26] ), .CO(
        \mult_22/CARRYB[38][25] ), .S(\mult_22/SUMB[38][25] ) );
  FA_X1 \mult_22/S2_38_24  ( .A(\mult_22/ab[38][24] ), .B(
        \mult_22/CARRYB[37][24] ), .CI(\mult_22/SUMB[37][25] ), .CO(
        \mult_22/CARRYB[38][24] ), .S(\mult_22/SUMB[38][24] ) );
  FA_X1 \mult_22/S2_38_23  ( .A(\mult_22/ab[38][23] ), .B(
        \mult_22/CARRYB[37][23] ), .CI(\mult_22/SUMB[37][24] ), .CO(
        \mult_22/CARRYB[38][23] ), .S(\mult_22/SUMB[38][23] ) );
  FA_X1 \mult_22/S2_38_22  ( .A(\mult_22/ab[38][22] ), .B(
        \mult_22/CARRYB[37][22] ), .CI(\mult_22/SUMB[37][23] ), .CO(
        \mult_22/CARRYB[38][22] ), .S(\mult_22/SUMB[38][22] ) );
  FA_X1 \mult_22/S2_38_21  ( .A(\mult_22/ab[38][21] ), .B(
        \mult_22/CARRYB[37][21] ), .CI(\mult_22/SUMB[37][22] ), .CO(
        \mult_22/CARRYB[38][21] ), .S(\mult_22/SUMB[38][21] ) );
  FA_X1 \mult_22/S2_38_20  ( .A(\mult_22/ab[38][20] ), .B(
        \mult_22/CARRYB[37][20] ), .CI(\mult_22/SUMB[37][21] ), .CO(
        \mult_22/CARRYB[38][20] ), .S(\mult_22/SUMB[38][20] ) );
  FA_X1 \mult_22/S2_38_19  ( .A(\mult_22/ab[38][19] ), .B(
        \mult_22/CARRYB[37][19] ), .CI(\mult_22/SUMB[37][20] ), .CO(
        \mult_22/CARRYB[38][19] ), .S(\mult_22/SUMB[38][19] ) );
  FA_X1 \mult_22/S2_38_18  ( .A(\mult_22/ab[38][18] ), .B(
        \mult_22/CARRYB[37][18] ), .CI(\mult_22/SUMB[37][19] ), .CO(
        \mult_22/CARRYB[38][18] ), .S(\mult_22/SUMB[38][18] ) );
  FA_X1 \mult_22/S2_38_17  ( .A(\mult_22/ab[38][17] ), .B(
        \mult_22/CARRYB[37][17] ), .CI(\mult_22/SUMB[37][18] ), .CO(
        \mult_22/CARRYB[38][17] ), .S(\mult_22/SUMB[38][17] ) );
  FA_X1 \mult_22/S2_38_16  ( .A(\mult_22/ab[38][16] ), .B(
        \mult_22/CARRYB[37][16] ), .CI(\mult_22/SUMB[37][17] ), .CO(
        \mult_22/CARRYB[38][16] ), .S(\mult_22/SUMB[38][16] ) );
  FA_X1 \mult_22/S2_38_15  ( .A(\mult_22/ab[38][15] ), .B(
        \mult_22/CARRYB[37][15] ), .CI(\mult_22/SUMB[37][16] ), .CO(
        \mult_22/CARRYB[38][15] ), .S(\mult_22/SUMB[38][15] ) );
  FA_X1 \mult_22/S2_38_14  ( .A(\mult_22/ab[38][14] ), .B(
        \mult_22/CARRYB[37][14] ), .CI(\mult_22/SUMB[37][15] ), .CO(
        \mult_22/CARRYB[38][14] ), .S(\mult_22/SUMB[38][14] ) );
  FA_X1 \mult_22/S2_38_13  ( .A(\mult_22/ab[38][13] ), .B(
        \mult_22/CARRYB[37][13] ), .CI(\mult_22/SUMB[37][14] ), .CO(
        \mult_22/CARRYB[38][13] ), .S(\mult_22/SUMB[38][13] ) );
  FA_X1 \mult_22/S2_38_12  ( .A(\mult_22/ab[38][12] ), .B(
        \mult_22/CARRYB[37][12] ), .CI(\mult_22/SUMB[37][13] ), .CO(
        \mult_22/CARRYB[38][12] ), .S(\mult_22/SUMB[38][12] ) );
  FA_X1 \mult_22/S2_38_11  ( .A(\mult_22/ab[38][11] ), .B(
        \mult_22/CARRYB[37][11] ), .CI(\mult_22/SUMB[37][12] ), .CO(
        \mult_22/CARRYB[38][11] ), .S(\mult_22/SUMB[38][11] ) );
  FA_X1 \mult_22/S2_38_10  ( .A(\mult_22/ab[38][10] ), .B(
        \mult_22/CARRYB[37][10] ), .CI(\mult_22/SUMB[37][11] ), .CO(
        \mult_22/CARRYB[38][10] ), .S(\mult_22/SUMB[38][10] ) );
  FA_X1 \mult_22/S2_38_9  ( .A(\mult_22/ab[38][9] ), .B(
        \mult_22/CARRYB[37][9] ), .CI(\mult_22/SUMB[37][10] ), .CO(
        \mult_22/CARRYB[38][9] ), .S(\mult_22/SUMB[38][9] ) );
  FA_X1 \mult_22/S2_38_8  ( .A(\mult_22/ab[38][8] ), .B(
        \mult_22/CARRYB[37][8] ), .CI(\mult_22/SUMB[37][9] ), .CO(
        \mult_22/CARRYB[38][8] ), .S(\mult_22/SUMB[38][8] ) );
  FA_X1 \mult_22/S2_38_7  ( .A(\mult_22/ab[38][7] ), .B(
        \mult_22/CARRYB[37][7] ), .CI(\mult_22/SUMB[37][8] ), .CO(
        \mult_22/CARRYB[38][7] ), .S(\mult_22/SUMB[38][7] ) );
  FA_X1 \mult_22/S2_38_6  ( .A(\mult_22/ab[38][6] ), .B(
        \mult_22/CARRYB[37][6] ), .CI(\mult_22/SUMB[37][7] ), .CO(
        \mult_22/CARRYB[38][6] ), .S(\mult_22/SUMB[38][6] ) );
  FA_X1 \mult_22/S2_38_5  ( .A(\mult_22/ab[38][5] ), .B(
        \mult_22/CARRYB[37][5] ), .CI(\mult_22/SUMB[37][6] ), .CO(
        \mult_22/CARRYB[38][5] ), .S(\mult_22/SUMB[38][5] ) );
  FA_X1 \mult_22/S2_38_4  ( .A(\mult_22/ab[38][4] ), .B(
        \mult_22/CARRYB[37][4] ), .CI(\mult_22/SUMB[37][5] ), .CO(
        \mult_22/CARRYB[38][4] ), .S(\mult_22/SUMB[38][4] ) );
  FA_X1 \mult_22/S2_38_3  ( .A(\mult_22/ab[38][3] ), .B(
        \mult_22/CARRYB[37][3] ), .CI(\mult_22/SUMB[37][4] ), .CO(
        \mult_22/CARRYB[38][3] ), .S(\mult_22/SUMB[38][3] ) );
  FA_X1 \mult_22/S2_38_2  ( .A(\mult_22/ab[38][2] ), .B(
        \mult_22/CARRYB[37][2] ), .CI(\mult_22/SUMB[37][3] ), .CO(
        \mult_22/CARRYB[38][2] ), .S(\mult_22/SUMB[38][2] ) );
  FA_X1 \mult_22/S2_38_1  ( .A(\mult_22/ab[38][1] ), .B(
        \mult_22/CARRYB[37][1] ), .CI(\mult_22/SUMB[37][2] ), .CO(
        \mult_22/CARRYB[38][1] ), .S(\mult_22/SUMB[38][1] ) );
  FA_X1 \mult_22/S1_38_0  ( .A(\mult_22/ab[38][0] ), .B(
        \mult_22/CARRYB[37][0] ), .CI(\mult_22/SUMB[37][1] ), .CO(
        \mult_22/CARRYB[38][0] ), .S(N166) );
  FA_X1 \mult_22/S3_39_62  ( .A(\mult_22/ab[39][62] ), .B(
        \mult_22/CARRYB[38][62] ), .CI(\mult_22/ab[38][63] ), .CO(
        \mult_22/CARRYB[39][62] ), .S(\mult_22/SUMB[39][62] ) );
  FA_X1 \mult_22/S2_39_61  ( .A(\mult_22/ab[39][61] ), .B(
        \mult_22/CARRYB[38][61] ), .CI(\mult_22/SUMB[38][62] ), .CO(
        \mult_22/CARRYB[39][61] ), .S(\mult_22/SUMB[39][61] ) );
  FA_X1 \mult_22/S2_39_60  ( .A(\mult_22/ab[39][60] ), .B(
        \mult_22/CARRYB[38][60] ), .CI(\mult_22/SUMB[38][61] ), .CO(
        \mult_22/CARRYB[39][60] ), .S(\mult_22/SUMB[39][60] ) );
  FA_X1 \mult_22/S2_39_59  ( .A(\mult_22/ab[39][59] ), .B(
        \mult_22/CARRYB[38][59] ), .CI(\mult_22/SUMB[38][60] ), .CO(
        \mult_22/CARRYB[39][59] ), .S(\mult_22/SUMB[39][59] ) );
  FA_X1 \mult_22/S2_39_58  ( .A(\mult_22/ab[39][58] ), .B(
        \mult_22/CARRYB[38][58] ), .CI(\mult_22/SUMB[38][59] ), .CO(
        \mult_22/CARRYB[39][58] ), .S(\mult_22/SUMB[39][58] ) );
  FA_X1 \mult_22/S2_39_57  ( .A(\mult_22/ab[39][57] ), .B(
        \mult_22/CARRYB[38][57] ), .CI(\mult_22/SUMB[38][58] ), .CO(
        \mult_22/CARRYB[39][57] ), .S(\mult_22/SUMB[39][57] ) );
  FA_X1 \mult_22/S2_39_56  ( .A(\mult_22/ab[39][56] ), .B(
        \mult_22/CARRYB[38][56] ), .CI(\mult_22/SUMB[38][57] ), .CO(
        \mult_22/CARRYB[39][56] ), .S(\mult_22/SUMB[39][56] ) );
  FA_X1 \mult_22/S2_39_55  ( .A(\mult_22/ab[39][55] ), .B(
        \mult_22/CARRYB[38][55] ), .CI(\mult_22/SUMB[38][56] ), .CO(
        \mult_22/CARRYB[39][55] ), .S(\mult_22/SUMB[39][55] ) );
  FA_X1 \mult_22/S2_39_54  ( .A(\mult_22/ab[39][54] ), .B(
        \mult_22/CARRYB[38][54] ), .CI(\mult_22/SUMB[38][55] ), .CO(
        \mult_22/CARRYB[39][54] ), .S(\mult_22/SUMB[39][54] ) );
  FA_X1 \mult_22/S2_39_53  ( .A(\mult_22/ab[39][53] ), .B(
        \mult_22/CARRYB[38][53] ), .CI(\mult_22/SUMB[38][54] ), .CO(
        \mult_22/CARRYB[39][53] ), .S(\mult_22/SUMB[39][53] ) );
  FA_X1 \mult_22/S2_39_52  ( .A(\mult_22/ab[39][52] ), .B(
        \mult_22/CARRYB[38][52] ), .CI(\mult_22/SUMB[38][53] ), .CO(
        \mult_22/CARRYB[39][52] ), .S(\mult_22/SUMB[39][52] ) );
  FA_X1 \mult_22/S2_39_51  ( .A(\mult_22/ab[39][51] ), .B(
        \mult_22/CARRYB[38][51] ), .CI(\mult_22/SUMB[38][52] ), .CO(
        \mult_22/CARRYB[39][51] ), .S(\mult_22/SUMB[39][51] ) );
  FA_X1 \mult_22/S2_39_50  ( .A(\mult_22/ab[39][50] ), .B(
        \mult_22/CARRYB[38][50] ), .CI(\mult_22/SUMB[38][51] ), .CO(
        \mult_22/CARRYB[39][50] ), .S(\mult_22/SUMB[39][50] ) );
  FA_X1 \mult_22/S2_39_49  ( .A(\mult_22/ab[39][49] ), .B(
        \mult_22/CARRYB[38][49] ), .CI(\mult_22/SUMB[38][50] ), .CO(
        \mult_22/CARRYB[39][49] ), .S(\mult_22/SUMB[39][49] ) );
  FA_X1 \mult_22/S2_39_48  ( .A(\mult_22/ab[39][48] ), .B(
        \mult_22/CARRYB[38][48] ), .CI(\mult_22/SUMB[38][49] ), .CO(
        \mult_22/CARRYB[39][48] ), .S(\mult_22/SUMB[39][48] ) );
  FA_X1 \mult_22/S2_39_47  ( .A(\mult_22/ab[39][47] ), .B(
        \mult_22/CARRYB[38][47] ), .CI(\mult_22/SUMB[38][48] ), .CO(
        \mult_22/CARRYB[39][47] ), .S(\mult_22/SUMB[39][47] ) );
  FA_X1 \mult_22/S2_39_46  ( .A(\mult_22/ab[39][46] ), .B(
        \mult_22/CARRYB[38][46] ), .CI(\mult_22/SUMB[38][47] ), .CO(
        \mult_22/CARRYB[39][46] ), .S(\mult_22/SUMB[39][46] ) );
  FA_X1 \mult_22/S2_39_45  ( .A(\mult_22/ab[39][45] ), .B(
        \mult_22/CARRYB[38][45] ), .CI(\mult_22/SUMB[38][46] ), .CO(
        \mult_22/CARRYB[39][45] ), .S(\mult_22/SUMB[39][45] ) );
  FA_X1 \mult_22/S2_39_44  ( .A(\mult_22/ab[39][44] ), .B(
        \mult_22/CARRYB[38][44] ), .CI(\mult_22/SUMB[38][45] ), .CO(
        \mult_22/CARRYB[39][44] ), .S(\mult_22/SUMB[39][44] ) );
  FA_X1 \mult_22/S2_39_43  ( .A(\mult_22/ab[39][43] ), .B(
        \mult_22/CARRYB[38][43] ), .CI(\mult_22/SUMB[38][44] ), .CO(
        \mult_22/CARRYB[39][43] ), .S(\mult_22/SUMB[39][43] ) );
  FA_X1 \mult_22/S2_39_42  ( .A(\mult_22/ab[39][42] ), .B(
        \mult_22/CARRYB[38][42] ), .CI(\mult_22/SUMB[38][43] ), .CO(
        \mult_22/CARRYB[39][42] ), .S(\mult_22/SUMB[39][42] ) );
  FA_X1 \mult_22/S2_39_41  ( .A(\mult_22/ab[39][41] ), .B(
        \mult_22/CARRYB[38][41] ), .CI(\mult_22/SUMB[38][42] ), .CO(
        \mult_22/CARRYB[39][41] ), .S(\mult_22/SUMB[39][41] ) );
  FA_X1 \mult_22/S2_39_40  ( .A(\mult_22/ab[39][40] ), .B(
        \mult_22/CARRYB[38][40] ), .CI(\mult_22/SUMB[38][41] ), .CO(
        \mult_22/CARRYB[39][40] ), .S(\mult_22/SUMB[39][40] ) );
  FA_X1 \mult_22/S2_39_39  ( .A(\mult_22/ab[39][39] ), .B(
        \mult_22/CARRYB[38][39] ), .CI(\mult_22/SUMB[38][40] ), .CO(
        \mult_22/CARRYB[39][39] ), .S(\mult_22/SUMB[39][39] ) );
  FA_X1 \mult_22/S2_39_38  ( .A(\mult_22/ab[39][38] ), .B(
        \mult_22/CARRYB[38][38] ), .CI(\mult_22/SUMB[38][39] ), .CO(
        \mult_22/CARRYB[39][38] ), .S(\mult_22/SUMB[39][38] ) );
  FA_X1 \mult_22/S2_39_37  ( .A(\mult_22/ab[39][37] ), .B(
        \mult_22/CARRYB[38][37] ), .CI(\mult_22/SUMB[38][38] ), .CO(
        \mult_22/CARRYB[39][37] ), .S(\mult_22/SUMB[39][37] ) );
  FA_X1 \mult_22/S2_39_36  ( .A(\mult_22/ab[39][36] ), .B(
        \mult_22/CARRYB[38][36] ), .CI(\mult_22/SUMB[38][37] ), .CO(
        \mult_22/CARRYB[39][36] ), .S(\mult_22/SUMB[39][36] ) );
  FA_X1 \mult_22/S2_39_35  ( .A(\mult_22/ab[39][35] ), .B(
        \mult_22/CARRYB[38][35] ), .CI(\mult_22/SUMB[38][36] ), .CO(
        \mult_22/CARRYB[39][35] ), .S(\mult_22/SUMB[39][35] ) );
  FA_X1 \mult_22/S2_39_34  ( .A(\mult_22/ab[39][34] ), .B(
        \mult_22/CARRYB[38][34] ), .CI(\mult_22/SUMB[38][35] ), .CO(
        \mult_22/CARRYB[39][34] ), .S(\mult_22/SUMB[39][34] ) );
  FA_X1 \mult_22/S2_39_33  ( .A(\mult_22/ab[39][33] ), .B(
        \mult_22/CARRYB[38][33] ), .CI(\mult_22/SUMB[38][34] ), .CO(
        \mult_22/CARRYB[39][33] ), .S(\mult_22/SUMB[39][33] ) );
  FA_X1 \mult_22/S2_39_32  ( .A(\mult_22/ab[39][32] ), .B(
        \mult_22/CARRYB[38][32] ), .CI(\mult_22/SUMB[38][33] ), .CO(
        \mult_22/CARRYB[39][32] ), .S(\mult_22/SUMB[39][32] ) );
  FA_X1 \mult_22/S2_39_31  ( .A(\mult_22/ab[39][31] ), .B(
        \mult_22/CARRYB[38][31] ), .CI(\mult_22/SUMB[38][32] ), .CO(
        \mult_22/CARRYB[39][31] ), .S(\mult_22/SUMB[39][31] ) );
  FA_X1 \mult_22/S2_39_30  ( .A(\mult_22/ab[39][30] ), .B(
        \mult_22/CARRYB[38][30] ), .CI(\mult_22/SUMB[38][31] ), .CO(
        \mult_22/CARRYB[39][30] ), .S(\mult_22/SUMB[39][30] ) );
  FA_X1 \mult_22/S2_39_29  ( .A(\mult_22/ab[39][29] ), .B(
        \mult_22/CARRYB[38][29] ), .CI(\mult_22/SUMB[38][30] ), .CO(
        \mult_22/CARRYB[39][29] ), .S(\mult_22/SUMB[39][29] ) );
  FA_X1 \mult_22/S2_39_28  ( .A(\mult_22/CARRYB[38][28] ), .B(
        \mult_22/ab[39][28] ), .CI(\mult_22/SUMB[38][29] ), .CO(
        \mult_22/CARRYB[39][28] ), .S(\mult_22/SUMB[39][28] ) );
  FA_X1 \mult_22/S2_39_27  ( .A(\mult_22/ab[39][27] ), .B(
        \mult_22/CARRYB[38][27] ), .CI(\mult_22/SUMB[38][28] ), .CO(
        \mult_22/CARRYB[39][27] ), .S(\mult_22/SUMB[39][27] ) );
  FA_X1 \mult_22/S2_39_26  ( .A(\mult_22/ab[39][26] ), .B(
        \mult_22/CARRYB[38][26] ), .CI(\mult_22/SUMB[38][27] ), .CO(
        \mult_22/CARRYB[39][26] ), .S(\mult_22/SUMB[39][26] ) );
  FA_X1 \mult_22/S2_39_25  ( .A(\mult_22/ab[39][25] ), .B(
        \mult_22/CARRYB[38][25] ), .CI(\mult_22/SUMB[38][26] ), .CO(
        \mult_22/CARRYB[39][25] ), .S(\mult_22/SUMB[39][25] ) );
  FA_X1 \mult_22/S2_39_24  ( .A(\mult_22/ab[39][24] ), .B(
        \mult_22/CARRYB[38][24] ), .CI(\mult_22/SUMB[38][25] ), .CO(
        \mult_22/CARRYB[39][24] ), .S(\mult_22/SUMB[39][24] ) );
  FA_X1 \mult_22/S2_39_23  ( .A(\mult_22/ab[39][23] ), .B(
        \mult_22/CARRYB[38][23] ), .CI(\mult_22/SUMB[38][24] ), .CO(
        \mult_22/CARRYB[39][23] ), .S(\mult_22/SUMB[39][23] ) );
  FA_X1 \mult_22/S2_39_22  ( .A(\mult_22/ab[39][22] ), .B(
        \mult_22/CARRYB[38][22] ), .CI(\mult_22/SUMB[38][23] ), .CO(
        \mult_22/CARRYB[39][22] ), .S(\mult_22/SUMB[39][22] ) );
  FA_X1 \mult_22/S2_39_21  ( .A(\mult_22/CARRYB[38][21] ), .B(
        \mult_22/ab[39][21] ), .CI(\mult_22/SUMB[38][22] ), .CO(
        \mult_22/CARRYB[39][21] ), .S(\mult_22/SUMB[39][21] ) );
  FA_X1 \mult_22/S2_39_20  ( .A(\mult_22/ab[39][20] ), .B(
        \mult_22/CARRYB[38][20] ), .CI(\mult_22/SUMB[38][21] ), .CO(
        \mult_22/CARRYB[39][20] ), .S(\mult_22/SUMB[39][20] ) );
  FA_X1 \mult_22/S2_39_19  ( .A(\mult_22/ab[39][19] ), .B(
        \mult_22/CARRYB[38][19] ), .CI(\mult_22/SUMB[38][20] ), .CO(
        \mult_22/CARRYB[39][19] ), .S(\mult_22/SUMB[39][19] ) );
  FA_X1 \mult_22/S2_39_18  ( .A(\mult_22/ab[39][18] ), .B(
        \mult_22/CARRYB[38][18] ), .CI(\mult_22/SUMB[38][19] ), .CO(
        \mult_22/CARRYB[39][18] ), .S(\mult_22/SUMB[39][18] ) );
  FA_X1 \mult_22/S2_39_17  ( .A(\mult_22/ab[39][17] ), .B(
        \mult_22/CARRYB[38][17] ), .CI(\mult_22/SUMB[38][18] ), .CO(
        \mult_22/CARRYB[39][17] ), .S(\mult_22/SUMB[39][17] ) );
  FA_X1 \mult_22/S2_39_16  ( .A(\mult_22/ab[39][16] ), .B(
        \mult_22/CARRYB[38][16] ), .CI(\mult_22/SUMB[38][17] ), .CO(
        \mult_22/CARRYB[39][16] ), .S(\mult_22/SUMB[39][16] ) );
  FA_X1 \mult_22/S2_39_15  ( .A(\mult_22/ab[39][15] ), .B(
        \mult_22/CARRYB[38][15] ), .CI(\mult_22/SUMB[38][16] ), .CO(
        \mult_22/CARRYB[39][15] ), .S(\mult_22/SUMB[39][15] ) );
  FA_X1 \mult_22/S2_39_14  ( .A(\mult_22/ab[39][14] ), .B(
        \mult_22/CARRYB[38][14] ), .CI(\mult_22/SUMB[38][15] ), .CO(
        \mult_22/CARRYB[39][14] ), .S(\mult_22/SUMB[39][14] ) );
  FA_X1 \mult_22/S2_39_13  ( .A(\mult_22/ab[39][13] ), .B(
        \mult_22/CARRYB[38][13] ), .CI(\mult_22/SUMB[38][14] ), .CO(
        \mult_22/CARRYB[39][13] ), .S(\mult_22/SUMB[39][13] ) );
  FA_X1 \mult_22/S2_39_12  ( .A(\mult_22/ab[39][12] ), .B(
        \mult_22/CARRYB[38][12] ), .CI(\mult_22/SUMB[38][13] ), .CO(
        \mult_22/CARRYB[39][12] ), .S(\mult_22/SUMB[39][12] ) );
  FA_X1 \mult_22/S2_39_11  ( .A(\mult_22/ab[39][11] ), .B(
        \mult_22/CARRYB[38][11] ), .CI(\mult_22/SUMB[38][12] ), .CO(
        \mult_22/CARRYB[39][11] ), .S(\mult_22/SUMB[39][11] ) );
  FA_X1 \mult_22/S2_39_10  ( .A(\mult_22/ab[39][10] ), .B(
        \mult_22/CARRYB[38][10] ), .CI(\mult_22/SUMB[38][11] ), .CO(
        \mult_22/CARRYB[39][10] ), .S(\mult_22/SUMB[39][10] ) );
  FA_X1 \mult_22/S2_39_9  ( .A(\mult_22/ab[39][9] ), .B(
        \mult_22/CARRYB[38][9] ), .CI(\mult_22/SUMB[38][10] ), .CO(
        \mult_22/CARRYB[39][9] ), .S(\mult_22/SUMB[39][9] ) );
  FA_X1 \mult_22/S2_39_8  ( .A(\mult_22/ab[39][8] ), .B(
        \mult_22/CARRYB[38][8] ), .CI(\mult_22/SUMB[38][9] ), .CO(
        \mult_22/CARRYB[39][8] ), .S(\mult_22/SUMB[39][8] ) );
  FA_X1 \mult_22/S2_39_7  ( .A(\mult_22/ab[39][7] ), .B(
        \mult_22/CARRYB[38][7] ), .CI(\mult_22/SUMB[38][8] ), .CO(
        \mult_22/CARRYB[39][7] ), .S(\mult_22/SUMB[39][7] ) );
  FA_X1 \mult_22/S2_39_6  ( .A(\mult_22/ab[39][6] ), .B(
        \mult_22/CARRYB[38][6] ), .CI(\mult_22/SUMB[38][7] ), .CO(
        \mult_22/CARRYB[39][6] ), .S(\mult_22/SUMB[39][6] ) );
  FA_X1 \mult_22/S2_39_5  ( .A(\mult_22/ab[39][5] ), .B(
        \mult_22/CARRYB[38][5] ), .CI(\mult_22/SUMB[38][6] ), .CO(
        \mult_22/CARRYB[39][5] ), .S(\mult_22/SUMB[39][5] ) );
  FA_X1 \mult_22/S2_39_4  ( .A(\mult_22/ab[39][4] ), .B(
        \mult_22/CARRYB[38][4] ), .CI(\mult_22/SUMB[38][5] ), .CO(
        \mult_22/CARRYB[39][4] ), .S(\mult_22/SUMB[39][4] ) );
  FA_X1 \mult_22/S2_39_3  ( .A(\mult_22/ab[39][3] ), .B(
        \mult_22/CARRYB[38][3] ), .CI(\mult_22/SUMB[38][4] ), .CO(
        \mult_22/CARRYB[39][3] ), .S(\mult_22/SUMB[39][3] ) );
  FA_X1 \mult_22/S2_39_2  ( .A(\mult_22/ab[39][2] ), .B(
        \mult_22/CARRYB[38][2] ), .CI(\mult_22/SUMB[38][3] ), .CO(
        \mult_22/CARRYB[39][2] ), .S(\mult_22/SUMB[39][2] ) );
  FA_X1 \mult_22/S2_39_1  ( .A(\mult_22/ab[39][1] ), .B(
        \mult_22/CARRYB[38][1] ), .CI(\mult_22/SUMB[38][2] ), .CO(
        \mult_22/CARRYB[39][1] ), .S(\mult_22/SUMB[39][1] ) );
  FA_X1 \mult_22/S1_39_0  ( .A(\mult_22/ab[39][0] ), .B(
        \mult_22/CARRYB[38][0] ), .CI(\mult_22/SUMB[38][1] ), .CO(
        \mult_22/CARRYB[39][0] ), .S(N167) );
  FA_X1 \mult_22/S3_40_62  ( .A(\mult_22/ab[40][62] ), .B(
        \mult_22/CARRYB[39][62] ), .CI(\mult_22/ab[39][63] ), .CO(
        \mult_22/CARRYB[40][62] ), .S(\mult_22/SUMB[40][62] ) );
  FA_X1 \mult_22/S2_40_61  ( .A(\mult_22/ab[40][61] ), .B(
        \mult_22/CARRYB[39][61] ), .CI(\mult_22/SUMB[39][62] ), .CO(
        \mult_22/CARRYB[40][61] ), .S(\mult_22/SUMB[40][61] ) );
  FA_X1 \mult_22/S2_40_60  ( .A(\mult_22/ab[40][60] ), .B(
        \mult_22/CARRYB[39][60] ), .CI(\mult_22/SUMB[39][61] ), .CO(
        \mult_22/CARRYB[40][60] ), .S(\mult_22/SUMB[40][60] ) );
  FA_X1 \mult_22/S2_40_59  ( .A(\mult_22/ab[40][59] ), .B(
        \mult_22/CARRYB[39][59] ), .CI(\mult_22/SUMB[39][60] ), .CO(
        \mult_22/CARRYB[40][59] ), .S(\mult_22/SUMB[40][59] ) );
  FA_X1 \mult_22/S2_40_58  ( .A(\mult_22/ab[40][58] ), .B(
        \mult_22/CARRYB[39][58] ), .CI(\mult_22/SUMB[39][59] ), .CO(
        \mult_22/CARRYB[40][58] ), .S(\mult_22/SUMB[40][58] ) );
  FA_X1 \mult_22/S2_40_57  ( .A(\mult_22/ab[40][57] ), .B(
        \mult_22/CARRYB[39][57] ), .CI(\mult_22/SUMB[39][58] ), .CO(
        \mult_22/CARRYB[40][57] ), .S(\mult_22/SUMB[40][57] ) );
  FA_X1 \mult_22/S2_40_56  ( .A(\mult_22/ab[40][56] ), .B(
        \mult_22/CARRYB[39][56] ), .CI(\mult_22/SUMB[39][57] ), .CO(
        \mult_22/CARRYB[40][56] ), .S(\mult_22/SUMB[40][56] ) );
  FA_X1 \mult_22/S2_40_55  ( .A(\mult_22/ab[40][55] ), .B(
        \mult_22/CARRYB[39][55] ), .CI(\mult_22/SUMB[39][56] ), .CO(
        \mult_22/CARRYB[40][55] ), .S(\mult_22/SUMB[40][55] ) );
  FA_X1 \mult_22/S2_40_54  ( .A(\mult_22/ab[40][54] ), .B(
        \mult_22/CARRYB[39][54] ), .CI(\mult_22/SUMB[39][55] ), .CO(
        \mult_22/CARRYB[40][54] ), .S(\mult_22/SUMB[40][54] ) );
  FA_X1 \mult_22/S2_40_53  ( .A(\mult_22/ab[40][53] ), .B(
        \mult_22/CARRYB[39][53] ), .CI(\mult_22/SUMB[39][54] ), .CO(
        \mult_22/CARRYB[40][53] ), .S(\mult_22/SUMB[40][53] ) );
  FA_X1 \mult_22/S2_40_52  ( .A(\mult_22/ab[40][52] ), .B(
        \mult_22/CARRYB[39][52] ), .CI(\mult_22/SUMB[39][53] ), .CO(
        \mult_22/CARRYB[40][52] ), .S(\mult_22/SUMB[40][52] ) );
  FA_X1 \mult_22/S2_40_51  ( .A(\mult_22/ab[40][51] ), .B(
        \mult_22/CARRYB[39][51] ), .CI(\mult_22/SUMB[39][52] ), .CO(
        \mult_22/CARRYB[40][51] ), .S(\mult_22/SUMB[40][51] ) );
  FA_X1 \mult_22/S2_40_50  ( .A(\mult_22/ab[40][50] ), .B(
        \mult_22/CARRYB[39][50] ), .CI(\mult_22/SUMB[39][51] ), .CO(
        \mult_22/CARRYB[40][50] ), .S(\mult_22/SUMB[40][50] ) );
  FA_X1 \mult_22/S2_40_49  ( .A(\mult_22/ab[40][49] ), .B(
        \mult_22/CARRYB[39][49] ), .CI(\mult_22/SUMB[39][50] ), .CO(
        \mult_22/CARRYB[40][49] ), .S(\mult_22/SUMB[40][49] ) );
  FA_X1 \mult_22/S2_40_48  ( .A(\mult_22/ab[40][48] ), .B(
        \mult_22/CARRYB[39][48] ), .CI(\mult_22/SUMB[39][49] ), .CO(
        \mult_22/CARRYB[40][48] ), .S(\mult_22/SUMB[40][48] ) );
  FA_X1 \mult_22/S2_40_47  ( .A(\mult_22/ab[40][47] ), .B(
        \mult_22/CARRYB[39][47] ), .CI(\mult_22/SUMB[39][48] ), .CO(
        \mult_22/CARRYB[40][47] ), .S(\mult_22/SUMB[40][47] ) );
  FA_X1 \mult_22/S2_40_46  ( .A(\mult_22/ab[40][46] ), .B(
        \mult_22/CARRYB[39][46] ), .CI(\mult_22/SUMB[39][47] ), .CO(
        \mult_22/CARRYB[40][46] ), .S(\mult_22/SUMB[40][46] ) );
  FA_X1 \mult_22/S2_40_45  ( .A(\mult_22/ab[40][45] ), .B(
        \mult_22/CARRYB[39][45] ), .CI(\mult_22/SUMB[39][46] ), .CO(
        \mult_22/CARRYB[40][45] ), .S(\mult_22/SUMB[40][45] ) );
  FA_X1 \mult_22/S2_40_44  ( .A(\mult_22/ab[40][44] ), .B(
        \mult_22/CARRYB[39][44] ), .CI(\mult_22/SUMB[39][45] ), .CO(
        \mult_22/CARRYB[40][44] ), .S(\mult_22/SUMB[40][44] ) );
  FA_X1 \mult_22/S2_40_43  ( .A(\mult_22/ab[40][43] ), .B(
        \mult_22/CARRYB[39][43] ), .CI(\mult_22/SUMB[39][44] ), .CO(
        \mult_22/CARRYB[40][43] ), .S(\mult_22/SUMB[40][43] ) );
  FA_X1 \mult_22/S2_40_42  ( .A(\mult_22/ab[40][42] ), .B(
        \mult_22/CARRYB[39][42] ), .CI(\mult_22/SUMB[39][43] ), .CO(
        \mult_22/CARRYB[40][42] ), .S(\mult_22/SUMB[40][42] ) );
  FA_X1 \mult_22/S2_40_41  ( .A(\mult_22/ab[40][41] ), .B(
        \mult_22/CARRYB[39][41] ), .CI(\mult_22/SUMB[39][42] ), .CO(
        \mult_22/CARRYB[40][41] ), .S(\mult_22/SUMB[40][41] ) );
  FA_X1 \mult_22/S2_40_40  ( .A(\mult_22/ab[40][40] ), .B(
        \mult_22/CARRYB[39][40] ), .CI(\mult_22/SUMB[39][41] ), .CO(
        \mult_22/CARRYB[40][40] ), .S(\mult_22/SUMB[40][40] ) );
  FA_X1 \mult_22/S2_40_39  ( .A(\mult_22/ab[40][39] ), .B(
        \mult_22/CARRYB[39][39] ), .CI(\mult_22/SUMB[39][40] ), .CO(
        \mult_22/CARRYB[40][39] ), .S(\mult_22/SUMB[40][39] ) );
  FA_X1 \mult_22/S2_40_38  ( .A(\mult_22/ab[40][38] ), .B(
        \mult_22/CARRYB[39][38] ), .CI(\mult_22/SUMB[39][39] ), .CO(
        \mult_22/CARRYB[40][38] ), .S(\mult_22/SUMB[40][38] ) );
  FA_X1 \mult_22/S2_40_37  ( .A(\mult_22/ab[40][37] ), .B(
        \mult_22/CARRYB[39][37] ), .CI(\mult_22/SUMB[39][38] ), .CO(
        \mult_22/CARRYB[40][37] ), .S(\mult_22/SUMB[40][37] ) );
  FA_X1 \mult_22/S2_40_36  ( .A(\mult_22/ab[40][36] ), .B(
        \mult_22/CARRYB[39][36] ), .CI(\mult_22/SUMB[39][37] ), .CO(
        \mult_22/CARRYB[40][36] ), .S(\mult_22/SUMB[40][36] ) );
  FA_X1 \mult_22/S2_40_35  ( .A(\mult_22/ab[40][35] ), .B(
        \mult_22/CARRYB[39][35] ), .CI(\mult_22/SUMB[39][36] ), .CO(
        \mult_22/CARRYB[40][35] ), .S(\mult_22/SUMB[40][35] ) );
  FA_X1 \mult_22/S2_40_34  ( .A(\mult_22/ab[40][34] ), .B(
        \mult_22/CARRYB[39][34] ), .CI(\mult_22/SUMB[39][35] ), .CO(
        \mult_22/CARRYB[40][34] ), .S(\mult_22/SUMB[40][34] ) );
  FA_X1 \mult_22/S2_40_33  ( .A(\mult_22/ab[40][33] ), .B(
        \mult_22/CARRYB[39][33] ), .CI(\mult_22/SUMB[39][34] ), .CO(
        \mult_22/CARRYB[40][33] ), .S(\mult_22/SUMB[40][33] ) );
  FA_X1 \mult_22/S2_40_32  ( .A(\mult_22/ab[40][32] ), .B(
        \mult_22/CARRYB[39][32] ), .CI(\mult_22/SUMB[39][33] ), .CO(
        \mult_22/CARRYB[40][32] ), .S(\mult_22/SUMB[40][32] ) );
  FA_X1 \mult_22/S2_40_31  ( .A(\mult_22/ab[40][31] ), .B(
        \mult_22/CARRYB[39][31] ), .CI(\mult_22/SUMB[39][32] ), .CO(
        \mult_22/CARRYB[40][31] ), .S(\mult_22/SUMB[40][31] ) );
  FA_X1 \mult_22/S2_40_30  ( .A(\mult_22/ab[40][30] ), .B(
        \mult_22/CARRYB[39][30] ), .CI(\mult_22/SUMB[39][31] ), .CO(
        \mult_22/CARRYB[40][30] ), .S(\mult_22/SUMB[40][30] ) );
  FA_X1 \mult_22/S2_40_29  ( .A(\mult_22/ab[40][29] ), .B(
        \mult_22/CARRYB[39][29] ), .CI(\mult_22/SUMB[39][30] ), .CO(
        \mult_22/CARRYB[40][29] ), .S(\mult_22/SUMB[40][29] ) );
  FA_X1 \mult_22/S2_40_28  ( .A(\mult_22/ab[40][28] ), .B(
        \mult_22/CARRYB[39][28] ), .CI(\mult_22/SUMB[39][29] ), .CO(
        \mult_22/CARRYB[40][28] ), .S(\mult_22/SUMB[40][28] ) );
  FA_X1 \mult_22/S2_40_27  ( .A(\mult_22/ab[40][27] ), .B(
        \mult_22/CARRYB[39][27] ), .CI(\mult_22/SUMB[39][28] ), .CO(
        \mult_22/CARRYB[40][27] ), .S(\mult_22/SUMB[40][27] ) );
  FA_X1 \mult_22/S2_40_26  ( .A(\mult_22/CARRYB[39][26] ), .B(
        \mult_22/ab[40][26] ), .CI(\mult_22/SUMB[39][27] ), .CO(
        \mult_22/CARRYB[40][26] ), .S(\mult_22/SUMB[40][26] ) );
  FA_X1 \mult_22/S2_40_25  ( .A(\mult_22/ab[40][25] ), .B(
        \mult_22/CARRYB[39][25] ), .CI(\mult_22/SUMB[39][26] ), .CO(
        \mult_22/CARRYB[40][25] ), .S(\mult_22/SUMB[40][25] ) );
  FA_X1 \mult_22/S2_40_24  ( .A(\mult_22/ab[40][24] ), .B(
        \mult_22/CARRYB[39][24] ), .CI(\mult_22/SUMB[39][25] ), .CO(
        \mult_22/CARRYB[40][24] ), .S(\mult_22/SUMB[40][24] ) );
  FA_X1 \mult_22/S2_40_23  ( .A(\mult_22/ab[40][23] ), .B(
        \mult_22/CARRYB[39][23] ), .CI(\mult_22/SUMB[39][24] ), .CO(
        \mult_22/CARRYB[40][23] ), .S(\mult_22/SUMB[40][23] ) );
  FA_X1 \mult_22/S2_40_22  ( .A(\mult_22/ab[40][22] ), .B(
        \mult_22/CARRYB[39][22] ), .CI(\mult_22/SUMB[39][23] ), .CO(
        \mult_22/CARRYB[40][22] ), .S(\mult_22/SUMB[40][22] ) );
  FA_X1 \mult_22/S2_40_21  ( .A(\mult_22/ab[40][21] ), .B(
        \mult_22/CARRYB[39][21] ), .CI(\mult_22/SUMB[39][22] ), .CO(
        \mult_22/CARRYB[40][21] ), .S(\mult_22/SUMB[40][21] ) );
  FA_X1 \mult_22/S2_40_20  ( .A(\mult_22/ab[40][20] ), .B(
        \mult_22/CARRYB[39][20] ), .CI(\mult_22/SUMB[39][21] ), .CO(
        \mult_22/CARRYB[40][20] ), .S(\mult_22/SUMB[40][20] ) );
  FA_X1 \mult_22/S2_40_19  ( .A(\mult_22/ab[40][19] ), .B(
        \mult_22/CARRYB[39][19] ), .CI(\mult_22/SUMB[39][20] ), .CO(
        \mult_22/CARRYB[40][19] ), .S(\mult_22/SUMB[40][19] ) );
  FA_X1 \mult_22/S2_40_18  ( .A(\mult_22/ab[40][18] ), .B(
        \mult_22/CARRYB[39][18] ), .CI(\mult_22/SUMB[39][19] ), .CO(
        \mult_22/CARRYB[40][18] ), .S(\mult_22/SUMB[40][18] ) );
  FA_X1 \mult_22/S2_40_17  ( .A(\mult_22/ab[40][17] ), .B(
        \mult_22/CARRYB[39][17] ), .CI(\mult_22/SUMB[39][18] ), .CO(
        \mult_22/CARRYB[40][17] ), .S(\mult_22/SUMB[40][17] ) );
  FA_X1 \mult_22/S2_40_16  ( .A(\mult_22/ab[40][16] ), .B(
        \mult_22/CARRYB[39][16] ), .CI(\mult_22/SUMB[39][17] ), .CO(
        \mult_22/CARRYB[40][16] ), .S(\mult_22/SUMB[40][16] ) );
  FA_X1 \mult_22/S2_40_15  ( .A(\mult_22/ab[40][15] ), .B(
        \mult_22/CARRYB[39][15] ), .CI(\mult_22/SUMB[39][16] ), .CO(
        \mult_22/CARRYB[40][15] ), .S(\mult_22/SUMB[40][15] ) );
  FA_X1 \mult_22/S2_40_14  ( .A(\mult_22/ab[40][14] ), .B(
        \mult_22/CARRYB[39][14] ), .CI(\mult_22/SUMB[39][15] ), .CO(
        \mult_22/CARRYB[40][14] ), .S(\mult_22/SUMB[40][14] ) );
  FA_X1 \mult_22/S2_40_13  ( .A(\mult_22/ab[40][13] ), .B(
        \mult_22/CARRYB[39][13] ), .CI(\mult_22/SUMB[39][14] ), .CO(
        \mult_22/CARRYB[40][13] ), .S(\mult_22/SUMB[40][13] ) );
  FA_X1 \mult_22/S2_40_12  ( .A(\mult_22/ab[40][12] ), .B(
        \mult_22/CARRYB[39][12] ), .CI(\mult_22/SUMB[39][13] ), .CO(
        \mult_22/CARRYB[40][12] ), .S(\mult_22/SUMB[40][12] ) );
  FA_X1 \mult_22/S2_40_11  ( .A(\mult_22/ab[40][11] ), .B(
        \mult_22/CARRYB[39][11] ), .CI(\mult_22/SUMB[39][12] ), .CO(
        \mult_22/CARRYB[40][11] ), .S(\mult_22/SUMB[40][11] ) );
  FA_X1 \mult_22/S2_40_10  ( .A(\mult_22/ab[40][10] ), .B(
        \mult_22/CARRYB[39][10] ), .CI(\mult_22/SUMB[39][11] ), .CO(
        \mult_22/CARRYB[40][10] ), .S(\mult_22/SUMB[40][10] ) );
  FA_X1 \mult_22/S2_40_9  ( .A(\mult_22/ab[40][9] ), .B(
        \mult_22/CARRYB[39][9] ), .CI(\mult_22/SUMB[39][10] ), .CO(
        \mult_22/CARRYB[40][9] ), .S(\mult_22/SUMB[40][9] ) );
  FA_X1 \mult_22/S2_40_8  ( .A(\mult_22/ab[40][8] ), .B(
        \mult_22/CARRYB[39][8] ), .CI(\mult_22/SUMB[39][9] ), .CO(
        \mult_22/CARRYB[40][8] ), .S(\mult_22/SUMB[40][8] ) );
  FA_X1 \mult_22/S2_40_7  ( .A(\mult_22/ab[40][7] ), .B(
        \mult_22/CARRYB[39][7] ), .CI(\mult_22/SUMB[39][8] ), .CO(
        \mult_22/CARRYB[40][7] ), .S(\mult_22/SUMB[40][7] ) );
  FA_X1 \mult_22/S2_40_6  ( .A(\mult_22/ab[40][6] ), .B(
        \mult_22/CARRYB[39][6] ), .CI(\mult_22/SUMB[39][7] ), .CO(
        \mult_22/CARRYB[40][6] ), .S(\mult_22/SUMB[40][6] ) );
  FA_X1 \mult_22/S2_40_5  ( .A(\mult_22/ab[40][5] ), .B(
        \mult_22/CARRYB[39][5] ), .CI(\mult_22/SUMB[39][6] ), .CO(
        \mult_22/CARRYB[40][5] ), .S(\mult_22/SUMB[40][5] ) );
  FA_X1 \mult_22/S2_40_4  ( .A(\mult_22/ab[40][4] ), .B(
        \mult_22/CARRYB[39][4] ), .CI(\mult_22/SUMB[39][5] ), .CO(
        \mult_22/CARRYB[40][4] ), .S(\mult_22/SUMB[40][4] ) );
  FA_X1 \mult_22/S2_40_3  ( .A(\mult_22/ab[40][3] ), .B(
        \mult_22/CARRYB[39][3] ), .CI(\mult_22/SUMB[39][4] ), .CO(
        \mult_22/CARRYB[40][3] ), .S(\mult_22/SUMB[40][3] ) );
  FA_X1 \mult_22/S2_40_2  ( .A(\mult_22/ab[40][2] ), .B(
        \mult_22/CARRYB[39][2] ), .CI(\mult_22/SUMB[39][3] ), .CO(
        \mult_22/CARRYB[40][2] ), .S(\mult_22/SUMB[40][2] ) );
  FA_X1 \mult_22/S2_40_1  ( .A(\mult_22/ab[40][1] ), .B(
        \mult_22/CARRYB[39][1] ), .CI(\mult_22/SUMB[39][2] ), .CO(
        \mult_22/CARRYB[40][1] ), .S(\mult_22/SUMB[40][1] ) );
  FA_X1 \mult_22/S1_40_0  ( .A(\mult_22/ab[40][0] ), .B(
        \mult_22/CARRYB[39][0] ), .CI(\mult_22/SUMB[39][1] ), .CO(
        \mult_22/CARRYB[40][0] ), .S(N168) );
  FA_X1 \mult_22/S3_41_62  ( .A(\mult_22/ab[41][62] ), .B(
        \mult_22/CARRYB[40][62] ), .CI(\mult_22/ab[40][63] ), .CO(
        \mult_22/CARRYB[41][62] ), .S(\mult_22/SUMB[41][62] ) );
  FA_X1 \mult_22/S2_41_61  ( .A(\mult_22/ab[41][61] ), .B(
        \mult_22/CARRYB[40][61] ), .CI(\mult_22/SUMB[40][62] ), .CO(
        \mult_22/CARRYB[41][61] ), .S(\mult_22/SUMB[41][61] ) );
  FA_X1 \mult_22/S2_41_60  ( .A(\mult_22/ab[41][60] ), .B(
        \mult_22/CARRYB[40][60] ), .CI(\mult_22/SUMB[40][61] ), .CO(
        \mult_22/CARRYB[41][60] ), .S(\mult_22/SUMB[41][60] ) );
  FA_X1 \mult_22/S2_41_59  ( .A(\mult_22/ab[41][59] ), .B(
        \mult_22/CARRYB[40][59] ), .CI(\mult_22/SUMB[40][60] ), .CO(
        \mult_22/CARRYB[41][59] ), .S(\mult_22/SUMB[41][59] ) );
  FA_X1 \mult_22/S2_41_58  ( .A(\mult_22/ab[41][58] ), .B(
        \mult_22/CARRYB[40][58] ), .CI(\mult_22/SUMB[40][59] ), .CO(
        \mult_22/CARRYB[41][58] ), .S(\mult_22/SUMB[41][58] ) );
  FA_X1 \mult_22/S2_41_57  ( .A(\mult_22/ab[41][57] ), .B(
        \mult_22/CARRYB[40][57] ), .CI(\mult_22/SUMB[40][58] ), .CO(
        \mult_22/CARRYB[41][57] ), .S(\mult_22/SUMB[41][57] ) );
  FA_X1 \mult_22/S2_41_56  ( .A(\mult_22/ab[41][56] ), .B(
        \mult_22/CARRYB[40][56] ), .CI(\mult_22/SUMB[40][57] ), .CO(
        \mult_22/CARRYB[41][56] ), .S(\mult_22/SUMB[41][56] ) );
  FA_X1 \mult_22/S2_41_55  ( .A(\mult_22/ab[41][55] ), .B(
        \mult_22/CARRYB[40][55] ), .CI(\mult_22/SUMB[40][56] ), .CO(
        \mult_22/CARRYB[41][55] ), .S(\mult_22/SUMB[41][55] ) );
  FA_X1 \mult_22/S2_41_54  ( .A(\mult_22/ab[41][54] ), .B(
        \mult_22/CARRYB[40][54] ), .CI(\mult_22/SUMB[40][55] ), .CO(
        \mult_22/CARRYB[41][54] ), .S(\mult_22/SUMB[41][54] ) );
  FA_X1 \mult_22/S2_41_53  ( .A(\mult_22/ab[41][53] ), .B(
        \mult_22/CARRYB[40][53] ), .CI(\mult_22/SUMB[40][54] ), .CO(
        \mult_22/CARRYB[41][53] ), .S(\mult_22/SUMB[41][53] ) );
  FA_X1 \mult_22/S2_41_52  ( .A(\mult_22/ab[41][52] ), .B(
        \mult_22/CARRYB[40][52] ), .CI(\mult_22/SUMB[40][53] ), .CO(
        \mult_22/CARRYB[41][52] ), .S(\mult_22/SUMB[41][52] ) );
  FA_X1 \mult_22/S2_41_51  ( .A(\mult_22/ab[41][51] ), .B(
        \mult_22/CARRYB[40][51] ), .CI(\mult_22/SUMB[40][52] ), .CO(
        \mult_22/CARRYB[41][51] ), .S(\mult_22/SUMB[41][51] ) );
  FA_X1 \mult_22/S2_41_50  ( .A(\mult_22/ab[41][50] ), .B(
        \mult_22/CARRYB[40][50] ), .CI(\mult_22/SUMB[40][51] ), .CO(
        \mult_22/CARRYB[41][50] ), .S(\mult_22/SUMB[41][50] ) );
  FA_X1 \mult_22/S2_41_49  ( .A(\mult_22/ab[41][49] ), .B(
        \mult_22/CARRYB[40][49] ), .CI(\mult_22/SUMB[40][50] ), .CO(
        \mult_22/CARRYB[41][49] ), .S(\mult_22/SUMB[41][49] ) );
  FA_X1 \mult_22/S2_41_48  ( .A(\mult_22/ab[41][48] ), .B(
        \mult_22/CARRYB[40][48] ), .CI(\mult_22/SUMB[40][49] ), .CO(
        \mult_22/CARRYB[41][48] ), .S(\mult_22/SUMB[41][48] ) );
  FA_X1 \mult_22/S2_41_47  ( .A(\mult_22/ab[41][47] ), .B(
        \mult_22/CARRYB[40][47] ), .CI(\mult_22/SUMB[40][48] ), .CO(
        \mult_22/CARRYB[41][47] ), .S(\mult_22/SUMB[41][47] ) );
  FA_X1 \mult_22/S2_41_46  ( .A(\mult_22/ab[41][46] ), .B(
        \mult_22/CARRYB[40][46] ), .CI(\mult_22/SUMB[40][47] ), .CO(
        \mult_22/CARRYB[41][46] ), .S(\mult_22/SUMB[41][46] ) );
  FA_X1 \mult_22/S2_41_45  ( .A(\mult_22/ab[41][45] ), .B(
        \mult_22/CARRYB[40][45] ), .CI(\mult_22/SUMB[40][46] ), .CO(
        \mult_22/CARRYB[41][45] ), .S(\mult_22/SUMB[41][45] ) );
  FA_X1 \mult_22/S2_41_44  ( .A(\mult_22/ab[41][44] ), .B(
        \mult_22/CARRYB[40][44] ), .CI(\mult_22/SUMB[40][45] ), .CO(
        \mult_22/CARRYB[41][44] ), .S(\mult_22/SUMB[41][44] ) );
  FA_X1 \mult_22/S2_41_43  ( .A(\mult_22/ab[41][43] ), .B(
        \mult_22/CARRYB[40][43] ), .CI(\mult_22/SUMB[40][44] ), .CO(
        \mult_22/CARRYB[41][43] ), .S(\mult_22/SUMB[41][43] ) );
  FA_X1 \mult_22/S2_41_42  ( .A(\mult_22/ab[41][42] ), .B(
        \mult_22/CARRYB[40][42] ), .CI(\mult_22/SUMB[40][43] ), .CO(
        \mult_22/CARRYB[41][42] ), .S(\mult_22/SUMB[41][42] ) );
  FA_X1 \mult_22/S2_41_41  ( .A(\mult_22/ab[41][41] ), .B(
        \mult_22/CARRYB[40][41] ), .CI(\mult_22/SUMB[40][42] ), .CO(
        \mult_22/CARRYB[41][41] ), .S(\mult_22/SUMB[41][41] ) );
  FA_X1 \mult_22/S2_41_40  ( .A(\mult_22/ab[41][40] ), .B(
        \mult_22/CARRYB[40][40] ), .CI(\mult_22/SUMB[40][41] ), .CO(
        \mult_22/CARRYB[41][40] ), .S(\mult_22/SUMB[41][40] ) );
  FA_X1 \mult_22/S2_41_39  ( .A(\mult_22/ab[41][39] ), .B(
        \mult_22/CARRYB[40][39] ), .CI(\mult_22/SUMB[40][40] ), .CO(
        \mult_22/CARRYB[41][39] ), .S(\mult_22/SUMB[41][39] ) );
  FA_X1 \mult_22/S2_41_38  ( .A(\mult_22/ab[41][38] ), .B(
        \mult_22/CARRYB[40][38] ), .CI(\mult_22/SUMB[40][39] ), .CO(
        \mult_22/CARRYB[41][38] ), .S(\mult_22/SUMB[41][38] ) );
  FA_X1 \mult_22/S2_41_37  ( .A(\mult_22/ab[41][37] ), .B(
        \mult_22/CARRYB[40][37] ), .CI(\mult_22/SUMB[40][38] ), .CO(
        \mult_22/CARRYB[41][37] ), .S(\mult_22/SUMB[41][37] ) );
  FA_X1 \mult_22/S2_41_36  ( .A(\mult_22/ab[41][36] ), .B(
        \mult_22/CARRYB[40][36] ), .CI(\mult_22/SUMB[40][37] ), .CO(
        \mult_22/CARRYB[41][36] ), .S(\mult_22/SUMB[41][36] ) );
  FA_X1 \mult_22/S2_41_35  ( .A(\mult_22/ab[41][35] ), .B(
        \mult_22/CARRYB[40][35] ), .CI(\mult_22/SUMB[40][36] ), .CO(
        \mult_22/CARRYB[41][35] ), .S(\mult_22/SUMB[41][35] ) );
  FA_X1 \mult_22/S2_41_34  ( .A(\mult_22/ab[41][34] ), .B(
        \mult_22/CARRYB[40][34] ), .CI(\mult_22/SUMB[40][35] ), .CO(
        \mult_22/CARRYB[41][34] ), .S(\mult_22/SUMB[41][34] ) );
  FA_X1 \mult_22/S2_41_33  ( .A(\mult_22/ab[41][33] ), .B(
        \mult_22/CARRYB[40][33] ), .CI(\mult_22/SUMB[40][34] ), .CO(
        \mult_22/CARRYB[41][33] ), .S(\mult_22/SUMB[41][33] ) );
  FA_X1 \mult_22/S2_41_32  ( .A(\mult_22/ab[41][32] ), .B(
        \mult_22/CARRYB[40][32] ), .CI(\mult_22/SUMB[40][33] ), .CO(
        \mult_22/CARRYB[41][32] ), .S(\mult_22/SUMB[41][32] ) );
  FA_X1 \mult_22/S2_41_31  ( .A(\mult_22/ab[41][31] ), .B(
        \mult_22/CARRYB[40][31] ), .CI(\mult_22/SUMB[40][32] ), .CO(
        \mult_22/CARRYB[41][31] ), .S(\mult_22/SUMB[41][31] ) );
  FA_X1 \mult_22/S2_41_30  ( .A(\mult_22/ab[41][30] ), .B(
        \mult_22/CARRYB[40][30] ), .CI(\mult_22/SUMB[40][31] ), .CO(
        \mult_22/CARRYB[41][30] ), .S(\mult_22/SUMB[41][30] ) );
  FA_X1 \mult_22/S2_41_29  ( .A(\mult_22/ab[41][29] ), .B(
        \mult_22/CARRYB[40][29] ), .CI(\mult_22/SUMB[40][30] ), .CO(
        \mult_22/CARRYB[41][29] ), .S(\mult_22/SUMB[41][29] ) );
  FA_X1 \mult_22/S2_41_28  ( .A(\mult_22/ab[41][28] ), .B(
        \mult_22/CARRYB[40][28] ), .CI(\mult_22/SUMB[40][29] ), .CO(
        \mult_22/CARRYB[41][28] ), .S(\mult_22/SUMB[41][28] ) );
  FA_X1 \mult_22/S2_41_27  ( .A(\mult_22/ab[41][27] ), .B(
        \mult_22/CARRYB[40][27] ), .CI(\mult_22/SUMB[40][28] ), .CO(
        \mult_22/CARRYB[41][27] ), .S(\mult_22/SUMB[41][27] ) );
  FA_X1 \mult_22/S2_41_26  ( .A(\mult_22/CARRYB[40][26] ), .B(
        \mult_22/ab[41][26] ), .CI(\mult_22/SUMB[40][27] ), .CO(
        \mult_22/CARRYB[41][26] ), .S(\mult_22/SUMB[41][26] ) );
  FA_X1 \mult_22/S2_41_25  ( .A(\mult_22/ab[41][25] ), .B(
        \mult_22/CARRYB[40][25] ), .CI(\mult_22/SUMB[40][26] ), .CO(
        \mult_22/CARRYB[41][25] ), .S(\mult_22/SUMB[41][25] ) );
  FA_X1 \mult_22/S2_41_24  ( .A(\mult_22/ab[41][24] ), .B(
        \mult_22/CARRYB[40][24] ), .CI(\mult_22/SUMB[40][25] ), .CO(
        \mult_22/CARRYB[41][24] ), .S(\mult_22/SUMB[41][24] ) );
  FA_X1 \mult_22/S2_41_23  ( .A(\mult_22/ab[41][23] ), .B(
        \mult_22/CARRYB[40][23] ), .CI(\mult_22/SUMB[40][24] ), .CO(
        \mult_22/CARRYB[41][23] ), .S(\mult_22/SUMB[41][23] ) );
  FA_X1 \mult_22/S2_41_22  ( .A(\mult_22/ab[41][22] ), .B(
        \mult_22/CARRYB[40][22] ), .CI(\mult_22/SUMB[40][23] ), .CO(
        \mult_22/CARRYB[41][22] ), .S(\mult_22/SUMB[41][22] ) );
  FA_X1 \mult_22/S2_41_21  ( .A(\mult_22/ab[41][21] ), .B(
        \mult_22/CARRYB[40][21] ), .CI(\mult_22/SUMB[40][22] ), .CO(
        \mult_22/CARRYB[41][21] ), .S(\mult_22/SUMB[41][21] ) );
  FA_X1 \mult_22/S2_41_20  ( .A(\mult_22/ab[41][20] ), .B(
        \mult_22/CARRYB[40][20] ), .CI(\mult_22/SUMB[40][21] ), .CO(
        \mult_22/CARRYB[41][20] ), .S(\mult_22/SUMB[41][20] ) );
  FA_X1 \mult_22/S2_41_19  ( .A(\mult_22/ab[41][19] ), .B(
        \mult_22/CARRYB[40][19] ), .CI(\mult_22/SUMB[40][20] ), .CO(
        \mult_22/CARRYB[41][19] ), .S(\mult_22/SUMB[41][19] ) );
  FA_X1 \mult_22/S2_41_18  ( .A(\mult_22/ab[41][18] ), .B(
        \mult_22/CARRYB[40][18] ), .CI(\mult_22/SUMB[40][19] ), .CO(
        \mult_22/CARRYB[41][18] ), .S(\mult_22/SUMB[41][18] ) );
  FA_X1 \mult_22/S2_41_17  ( .A(\mult_22/ab[41][17] ), .B(
        \mult_22/CARRYB[40][17] ), .CI(\mult_22/SUMB[40][18] ), .CO(
        \mult_22/CARRYB[41][17] ), .S(\mult_22/SUMB[41][17] ) );
  FA_X1 \mult_22/S2_41_16  ( .A(\mult_22/ab[41][16] ), .B(
        \mult_22/CARRYB[40][16] ), .CI(\mult_22/SUMB[40][17] ), .CO(
        \mult_22/CARRYB[41][16] ), .S(\mult_22/SUMB[41][16] ) );
  FA_X1 \mult_22/S2_41_15  ( .A(\mult_22/ab[41][15] ), .B(
        \mult_22/CARRYB[40][15] ), .CI(\mult_22/SUMB[40][16] ), .CO(
        \mult_22/CARRYB[41][15] ), .S(\mult_22/SUMB[41][15] ) );
  FA_X1 \mult_22/S2_41_14  ( .A(\mult_22/ab[41][14] ), .B(
        \mult_22/CARRYB[40][14] ), .CI(\mult_22/SUMB[40][15] ), .CO(
        \mult_22/CARRYB[41][14] ), .S(\mult_22/SUMB[41][14] ) );
  FA_X1 \mult_22/S2_41_13  ( .A(\mult_22/ab[41][13] ), .B(
        \mult_22/CARRYB[40][13] ), .CI(\mult_22/SUMB[40][14] ), .CO(
        \mult_22/CARRYB[41][13] ), .S(\mult_22/SUMB[41][13] ) );
  FA_X1 \mult_22/S2_41_12  ( .A(\mult_22/ab[41][12] ), .B(
        \mult_22/CARRYB[40][12] ), .CI(\mult_22/SUMB[40][13] ), .CO(
        \mult_22/CARRYB[41][12] ), .S(\mult_22/SUMB[41][12] ) );
  FA_X1 \mult_22/S2_41_11  ( .A(\mult_22/ab[41][11] ), .B(
        \mult_22/CARRYB[40][11] ), .CI(\mult_22/SUMB[40][12] ), .CO(
        \mult_22/CARRYB[41][11] ), .S(\mult_22/SUMB[41][11] ) );
  FA_X1 \mult_22/S2_41_10  ( .A(\mult_22/ab[41][10] ), .B(
        \mult_22/CARRYB[40][10] ), .CI(\mult_22/SUMB[40][11] ), .CO(
        \mult_22/CARRYB[41][10] ), .S(\mult_22/SUMB[41][10] ) );
  FA_X1 \mult_22/S2_41_9  ( .A(\mult_22/ab[41][9] ), .B(
        \mult_22/CARRYB[40][9] ), .CI(\mult_22/SUMB[40][10] ), .CO(
        \mult_22/CARRYB[41][9] ), .S(\mult_22/SUMB[41][9] ) );
  FA_X1 \mult_22/S2_41_8  ( .A(\mult_22/ab[41][8] ), .B(
        \mult_22/CARRYB[40][8] ), .CI(\mult_22/SUMB[40][9] ), .CO(
        \mult_22/CARRYB[41][8] ), .S(\mult_22/SUMB[41][8] ) );
  FA_X1 \mult_22/S2_41_7  ( .A(\mult_22/ab[41][7] ), .B(
        \mult_22/CARRYB[40][7] ), .CI(\mult_22/SUMB[40][8] ), .CO(
        \mult_22/CARRYB[41][7] ), .S(\mult_22/SUMB[41][7] ) );
  FA_X1 \mult_22/S2_41_6  ( .A(\mult_22/ab[41][6] ), .B(
        \mult_22/CARRYB[40][6] ), .CI(\mult_22/SUMB[40][7] ), .CO(
        \mult_22/CARRYB[41][6] ), .S(\mult_22/SUMB[41][6] ) );
  FA_X1 \mult_22/S2_41_5  ( .A(\mult_22/ab[41][5] ), .B(
        \mult_22/CARRYB[40][5] ), .CI(\mult_22/SUMB[40][6] ), .CO(
        \mult_22/CARRYB[41][5] ), .S(\mult_22/SUMB[41][5] ) );
  FA_X1 \mult_22/S2_41_4  ( .A(\mult_22/ab[41][4] ), .B(
        \mult_22/CARRYB[40][4] ), .CI(\mult_22/SUMB[40][5] ), .CO(
        \mult_22/CARRYB[41][4] ), .S(\mult_22/SUMB[41][4] ) );
  FA_X1 \mult_22/S2_41_3  ( .A(\mult_22/ab[41][3] ), .B(
        \mult_22/CARRYB[40][3] ), .CI(\mult_22/SUMB[40][4] ), .CO(
        \mult_22/CARRYB[41][3] ), .S(\mult_22/SUMB[41][3] ) );
  FA_X1 \mult_22/S2_41_2  ( .A(\mult_22/ab[41][2] ), .B(
        \mult_22/CARRYB[40][2] ), .CI(\mult_22/SUMB[40][3] ), .CO(
        \mult_22/CARRYB[41][2] ), .S(\mult_22/SUMB[41][2] ) );
  FA_X1 \mult_22/S2_41_1  ( .A(\mult_22/ab[41][1] ), .B(
        \mult_22/CARRYB[40][1] ), .CI(\mult_22/SUMB[40][2] ), .CO(
        \mult_22/CARRYB[41][1] ), .S(\mult_22/SUMB[41][1] ) );
  FA_X1 \mult_22/S1_41_0  ( .A(\mult_22/ab[41][0] ), .B(
        \mult_22/CARRYB[40][0] ), .CI(\mult_22/SUMB[40][1] ), .CO(
        \mult_22/CARRYB[41][0] ), .S(N169) );
  FA_X1 \mult_22/S3_42_62  ( .A(\mult_22/ab[42][62] ), .B(
        \mult_22/CARRYB[41][62] ), .CI(\mult_22/ab[41][63] ), .CO(
        \mult_22/CARRYB[42][62] ), .S(\mult_22/SUMB[42][62] ) );
  FA_X1 \mult_22/S2_42_61  ( .A(\mult_22/ab[42][61] ), .B(
        \mult_22/CARRYB[41][61] ), .CI(\mult_22/SUMB[41][62] ), .CO(
        \mult_22/CARRYB[42][61] ), .S(\mult_22/SUMB[42][61] ) );
  FA_X1 \mult_22/S2_42_60  ( .A(\mult_22/ab[42][60] ), .B(
        \mult_22/CARRYB[41][60] ), .CI(\mult_22/SUMB[41][61] ), .CO(
        \mult_22/CARRYB[42][60] ), .S(\mult_22/SUMB[42][60] ) );
  FA_X1 \mult_22/S2_42_59  ( .A(\mult_22/ab[42][59] ), .B(
        \mult_22/CARRYB[41][59] ), .CI(\mult_22/SUMB[41][60] ), .CO(
        \mult_22/CARRYB[42][59] ), .S(\mult_22/SUMB[42][59] ) );
  FA_X1 \mult_22/S2_42_58  ( .A(\mult_22/ab[42][58] ), .B(
        \mult_22/CARRYB[41][58] ), .CI(\mult_22/SUMB[41][59] ), .CO(
        \mult_22/CARRYB[42][58] ), .S(\mult_22/SUMB[42][58] ) );
  FA_X1 \mult_22/S2_42_57  ( .A(\mult_22/ab[42][57] ), .B(
        \mult_22/CARRYB[41][57] ), .CI(\mult_22/SUMB[41][58] ), .CO(
        \mult_22/CARRYB[42][57] ), .S(\mult_22/SUMB[42][57] ) );
  FA_X1 \mult_22/S2_42_56  ( .A(\mult_22/ab[42][56] ), .B(
        \mult_22/CARRYB[41][56] ), .CI(\mult_22/SUMB[41][57] ), .CO(
        \mult_22/CARRYB[42][56] ), .S(\mult_22/SUMB[42][56] ) );
  FA_X1 \mult_22/S2_42_55  ( .A(\mult_22/ab[42][55] ), .B(
        \mult_22/CARRYB[41][55] ), .CI(\mult_22/SUMB[41][56] ), .CO(
        \mult_22/CARRYB[42][55] ), .S(\mult_22/SUMB[42][55] ) );
  FA_X1 \mult_22/S2_42_54  ( .A(\mult_22/ab[42][54] ), .B(
        \mult_22/CARRYB[41][54] ), .CI(\mult_22/SUMB[41][55] ), .CO(
        \mult_22/CARRYB[42][54] ), .S(\mult_22/SUMB[42][54] ) );
  FA_X1 \mult_22/S2_42_53  ( .A(\mult_22/ab[42][53] ), .B(
        \mult_22/CARRYB[41][53] ), .CI(\mult_22/SUMB[41][54] ), .CO(
        \mult_22/CARRYB[42][53] ), .S(\mult_22/SUMB[42][53] ) );
  FA_X1 \mult_22/S2_42_52  ( .A(\mult_22/ab[42][52] ), .B(
        \mult_22/CARRYB[41][52] ), .CI(\mult_22/SUMB[41][53] ), .CO(
        \mult_22/CARRYB[42][52] ), .S(\mult_22/SUMB[42][52] ) );
  FA_X1 \mult_22/S2_42_51  ( .A(\mult_22/ab[42][51] ), .B(
        \mult_22/CARRYB[41][51] ), .CI(\mult_22/SUMB[41][52] ), .CO(
        \mult_22/CARRYB[42][51] ), .S(\mult_22/SUMB[42][51] ) );
  FA_X1 \mult_22/S2_42_50  ( .A(\mult_22/ab[42][50] ), .B(
        \mult_22/CARRYB[41][50] ), .CI(\mult_22/SUMB[41][51] ), .CO(
        \mult_22/CARRYB[42][50] ), .S(\mult_22/SUMB[42][50] ) );
  FA_X1 \mult_22/S2_42_49  ( .A(\mult_22/ab[42][49] ), .B(
        \mult_22/CARRYB[41][49] ), .CI(\mult_22/SUMB[41][50] ), .CO(
        \mult_22/CARRYB[42][49] ), .S(\mult_22/SUMB[42][49] ) );
  FA_X1 \mult_22/S2_42_48  ( .A(\mult_22/ab[42][48] ), .B(
        \mult_22/CARRYB[41][48] ), .CI(\mult_22/SUMB[41][49] ), .CO(
        \mult_22/CARRYB[42][48] ), .S(\mult_22/SUMB[42][48] ) );
  FA_X1 \mult_22/S2_42_47  ( .A(\mult_22/ab[42][47] ), .B(
        \mult_22/CARRYB[41][47] ), .CI(\mult_22/SUMB[41][48] ), .CO(
        \mult_22/CARRYB[42][47] ), .S(\mult_22/SUMB[42][47] ) );
  FA_X1 \mult_22/S2_42_46  ( .A(\mult_22/ab[42][46] ), .B(
        \mult_22/CARRYB[41][46] ), .CI(\mult_22/SUMB[41][47] ), .CO(
        \mult_22/CARRYB[42][46] ), .S(\mult_22/SUMB[42][46] ) );
  FA_X1 \mult_22/S2_42_45  ( .A(\mult_22/ab[42][45] ), .B(
        \mult_22/CARRYB[41][45] ), .CI(\mult_22/SUMB[41][46] ), .CO(
        \mult_22/CARRYB[42][45] ), .S(\mult_22/SUMB[42][45] ) );
  FA_X1 \mult_22/S2_42_44  ( .A(\mult_22/ab[42][44] ), .B(
        \mult_22/CARRYB[41][44] ), .CI(\mult_22/SUMB[41][45] ), .CO(
        \mult_22/CARRYB[42][44] ), .S(\mult_22/SUMB[42][44] ) );
  FA_X1 \mult_22/S2_42_43  ( .A(\mult_22/ab[42][43] ), .B(
        \mult_22/CARRYB[41][43] ), .CI(\mult_22/SUMB[41][44] ), .CO(
        \mult_22/CARRYB[42][43] ), .S(\mult_22/SUMB[42][43] ) );
  FA_X1 \mult_22/S2_42_42  ( .A(\mult_22/ab[42][42] ), .B(
        \mult_22/CARRYB[41][42] ), .CI(\mult_22/SUMB[41][43] ), .CO(
        \mult_22/CARRYB[42][42] ), .S(\mult_22/SUMB[42][42] ) );
  FA_X1 \mult_22/S2_42_41  ( .A(\mult_22/ab[42][41] ), .B(
        \mult_22/CARRYB[41][41] ), .CI(\mult_22/SUMB[41][42] ), .CO(
        \mult_22/CARRYB[42][41] ), .S(\mult_22/SUMB[42][41] ) );
  FA_X1 \mult_22/S2_42_40  ( .A(\mult_22/ab[42][40] ), .B(
        \mult_22/CARRYB[41][40] ), .CI(\mult_22/SUMB[41][41] ), .CO(
        \mult_22/CARRYB[42][40] ), .S(\mult_22/SUMB[42][40] ) );
  FA_X1 \mult_22/S2_42_39  ( .A(\mult_22/ab[42][39] ), .B(
        \mult_22/CARRYB[41][39] ), .CI(\mult_22/SUMB[41][40] ), .CO(
        \mult_22/CARRYB[42][39] ), .S(\mult_22/SUMB[42][39] ) );
  FA_X1 \mult_22/S2_42_38  ( .A(\mult_22/ab[42][38] ), .B(
        \mult_22/CARRYB[41][38] ), .CI(\mult_22/SUMB[41][39] ), .CO(
        \mult_22/CARRYB[42][38] ), .S(\mult_22/SUMB[42][38] ) );
  FA_X1 \mult_22/S2_42_37  ( .A(\mult_22/ab[42][37] ), .B(
        \mult_22/CARRYB[41][37] ), .CI(\mult_22/SUMB[41][38] ), .CO(
        \mult_22/CARRYB[42][37] ), .S(\mult_22/SUMB[42][37] ) );
  FA_X1 \mult_22/S2_42_36  ( .A(\mult_22/ab[42][36] ), .B(
        \mult_22/CARRYB[41][36] ), .CI(\mult_22/SUMB[41][37] ), .CO(
        \mult_22/CARRYB[42][36] ), .S(\mult_22/SUMB[42][36] ) );
  FA_X1 \mult_22/S2_42_35  ( .A(\mult_22/ab[42][35] ), .B(
        \mult_22/CARRYB[41][35] ), .CI(\mult_22/SUMB[41][36] ), .CO(
        \mult_22/CARRYB[42][35] ), .S(\mult_22/SUMB[42][35] ) );
  FA_X1 \mult_22/S2_42_34  ( .A(\mult_22/ab[42][34] ), .B(
        \mult_22/CARRYB[41][34] ), .CI(\mult_22/SUMB[41][35] ), .CO(
        \mult_22/CARRYB[42][34] ), .S(\mult_22/SUMB[42][34] ) );
  FA_X1 \mult_22/S2_42_33  ( .A(\mult_22/ab[42][33] ), .B(
        \mult_22/CARRYB[41][33] ), .CI(\mult_22/SUMB[41][34] ), .CO(
        \mult_22/CARRYB[42][33] ), .S(\mult_22/SUMB[42][33] ) );
  FA_X1 \mult_22/S2_42_32  ( .A(\mult_22/ab[42][32] ), .B(
        \mult_22/CARRYB[41][32] ), .CI(\mult_22/SUMB[41][33] ), .CO(
        \mult_22/CARRYB[42][32] ), .S(\mult_22/SUMB[42][32] ) );
  FA_X1 \mult_22/S2_42_31  ( .A(\mult_22/ab[42][31] ), .B(
        \mult_22/CARRYB[41][31] ), .CI(\mult_22/SUMB[41][32] ), .CO(
        \mult_22/CARRYB[42][31] ), .S(\mult_22/SUMB[42][31] ) );
  FA_X1 \mult_22/S2_42_30  ( .A(\mult_22/ab[42][30] ), .B(
        \mult_22/CARRYB[41][30] ), .CI(\mult_22/SUMB[41][31] ), .CO(
        \mult_22/CARRYB[42][30] ), .S(\mult_22/SUMB[42][30] ) );
  FA_X1 \mult_22/S2_42_29  ( .A(\mult_22/ab[42][29] ), .B(
        \mult_22/CARRYB[41][29] ), .CI(\mult_22/SUMB[41][30] ), .CO(
        \mult_22/CARRYB[42][29] ), .S(\mult_22/SUMB[42][29] ) );
  FA_X1 \mult_22/S2_42_28  ( .A(\mult_22/ab[42][28] ), .B(
        \mult_22/CARRYB[41][28] ), .CI(\mult_22/SUMB[41][29] ), .CO(
        \mult_22/CARRYB[42][28] ), .S(\mult_22/SUMB[42][28] ) );
  FA_X1 \mult_22/S2_42_27  ( .A(\mult_22/ab[42][27] ), .B(
        \mult_22/CARRYB[41][27] ), .CI(\mult_22/SUMB[41][28] ), .CO(
        \mult_22/CARRYB[42][27] ), .S(\mult_22/SUMB[42][27] ) );
  FA_X1 \mult_22/S2_42_26  ( .A(\mult_22/ab[42][26] ), .B(
        \mult_22/CARRYB[41][26] ), .CI(\mult_22/SUMB[41][27] ), .CO(
        \mult_22/CARRYB[42][26] ), .S(\mult_22/SUMB[42][26] ) );
  FA_X1 \mult_22/S2_42_25  ( .A(\mult_22/ab[42][25] ), .B(
        \mult_22/CARRYB[41][25] ), .CI(\mult_22/SUMB[41][26] ), .CO(
        \mult_22/CARRYB[42][25] ), .S(\mult_22/SUMB[42][25] ) );
  FA_X1 \mult_22/S2_42_24  ( .A(\mult_22/ab[42][24] ), .B(
        \mult_22/CARRYB[41][24] ), .CI(\mult_22/SUMB[41][25] ), .CO(
        \mult_22/CARRYB[42][24] ), .S(\mult_22/SUMB[42][24] ) );
  FA_X1 \mult_22/S2_42_23  ( .A(\mult_22/ab[42][23] ), .B(
        \mult_22/CARRYB[41][23] ), .CI(\mult_22/SUMB[41][24] ), .CO(
        \mult_22/CARRYB[42][23] ), .S(\mult_22/SUMB[42][23] ) );
  FA_X1 \mult_22/S2_42_22  ( .A(\mult_22/CARRYB[41][22] ), .B(
        \mult_22/ab[42][22] ), .CI(\mult_22/SUMB[41][23] ), .CO(
        \mult_22/CARRYB[42][22] ), .S(\mult_22/SUMB[42][22] ) );
  FA_X1 \mult_22/S2_42_21  ( .A(\mult_22/ab[42][21] ), .B(
        \mult_22/CARRYB[41][21] ), .CI(\mult_22/SUMB[41][22] ), .CO(
        \mult_22/CARRYB[42][21] ), .S(\mult_22/SUMB[42][21] ) );
  FA_X1 \mult_22/S2_42_20  ( .A(\mult_22/ab[42][20] ), .B(
        \mult_22/CARRYB[41][20] ), .CI(\mult_22/SUMB[41][21] ), .CO(
        \mult_22/CARRYB[42][20] ), .S(\mult_22/SUMB[42][20] ) );
  FA_X1 \mult_22/S2_42_19  ( .A(\mult_22/ab[42][19] ), .B(
        \mult_22/CARRYB[41][19] ), .CI(\mult_22/SUMB[41][20] ), .CO(
        \mult_22/CARRYB[42][19] ), .S(\mult_22/SUMB[42][19] ) );
  FA_X1 \mult_22/S2_42_18  ( .A(\mult_22/ab[42][18] ), .B(
        \mult_22/CARRYB[41][18] ), .CI(\mult_22/SUMB[41][19] ), .CO(
        \mult_22/CARRYB[42][18] ), .S(\mult_22/SUMB[42][18] ) );
  FA_X1 \mult_22/S2_42_17  ( .A(\mult_22/ab[42][17] ), .B(
        \mult_22/CARRYB[41][17] ), .CI(\mult_22/SUMB[41][18] ), .CO(
        \mult_22/CARRYB[42][17] ), .S(\mult_22/SUMB[42][17] ) );
  FA_X1 \mult_22/S2_42_16  ( .A(\mult_22/ab[42][16] ), .B(
        \mult_22/CARRYB[41][16] ), .CI(\mult_22/SUMB[41][17] ), .CO(
        \mult_22/CARRYB[42][16] ), .S(\mult_22/SUMB[42][16] ) );
  FA_X1 \mult_22/S2_42_15  ( .A(\mult_22/ab[42][15] ), .B(
        \mult_22/CARRYB[41][15] ), .CI(\mult_22/SUMB[41][16] ), .CO(
        \mult_22/CARRYB[42][15] ), .S(\mult_22/SUMB[42][15] ) );
  FA_X1 \mult_22/S2_42_14  ( .A(\mult_22/ab[42][14] ), .B(
        \mult_22/CARRYB[41][14] ), .CI(\mult_22/SUMB[41][15] ), .CO(
        \mult_22/CARRYB[42][14] ), .S(\mult_22/SUMB[42][14] ) );
  FA_X1 \mult_22/S2_42_13  ( .A(\mult_22/ab[42][13] ), .B(
        \mult_22/CARRYB[41][13] ), .CI(\mult_22/SUMB[41][14] ), .CO(
        \mult_22/CARRYB[42][13] ), .S(\mult_22/SUMB[42][13] ) );
  FA_X1 \mult_22/S2_42_12  ( .A(\mult_22/ab[42][12] ), .B(
        \mult_22/CARRYB[41][12] ), .CI(\mult_22/SUMB[41][13] ), .CO(
        \mult_22/CARRYB[42][12] ), .S(\mult_22/SUMB[42][12] ) );
  FA_X1 \mult_22/S2_42_11  ( .A(\mult_22/ab[42][11] ), .B(
        \mult_22/CARRYB[41][11] ), .CI(\mult_22/SUMB[41][12] ), .CO(
        \mult_22/CARRYB[42][11] ), .S(\mult_22/SUMB[42][11] ) );
  FA_X1 \mult_22/S2_42_10  ( .A(\mult_22/ab[42][10] ), .B(
        \mult_22/CARRYB[41][10] ), .CI(\mult_22/SUMB[41][11] ), .CO(
        \mult_22/CARRYB[42][10] ), .S(\mult_22/SUMB[42][10] ) );
  FA_X1 \mult_22/S2_42_9  ( .A(\mult_22/ab[42][9] ), .B(
        \mult_22/CARRYB[41][9] ), .CI(\mult_22/SUMB[41][10] ), .CO(
        \mult_22/CARRYB[42][9] ), .S(\mult_22/SUMB[42][9] ) );
  FA_X1 \mult_22/S2_42_8  ( .A(\mult_22/ab[42][8] ), .B(
        \mult_22/CARRYB[41][8] ), .CI(\mult_22/SUMB[41][9] ), .CO(
        \mult_22/CARRYB[42][8] ), .S(\mult_22/SUMB[42][8] ) );
  FA_X1 \mult_22/S2_42_7  ( .A(\mult_22/ab[42][7] ), .B(
        \mult_22/CARRYB[41][7] ), .CI(\mult_22/SUMB[41][8] ), .CO(
        \mult_22/CARRYB[42][7] ), .S(\mult_22/SUMB[42][7] ) );
  FA_X1 \mult_22/S2_42_6  ( .A(\mult_22/ab[42][6] ), .B(
        \mult_22/CARRYB[41][6] ), .CI(\mult_22/SUMB[41][7] ), .CO(
        \mult_22/CARRYB[42][6] ), .S(\mult_22/SUMB[42][6] ) );
  FA_X1 \mult_22/S2_42_5  ( .A(\mult_22/ab[42][5] ), .B(
        \mult_22/CARRYB[41][5] ), .CI(\mult_22/SUMB[41][6] ), .CO(
        \mult_22/CARRYB[42][5] ), .S(\mult_22/SUMB[42][5] ) );
  FA_X1 \mult_22/S2_42_4  ( .A(\mult_22/ab[42][4] ), .B(
        \mult_22/CARRYB[41][4] ), .CI(\mult_22/SUMB[41][5] ), .CO(
        \mult_22/CARRYB[42][4] ), .S(\mult_22/SUMB[42][4] ) );
  FA_X1 \mult_22/S2_42_3  ( .A(\mult_22/ab[42][3] ), .B(
        \mult_22/CARRYB[41][3] ), .CI(\mult_22/SUMB[41][4] ), .CO(
        \mult_22/CARRYB[42][3] ), .S(\mult_22/SUMB[42][3] ) );
  FA_X1 \mult_22/S2_42_2  ( .A(\mult_22/ab[42][2] ), .B(
        \mult_22/CARRYB[41][2] ), .CI(\mult_22/SUMB[41][3] ), .CO(
        \mult_22/CARRYB[42][2] ), .S(\mult_22/SUMB[42][2] ) );
  FA_X1 \mult_22/S2_42_1  ( .A(\mult_22/ab[42][1] ), .B(
        \mult_22/CARRYB[41][1] ), .CI(\mult_22/SUMB[41][2] ), .CO(
        \mult_22/CARRYB[42][1] ), .S(\mult_22/SUMB[42][1] ) );
  FA_X1 \mult_22/S1_42_0  ( .A(\mult_22/ab[42][0] ), .B(
        \mult_22/CARRYB[41][0] ), .CI(\mult_22/SUMB[41][1] ), .CO(
        \mult_22/CARRYB[42][0] ), .S(N170) );
  FA_X1 \mult_22/S3_43_62  ( .A(\mult_22/ab[43][62] ), .B(
        \mult_22/CARRYB[42][62] ), .CI(\mult_22/ab[42][63] ), .CO(
        \mult_22/CARRYB[43][62] ), .S(\mult_22/SUMB[43][62] ) );
  FA_X1 \mult_22/S2_43_61  ( .A(\mult_22/ab[43][61] ), .B(
        \mult_22/CARRYB[42][61] ), .CI(\mult_22/SUMB[42][62] ), .CO(
        \mult_22/CARRYB[43][61] ), .S(\mult_22/SUMB[43][61] ) );
  FA_X1 \mult_22/S2_43_60  ( .A(\mult_22/ab[43][60] ), .B(
        \mult_22/CARRYB[42][60] ), .CI(\mult_22/SUMB[42][61] ), .CO(
        \mult_22/CARRYB[43][60] ), .S(\mult_22/SUMB[43][60] ) );
  FA_X1 \mult_22/S2_43_59  ( .A(\mult_22/ab[43][59] ), .B(
        \mult_22/CARRYB[42][59] ), .CI(\mult_22/SUMB[42][60] ), .CO(
        \mult_22/CARRYB[43][59] ), .S(\mult_22/SUMB[43][59] ) );
  FA_X1 \mult_22/S2_43_58  ( .A(\mult_22/ab[43][58] ), .B(
        \mult_22/CARRYB[42][58] ), .CI(\mult_22/SUMB[42][59] ), .CO(
        \mult_22/CARRYB[43][58] ), .S(\mult_22/SUMB[43][58] ) );
  FA_X1 \mult_22/S2_43_57  ( .A(\mult_22/ab[43][57] ), .B(
        \mult_22/CARRYB[42][57] ), .CI(\mult_22/SUMB[42][58] ), .CO(
        \mult_22/CARRYB[43][57] ), .S(\mult_22/SUMB[43][57] ) );
  FA_X1 \mult_22/S2_43_56  ( .A(\mult_22/ab[43][56] ), .B(
        \mult_22/CARRYB[42][56] ), .CI(\mult_22/SUMB[42][57] ), .CO(
        \mult_22/CARRYB[43][56] ), .S(\mult_22/SUMB[43][56] ) );
  FA_X1 \mult_22/S2_43_55  ( .A(\mult_22/ab[43][55] ), .B(
        \mult_22/CARRYB[42][55] ), .CI(\mult_22/SUMB[42][56] ), .CO(
        \mult_22/CARRYB[43][55] ), .S(\mult_22/SUMB[43][55] ) );
  FA_X1 \mult_22/S2_43_54  ( .A(\mult_22/ab[43][54] ), .B(
        \mult_22/CARRYB[42][54] ), .CI(\mult_22/SUMB[42][55] ), .CO(
        \mult_22/CARRYB[43][54] ), .S(\mult_22/SUMB[43][54] ) );
  FA_X1 \mult_22/S2_43_53  ( .A(\mult_22/ab[43][53] ), .B(
        \mult_22/CARRYB[42][53] ), .CI(\mult_22/SUMB[42][54] ), .CO(
        \mult_22/CARRYB[43][53] ), .S(\mult_22/SUMB[43][53] ) );
  FA_X1 \mult_22/S2_43_52  ( .A(\mult_22/ab[43][52] ), .B(
        \mult_22/CARRYB[42][52] ), .CI(\mult_22/SUMB[42][53] ), .CO(
        \mult_22/CARRYB[43][52] ), .S(\mult_22/SUMB[43][52] ) );
  FA_X1 \mult_22/S2_43_51  ( .A(\mult_22/ab[43][51] ), .B(
        \mult_22/CARRYB[42][51] ), .CI(\mult_22/SUMB[42][52] ), .CO(
        \mult_22/CARRYB[43][51] ), .S(\mult_22/SUMB[43][51] ) );
  FA_X1 \mult_22/S2_43_50  ( .A(\mult_22/ab[43][50] ), .B(
        \mult_22/CARRYB[42][50] ), .CI(\mult_22/SUMB[42][51] ), .CO(
        \mult_22/CARRYB[43][50] ), .S(\mult_22/SUMB[43][50] ) );
  FA_X1 \mult_22/S2_43_49  ( .A(\mult_22/ab[43][49] ), .B(
        \mult_22/CARRYB[42][49] ), .CI(\mult_22/SUMB[42][50] ), .CO(
        \mult_22/CARRYB[43][49] ), .S(\mult_22/SUMB[43][49] ) );
  FA_X1 \mult_22/S2_43_48  ( .A(\mult_22/ab[43][48] ), .B(
        \mult_22/CARRYB[42][48] ), .CI(\mult_22/SUMB[42][49] ), .CO(
        \mult_22/CARRYB[43][48] ), .S(\mult_22/SUMB[43][48] ) );
  FA_X1 \mult_22/S2_43_47  ( .A(\mult_22/ab[43][47] ), .B(
        \mult_22/CARRYB[42][47] ), .CI(\mult_22/SUMB[42][48] ), .CO(
        \mult_22/CARRYB[43][47] ), .S(\mult_22/SUMB[43][47] ) );
  FA_X1 \mult_22/S2_43_46  ( .A(\mult_22/ab[43][46] ), .B(
        \mult_22/CARRYB[42][46] ), .CI(\mult_22/SUMB[42][47] ), .CO(
        \mult_22/CARRYB[43][46] ), .S(\mult_22/SUMB[43][46] ) );
  FA_X1 \mult_22/S2_43_45  ( .A(\mult_22/ab[43][45] ), .B(
        \mult_22/CARRYB[42][45] ), .CI(\mult_22/SUMB[42][46] ), .CO(
        \mult_22/CARRYB[43][45] ), .S(\mult_22/SUMB[43][45] ) );
  FA_X1 \mult_22/S2_43_44  ( .A(\mult_22/ab[43][44] ), .B(
        \mult_22/CARRYB[42][44] ), .CI(\mult_22/SUMB[42][45] ), .CO(
        \mult_22/CARRYB[43][44] ), .S(\mult_22/SUMB[43][44] ) );
  FA_X1 \mult_22/S2_43_43  ( .A(\mult_22/ab[43][43] ), .B(
        \mult_22/CARRYB[42][43] ), .CI(\mult_22/SUMB[42][44] ), .CO(
        \mult_22/CARRYB[43][43] ), .S(\mult_22/SUMB[43][43] ) );
  FA_X1 \mult_22/S2_43_42  ( .A(\mult_22/ab[43][42] ), .B(
        \mult_22/CARRYB[42][42] ), .CI(\mult_22/SUMB[42][43] ), .CO(
        \mult_22/CARRYB[43][42] ), .S(\mult_22/SUMB[43][42] ) );
  FA_X1 \mult_22/S2_43_41  ( .A(\mult_22/ab[43][41] ), .B(
        \mult_22/CARRYB[42][41] ), .CI(\mult_22/SUMB[42][42] ), .CO(
        \mult_22/CARRYB[43][41] ), .S(\mult_22/SUMB[43][41] ) );
  FA_X1 \mult_22/S2_43_40  ( .A(\mult_22/ab[43][40] ), .B(
        \mult_22/CARRYB[42][40] ), .CI(\mult_22/SUMB[42][41] ), .CO(
        \mult_22/CARRYB[43][40] ), .S(\mult_22/SUMB[43][40] ) );
  FA_X1 \mult_22/S2_43_39  ( .A(\mult_22/ab[43][39] ), .B(
        \mult_22/CARRYB[42][39] ), .CI(\mult_22/SUMB[42][40] ), .CO(
        \mult_22/CARRYB[43][39] ), .S(\mult_22/SUMB[43][39] ) );
  FA_X1 \mult_22/S2_43_38  ( .A(\mult_22/ab[43][38] ), .B(
        \mult_22/CARRYB[42][38] ), .CI(\mult_22/SUMB[42][39] ), .CO(
        \mult_22/CARRYB[43][38] ), .S(\mult_22/SUMB[43][38] ) );
  FA_X1 \mult_22/S2_43_37  ( .A(\mult_22/ab[43][37] ), .B(
        \mult_22/CARRYB[42][37] ), .CI(\mult_22/SUMB[42][38] ), .CO(
        \mult_22/CARRYB[43][37] ), .S(\mult_22/SUMB[43][37] ) );
  FA_X1 \mult_22/S2_43_36  ( .A(\mult_22/ab[43][36] ), .B(
        \mult_22/CARRYB[42][36] ), .CI(\mult_22/SUMB[42][37] ), .CO(
        \mult_22/CARRYB[43][36] ), .S(\mult_22/SUMB[43][36] ) );
  FA_X1 \mult_22/S2_43_35  ( .A(\mult_22/ab[43][35] ), .B(
        \mult_22/CARRYB[42][35] ), .CI(\mult_22/SUMB[42][36] ), .CO(
        \mult_22/CARRYB[43][35] ), .S(\mult_22/SUMB[43][35] ) );
  FA_X1 \mult_22/S2_43_34  ( .A(\mult_22/ab[43][34] ), .B(
        \mult_22/CARRYB[42][34] ), .CI(\mult_22/SUMB[42][35] ), .CO(
        \mult_22/CARRYB[43][34] ), .S(\mult_22/SUMB[43][34] ) );
  FA_X1 \mult_22/S2_43_33  ( .A(\mult_22/ab[43][33] ), .B(
        \mult_22/CARRYB[42][33] ), .CI(\mult_22/SUMB[42][34] ), .CO(
        \mult_22/CARRYB[43][33] ), .S(\mult_22/SUMB[43][33] ) );
  FA_X1 \mult_22/S2_43_32  ( .A(\mult_22/ab[43][32] ), .B(
        \mult_22/CARRYB[42][32] ), .CI(\mult_22/SUMB[42][33] ), .CO(
        \mult_22/CARRYB[43][32] ), .S(\mult_22/SUMB[43][32] ) );
  FA_X1 \mult_22/S2_43_31  ( .A(\mult_22/ab[43][31] ), .B(
        \mult_22/CARRYB[42][31] ), .CI(\mult_22/SUMB[42][32] ), .CO(
        \mult_22/CARRYB[43][31] ), .S(\mult_22/SUMB[43][31] ) );
  FA_X1 \mult_22/S2_43_30  ( .A(\mult_22/ab[43][30] ), .B(
        \mult_22/CARRYB[42][30] ), .CI(\mult_22/SUMB[42][31] ), .CO(
        \mult_22/CARRYB[43][30] ), .S(\mult_22/SUMB[43][30] ) );
  FA_X1 \mult_22/S2_43_29  ( .A(\mult_22/ab[43][29] ), .B(
        \mult_22/CARRYB[42][29] ), .CI(\mult_22/SUMB[42][30] ), .CO(
        \mult_22/CARRYB[43][29] ), .S(\mult_22/SUMB[43][29] ) );
  FA_X1 \mult_22/S2_43_28  ( .A(\mult_22/ab[43][28] ), .B(
        \mult_22/CARRYB[42][28] ), .CI(\mult_22/SUMB[42][29] ), .CO(
        \mult_22/CARRYB[43][28] ), .S(\mult_22/SUMB[43][28] ) );
  FA_X1 \mult_22/S2_43_27  ( .A(\mult_22/ab[43][27] ), .B(
        \mult_22/CARRYB[42][27] ), .CI(\mult_22/SUMB[42][28] ), .CO(
        \mult_22/CARRYB[43][27] ), .S(\mult_22/SUMB[43][27] ) );
  FA_X1 \mult_22/S2_43_26  ( .A(\mult_22/ab[43][26] ), .B(
        \mult_22/CARRYB[42][26] ), .CI(\mult_22/SUMB[42][27] ), .CO(
        \mult_22/CARRYB[43][26] ), .S(\mult_22/SUMB[43][26] ) );
  FA_X1 \mult_22/S2_43_25  ( .A(\mult_22/ab[43][25] ), .B(
        \mult_22/CARRYB[42][25] ), .CI(\mult_22/SUMB[42][26] ), .CO(
        \mult_22/CARRYB[43][25] ), .S(\mult_22/SUMB[43][25] ) );
  FA_X1 \mult_22/S2_43_24  ( .A(\mult_22/CARRYB[42][24] ), .B(
        \mult_22/ab[43][24] ), .CI(\mult_22/SUMB[42][25] ), .CO(
        \mult_22/CARRYB[43][24] ), .S(\mult_22/SUMB[43][24] ) );
  FA_X1 \mult_22/S2_43_23  ( .A(\mult_22/ab[43][23] ), .B(
        \mult_22/CARRYB[42][23] ), .CI(\mult_22/SUMB[42][24] ), .CO(
        \mult_22/CARRYB[43][23] ), .S(\mult_22/SUMB[43][23] ) );
  FA_X1 \mult_22/S2_43_22  ( .A(\mult_22/ab[43][22] ), .B(
        \mult_22/CARRYB[42][22] ), .CI(\mult_22/SUMB[42][23] ), .CO(
        \mult_22/CARRYB[43][22] ), .S(\mult_22/SUMB[43][22] ) );
  FA_X1 \mult_22/S2_43_21  ( .A(\mult_22/ab[43][21] ), .B(
        \mult_22/CARRYB[42][21] ), .CI(\mult_22/SUMB[42][22] ), .CO(
        \mult_22/CARRYB[43][21] ), .S(\mult_22/SUMB[43][21] ) );
  FA_X1 \mult_22/S2_43_20  ( .A(\mult_22/ab[43][20] ), .B(
        \mult_22/CARRYB[42][20] ), .CI(\mult_22/SUMB[42][21] ), .CO(
        \mult_22/CARRYB[43][20] ), .S(\mult_22/SUMB[43][20] ) );
  FA_X1 \mult_22/S2_43_19  ( .A(\mult_22/ab[43][19] ), .B(
        \mult_22/CARRYB[42][19] ), .CI(\mult_22/SUMB[42][20] ), .CO(
        \mult_22/CARRYB[43][19] ), .S(\mult_22/SUMB[43][19] ) );
  FA_X1 \mult_22/S2_43_18  ( .A(\mult_22/ab[43][18] ), .B(
        \mult_22/CARRYB[42][18] ), .CI(\mult_22/SUMB[42][19] ), .CO(
        \mult_22/CARRYB[43][18] ), .S(\mult_22/SUMB[43][18] ) );
  FA_X1 \mult_22/S2_43_17  ( .A(\mult_22/ab[43][17] ), .B(
        \mult_22/CARRYB[42][17] ), .CI(\mult_22/SUMB[42][18] ), .CO(
        \mult_22/CARRYB[43][17] ), .S(\mult_22/SUMB[43][17] ) );
  FA_X1 \mult_22/S2_43_16  ( .A(\mult_22/ab[43][16] ), .B(
        \mult_22/CARRYB[42][16] ), .CI(\mult_22/SUMB[42][17] ), .CO(
        \mult_22/CARRYB[43][16] ), .S(\mult_22/SUMB[43][16] ) );
  FA_X1 \mult_22/S2_43_15  ( .A(\mult_22/ab[43][15] ), .B(
        \mult_22/CARRYB[42][15] ), .CI(\mult_22/SUMB[42][16] ), .CO(
        \mult_22/CARRYB[43][15] ), .S(\mult_22/SUMB[43][15] ) );
  FA_X1 \mult_22/S2_43_14  ( .A(\mult_22/ab[43][14] ), .B(
        \mult_22/CARRYB[42][14] ), .CI(\mult_22/SUMB[42][15] ), .CO(
        \mult_22/CARRYB[43][14] ), .S(\mult_22/SUMB[43][14] ) );
  FA_X1 \mult_22/S2_43_13  ( .A(\mult_22/ab[43][13] ), .B(
        \mult_22/CARRYB[42][13] ), .CI(\mult_22/SUMB[42][14] ), .CO(
        \mult_22/CARRYB[43][13] ), .S(\mult_22/SUMB[43][13] ) );
  FA_X1 \mult_22/S2_43_12  ( .A(\mult_22/ab[43][12] ), .B(
        \mult_22/CARRYB[42][12] ), .CI(\mult_22/SUMB[42][13] ), .CO(
        \mult_22/CARRYB[43][12] ), .S(\mult_22/SUMB[43][12] ) );
  FA_X1 \mult_22/S2_43_11  ( .A(\mult_22/ab[43][11] ), .B(
        \mult_22/CARRYB[42][11] ), .CI(\mult_22/SUMB[42][12] ), .CO(
        \mult_22/CARRYB[43][11] ), .S(\mult_22/SUMB[43][11] ) );
  FA_X1 \mult_22/S2_43_10  ( .A(\mult_22/ab[43][10] ), .B(
        \mult_22/CARRYB[42][10] ), .CI(\mult_22/SUMB[42][11] ), .CO(
        \mult_22/CARRYB[43][10] ), .S(\mult_22/SUMB[43][10] ) );
  FA_X1 \mult_22/S2_43_9  ( .A(\mult_22/ab[43][9] ), .B(
        \mult_22/CARRYB[42][9] ), .CI(\mult_22/SUMB[42][10] ), .CO(
        \mult_22/CARRYB[43][9] ), .S(\mult_22/SUMB[43][9] ) );
  FA_X1 \mult_22/S2_43_8  ( .A(\mult_22/ab[43][8] ), .B(
        \mult_22/CARRYB[42][8] ), .CI(\mult_22/SUMB[42][9] ), .CO(
        \mult_22/CARRYB[43][8] ), .S(\mult_22/SUMB[43][8] ) );
  FA_X1 \mult_22/S2_43_7  ( .A(\mult_22/ab[43][7] ), .B(
        \mult_22/CARRYB[42][7] ), .CI(\mult_22/SUMB[42][8] ), .CO(
        \mult_22/CARRYB[43][7] ), .S(\mult_22/SUMB[43][7] ) );
  FA_X1 \mult_22/S2_43_6  ( .A(\mult_22/ab[43][6] ), .B(
        \mult_22/CARRYB[42][6] ), .CI(\mult_22/SUMB[42][7] ), .CO(
        \mult_22/CARRYB[43][6] ), .S(\mult_22/SUMB[43][6] ) );
  FA_X1 \mult_22/S2_43_5  ( .A(\mult_22/ab[43][5] ), .B(
        \mult_22/CARRYB[42][5] ), .CI(\mult_22/SUMB[42][6] ), .CO(
        \mult_22/CARRYB[43][5] ), .S(\mult_22/SUMB[43][5] ) );
  FA_X1 \mult_22/S2_43_4  ( .A(\mult_22/ab[43][4] ), .B(
        \mult_22/CARRYB[42][4] ), .CI(\mult_22/SUMB[42][5] ), .CO(
        \mult_22/CARRYB[43][4] ), .S(\mult_22/SUMB[43][4] ) );
  FA_X1 \mult_22/S2_43_3  ( .A(\mult_22/ab[43][3] ), .B(
        \mult_22/CARRYB[42][3] ), .CI(\mult_22/SUMB[42][4] ), .CO(
        \mult_22/CARRYB[43][3] ), .S(\mult_22/SUMB[43][3] ) );
  FA_X1 \mult_22/S2_43_2  ( .A(\mult_22/ab[43][2] ), .B(
        \mult_22/CARRYB[42][2] ), .CI(\mult_22/SUMB[42][3] ), .CO(
        \mult_22/CARRYB[43][2] ), .S(\mult_22/SUMB[43][2] ) );
  FA_X1 \mult_22/S2_43_1  ( .A(\mult_22/ab[43][1] ), .B(
        \mult_22/CARRYB[42][1] ), .CI(\mult_22/SUMB[42][2] ), .CO(
        \mult_22/CARRYB[43][1] ), .S(\mult_22/SUMB[43][1] ) );
  FA_X1 \mult_22/S1_43_0  ( .A(\mult_22/ab[43][0] ), .B(
        \mult_22/CARRYB[42][0] ), .CI(\mult_22/SUMB[42][1] ), .CO(
        \mult_22/CARRYB[43][0] ), .S(N171) );
  FA_X1 \mult_22/S3_44_62  ( .A(\mult_22/ab[44][62] ), .B(
        \mult_22/CARRYB[43][62] ), .CI(\mult_22/ab[43][63] ), .CO(
        \mult_22/CARRYB[44][62] ), .S(\mult_22/SUMB[44][62] ) );
  FA_X1 \mult_22/S2_44_61  ( .A(\mult_22/ab[44][61] ), .B(
        \mult_22/CARRYB[43][61] ), .CI(\mult_22/SUMB[43][62] ), .CO(
        \mult_22/CARRYB[44][61] ), .S(\mult_22/SUMB[44][61] ) );
  FA_X1 \mult_22/S2_44_60  ( .A(\mult_22/ab[44][60] ), .B(
        \mult_22/CARRYB[43][60] ), .CI(\mult_22/SUMB[43][61] ), .CO(
        \mult_22/CARRYB[44][60] ), .S(\mult_22/SUMB[44][60] ) );
  FA_X1 \mult_22/S2_44_59  ( .A(\mult_22/ab[44][59] ), .B(
        \mult_22/CARRYB[43][59] ), .CI(\mult_22/SUMB[43][60] ), .CO(
        \mult_22/CARRYB[44][59] ), .S(\mult_22/SUMB[44][59] ) );
  FA_X1 \mult_22/S2_44_58  ( .A(\mult_22/ab[44][58] ), .B(
        \mult_22/CARRYB[43][58] ), .CI(\mult_22/SUMB[43][59] ), .CO(
        \mult_22/CARRYB[44][58] ), .S(\mult_22/SUMB[44][58] ) );
  FA_X1 \mult_22/S2_44_57  ( .A(\mult_22/ab[44][57] ), .B(
        \mult_22/CARRYB[43][57] ), .CI(\mult_22/SUMB[43][58] ), .CO(
        \mult_22/CARRYB[44][57] ), .S(\mult_22/SUMB[44][57] ) );
  FA_X1 \mult_22/S2_44_56  ( .A(\mult_22/ab[44][56] ), .B(
        \mult_22/CARRYB[43][56] ), .CI(\mult_22/SUMB[43][57] ), .CO(
        \mult_22/CARRYB[44][56] ), .S(\mult_22/SUMB[44][56] ) );
  FA_X1 \mult_22/S2_44_55  ( .A(\mult_22/ab[44][55] ), .B(
        \mult_22/CARRYB[43][55] ), .CI(\mult_22/SUMB[43][56] ), .CO(
        \mult_22/CARRYB[44][55] ), .S(\mult_22/SUMB[44][55] ) );
  FA_X1 \mult_22/S2_44_54  ( .A(\mult_22/ab[44][54] ), .B(
        \mult_22/CARRYB[43][54] ), .CI(\mult_22/SUMB[43][55] ), .CO(
        \mult_22/CARRYB[44][54] ), .S(\mult_22/SUMB[44][54] ) );
  FA_X1 \mult_22/S2_44_53  ( .A(\mult_22/ab[44][53] ), .B(
        \mult_22/CARRYB[43][53] ), .CI(\mult_22/SUMB[43][54] ), .CO(
        \mult_22/CARRYB[44][53] ), .S(\mult_22/SUMB[44][53] ) );
  FA_X1 \mult_22/S2_44_52  ( .A(\mult_22/ab[44][52] ), .B(
        \mult_22/CARRYB[43][52] ), .CI(\mult_22/SUMB[43][53] ), .CO(
        \mult_22/CARRYB[44][52] ), .S(\mult_22/SUMB[44][52] ) );
  FA_X1 \mult_22/S2_44_51  ( .A(\mult_22/ab[44][51] ), .B(
        \mult_22/CARRYB[43][51] ), .CI(\mult_22/SUMB[43][52] ), .CO(
        \mult_22/CARRYB[44][51] ), .S(\mult_22/SUMB[44][51] ) );
  FA_X1 \mult_22/S2_44_50  ( .A(\mult_22/ab[44][50] ), .B(
        \mult_22/CARRYB[43][50] ), .CI(\mult_22/SUMB[43][51] ), .CO(
        \mult_22/CARRYB[44][50] ), .S(\mult_22/SUMB[44][50] ) );
  FA_X1 \mult_22/S2_44_49  ( .A(\mult_22/ab[44][49] ), .B(
        \mult_22/CARRYB[43][49] ), .CI(\mult_22/SUMB[43][50] ), .CO(
        \mult_22/CARRYB[44][49] ), .S(\mult_22/SUMB[44][49] ) );
  FA_X1 \mult_22/S2_44_48  ( .A(\mult_22/ab[44][48] ), .B(
        \mult_22/CARRYB[43][48] ), .CI(\mult_22/SUMB[43][49] ), .CO(
        \mult_22/CARRYB[44][48] ), .S(\mult_22/SUMB[44][48] ) );
  FA_X1 \mult_22/S2_44_47  ( .A(\mult_22/ab[44][47] ), .B(
        \mult_22/CARRYB[43][47] ), .CI(\mult_22/SUMB[43][48] ), .CO(
        \mult_22/CARRYB[44][47] ), .S(\mult_22/SUMB[44][47] ) );
  FA_X1 \mult_22/S2_44_46  ( .A(\mult_22/ab[44][46] ), .B(
        \mult_22/CARRYB[43][46] ), .CI(\mult_22/SUMB[43][47] ), .CO(
        \mult_22/CARRYB[44][46] ), .S(\mult_22/SUMB[44][46] ) );
  FA_X1 \mult_22/S2_44_45  ( .A(\mult_22/ab[44][45] ), .B(
        \mult_22/CARRYB[43][45] ), .CI(\mult_22/SUMB[43][46] ), .CO(
        \mult_22/CARRYB[44][45] ), .S(\mult_22/SUMB[44][45] ) );
  FA_X1 \mult_22/S2_44_44  ( .A(\mult_22/ab[44][44] ), .B(
        \mult_22/CARRYB[43][44] ), .CI(\mult_22/SUMB[43][45] ), .CO(
        \mult_22/CARRYB[44][44] ), .S(\mult_22/SUMB[44][44] ) );
  FA_X1 \mult_22/S2_44_43  ( .A(\mult_22/ab[44][43] ), .B(
        \mult_22/CARRYB[43][43] ), .CI(\mult_22/SUMB[43][44] ), .CO(
        \mult_22/CARRYB[44][43] ), .S(\mult_22/SUMB[44][43] ) );
  FA_X1 \mult_22/S2_44_42  ( .A(\mult_22/ab[44][42] ), .B(
        \mult_22/CARRYB[43][42] ), .CI(\mult_22/SUMB[43][43] ), .CO(
        \mult_22/CARRYB[44][42] ), .S(\mult_22/SUMB[44][42] ) );
  FA_X1 \mult_22/S2_44_41  ( .A(\mult_22/ab[44][41] ), .B(
        \mult_22/CARRYB[43][41] ), .CI(\mult_22/SUMB[43][42] ), .CO(
        \mult_22/CARRYB[44][41] ), .S(\mult_22/SUMB[44][41] ) );
  FA_X1 \mult_22/S2_44_40  ( .A(\mult_22/ab[44][40] ), .B(
        \mult_22/CARRYB[43][40] ), .CI(\mult_22/SUMB[43][41] ), .CO(
        \mult_22/CARRYB[44][40] ), .S(\mult_22/SUMB[44][40] ) );
  FA_X1 \mult_22/S2_44_39  ( .A(\mult_22/ab[44][39] ), .B(
        \mult_22/CARRYB[43][39] ), .CI(\mult_22/SUMB[43][40] ), .CO(
        \mult_22/CARRYB[44][39] ), .S(\mult_22/SUMB[44][39] ) );
  FA_X1 \mult_22/S2_44_38  ( .A(\mult_22/ab[44][38] ), .B(
        \mult_22/CARRYB[43][38] ), .CI(\mult_22/SUMB[43][39] ), .CO(
        \mult_22/CARRYB[44][38] ), .S(\mult_22/SUMB[44][38] ) );
  FA_X1 \mult_22/S2_44_37  ( .A(\mult_22/ab[44][37] ), .B(
        \mult_22/CARRYB[43][37] ), .CI(\mult_22/SUMB[43][38] ), .CO(
        \mult_22/CARRYB[44][37] ), .S(\mult_22/SUMB[44][37] ) );
  FA_X1 \mult_22/S2_44_36  ( .A(\mult_22/ab[44][36] ), .B(
        \mult_22/CARRYB[43][36] ), .CI(\mult_22/SUMB[43][37] ), .CO(
        \mult_22/CARRYB[44][36] ), .S(\mult_22/SUMB[44][36] ) );
  FA_X1 \mult_22/S2_44_35  ( .A(\mult_22/ab[44][35] ), .B(
        \mult_22/CARRYB[43][35] ), .CI(\mult_22/SUMB[43][36] ), .CO(
        \mult_22/CARRYB[44][35] ), .S(\mult_22/SUMB[44][35] ) );
  FA_X1 \mult_22/S2_44_34  ( .A(\mult_22/ab[44][34] ), .B(
        \mult_22/CARRYB[43][34] ), .CI(\mult_22/SUMB[43][35] ), .CO(
        \mult_22/CARRYB[44][34] ), .S(\mult_22/SUMB[44][34] ) );
  FA_X1 \mult_22/S2_44_33  ( .A(\mult_22/ab[44][33] ), .B(
        \mult_22/CARRYB[43][33] ), .CI(\mult_22/SUMB[43][34] ), .CO(
        \mult_22/CARRYB[44][33] ), .S(\mult_22/SUMB[44][33] ) );
  FA_X1 \mult_22/S2_44_32  ( .A(\mult_22/ab[44][32] ), .B(
        \mult_22/CARRYB[43][32] ), .CI(\mult_22/SUMB[43][33] ), .CO(
        \mult_22/CARRYB[44][32] ), .S(\mult_22/SUMB[44][32] ) );
  FA_X1 \mult_22/S2_44_31  ( .A(\mult_22/ab[44][31] ), .B(
        \mult_22/CARRYB[43][31] ), .CI(\mult_22/SUMB[43][32] ), .CO(
        \mult_22/CARRYB[44][31] ), .S(\mult_22/SUMB[44][31] ) );
  FA_X1 \mult_22/S2_44_30  ( .A(\mult_22/ab[44][30] ), .B(
        \mult_22/CARRYB[43][30] ), .CI(\mult_22/SUMB[43][31] ), .CO(
        \mult_22/CARRYB[44][30] ), .S(\mult_22/SUMB[44][30] ) );
  FA_X1 \mult_22/S2_44_29  ( .A(\mult_22/ab[44][29] ), .B(
        \mult_22/CARRYB[43][29] ), .CI(\mult_22/SUMB[43][30] ), .CO(
        \mult_22/CARRYB[44][29] ), .S(\mult_22/SUMB[44][29] ) );
  FA_X1 \mult_22/S2_44_28  ( .A(\mult_22/ab[44][28] ), .B(
        \mult_22/CARRYB[43][28] ), .CI(\mult_22/SUMB[43][29] ), .CO(
        \mult_22/CARRYB[44][28] ), .S(\mult_22/SUMB[44][28] ) );
  FA_X1 \mult_22/S2_44_27  ( .A(\mult_22/ab[44][27] ), .B(
        \mult_22/CARRYB[43][27] ), .CI(\mult_22/SUMB[43][28] ), .CO(
        \mult_22/CARRYB[44][27] ), .S(\mult_22/SUMB[44][27] ) );
  FA_X1 \mult_22/S2_44_26  ( .A(\mult_22/ab[44][26] ), .B(
        \mult_22/CARRYB[43][26] ), .CI(\mult_22/SUMB[43][27] ), .CO(
        \mult_22/CARRYB[44][26] ), .S(\mult_22/SUMB[44][26] ) );
  FA_X1 \mult_22/S2_44_25  ( .A(\mult_22/ab[44][25] ), .B(
        \mult_22/CARRYB[43][25] ), .CI(\mult_22/SUMB[43][26] ), .CO(
        \mult_22/CARRYB[44][25] ), .S(\mult_22/SUMB[44][25] ) );
  FA_X1 \mult_22/S2_44_24  ( .A(\mult_22/ab[44][24] ), .B(
        \mult_22/CARRYB[43][24] ), .CI(\mult_22/SUMB[43][25] ), .CO(
        \mult_22/CARRYB[44][24] ), .S(\mult_22/SUMB[44][24] ) );
  FA_X1 \mult_22/S2_44_23  ( .A(\mult_22/ab[44][23] ), .B(
        \mult_22/CARRYB[43][23] ), .CI(\mult_22/SUMB[43][24] ), .CO(
        \mult_22/CARRYB[44][23] ), .S(\mult_22/SUMB[44][23] ) );
  FA_X1 \mult_22/S2_44_22  ( .A(\mult_22/CARRYB[43][22] ), .B(
        \mult_22/ab[44][22] ), .CI(\mult_22/SUMB[43][23] ), .CO(
        \mult_22/CARRYB[44][22] ), .S(\mult_22/SUMB[44][22] ) );
  FA_X1 \mult_22/S2_44_21  ( .A(\mult_22/ab[44][21] ), .B(
        \mult_22/CARRYB[43][21] ), .CI(\mult_22/SUMB[43][22] ), .CO(
        \mult_22/CARRYB[44][21] ), .S(\mult_22/SUMB[44][21] ) );
  FA_X1 \mult_22/S2_44_20  ( .A(\mult_22/ab[44][20] ), .B(
        \mult_22/CARRYB[43][20] ), .CI(\mult_22/SUMB[43][21] ), .CO(
        \mult_22/CARRYB[44][20] ), .S(\mult_22/SUMB[44][20] ) );
  FA_X1 \mult_22/S2_44_19  ( .A(\mult_22/ab[44][19] ), .B(
        \mult_22/CARRYB[43][19] ), .CI(\mult_22/SUMB[43][20] ), .CO(
        \mult_22/CARRYB[44][19] ), .S(\mult_22/SUMB[44][19] ) );
  FA_X1 \mult_22/S2_44_18  ( .A(\mult_22/ab[44][18] ), .B(
        \mult_22/CARRYB[43][18] ), .CI(\mult_22/SUMB[43][19] ), .CO(
        \mult_22/CARRYB[44][18] ), .S(\mult_22/SUMB[44][18] ) );
  FA_X1 \mult_22/S2_44_17  ( .A(\mult_22/ab[44][17] ), .B(
        \mult_22/CARRYB[43][17] ), .CI(\mult_22/SUMB[43][18] ), .CO(
        \mult_22/CARRYB[44][17] ), .S(\mult_22/SUMB[44][17] ) );
  FA_X1 \mult_22/S2_44_16  ( .A(\mult_22/ab[44][16] ), .B(
        \mult_22/CARRYB[43][16] ), .CI(\mult_22/SUMB[43][17] ), .CO(
        \mult_22/CARRYB[44][16] ), .S(\mult_22/SUMB[44][16] ) );
  FA_X1 \mult_22/S2_44_15  ( .A(\mult_22/ab[44][15] ), .B(
        \mult_22/CARRYB[43][15] ), .CI(\mult_22/SUMB[43][16] ), .CO(
        \mult_22/CARRYB[44][15] ), .S(\mult_22/SUMB[44][15] ) );
  FA_X1 \mult_22/S2_44_14  ( .A(\mult_22/ab[44][14] ), .B(
        \mult_22/CARRYB[43][14] ), .CI(\mult_22/SUMB[43][15] ), .CO(
        \mult_22/CARRYB[44][14] ), .S(\mult_22/SUMB[44][14] ) );
  FA_X1 \mult_22/S2_44_13  ( .A(\mult_22/ab[44][13] ), .B(
        \mult_22/CARRYB[43][13] ), .CI(\mult_22/SUMB[43][14] ), .CO(
        \mult_22/CARRYB[44][13] ), .S(\mult_22/SUMB[44][13] ) );
  FA_X1 \mult_22/S2_44_12  ( .A(\mult_22/ab[44][12] ), .B(
        \mult_22/CARRYB[43][12] ), .CI(\mult_22/SUMB[43][13] ), .CO(
        \mult_22/CARRYB[44][12] ), .S(\mult_22/SUMB[44][12] ) );
  FA_X1 \mult_22/S2_44_11  ( .A(\mult_22/ab[44][11] ), .B(
        \mult_22/CARRYB[43][11] ), .CI(\mult_22/SUMB[43][12] ), .CO(
        \mult_22/CARRYB[44][11] ), .S(\mult_22/SUMB[44][11] ) );
  FA_X1 \mult_22/S2_44_10  ( .A(\mult_22/ab[44][10] ), .B(
        \mult_22/CARRYB[43][10] ), .CI(\mult_22/SUMB[43][11] ), .CO(
        \mult_22/CARRYB[44][10] ), .S(\mult_22/SUMB[44][10] ) );
  FA_X1 \mult_22/S2_44_9  ( .A(\mult_22/ab[44][9] ), .B(
        \mult_22/CARRYB[43][9] ), .CI(\mult_22/SUMB[43][10] ), .CO(
        \mult_22/CARRYB[44][9] ), .S(\mult_22/SUMB[44][9] ) );
  FA_X1 \mult_22/S2_44_8  ( .A(\mult_22/ab[44][8] ), .B(
        \mult_22/CARRYB[43][8] ), .CI(\mult_22/SUMB[43][9] ), .CO(
        \mult_22/CARRYB[44][8] ), .S(\mult_22/SUMB[44][8] ) );
  FA_X1 \mult_22/S2_44_7  ( .A(\mult_22/ab[44][7] ), .B(
        \mult_22/CARRYB[43][7] ), .CI(\mult_22/SUMB[43][8] ), .CO(
        \mult_22/CARRYB[44][7] ), .S(\mult_22/SUMB[44][7] ) );
  FA_X1 \mult_22/S2_44_6  ( .A(\mult_22/ab[44][6] ), .B(
        \mult_22/CARRYB[43][6] ), .CI(\mult_22/SUMB[43][7] ), .CO(
        \mult_22/CARRYB[44][6] ), .S(\mult_22/SUMB[44][6] ) );
  FA_X1 \mult_22/S2_44_5  ( .A(\mult_22/ab[44][5] ), .B(
        \mult_22/CARRYB[43][5] ), .CI(\mult_22/SUMB[43][6] ), .CO(
        \mult_22/CARRYB[44][5] ), .S(\mult_22/SUMB[44][5] ) );
  FA_X1 \mult_22/S2_44_4  ( .A(\mult_22/ab[44][4] ), .B(
        \mult_22/CARRYB[43][4] ), .CI(\mult_22/SUMB[43][5] ), .CO(
        \mult_22/CARRYB[44][4] ), .S(\mult_22/SUMB[44][4] ) );
  FA_X1 \mult_22/S2_44_3  ( .A(\mult_22/ab[44][3] ), .B(
        \mult_22/CARRYB[43][3] ), .CI(\mult_22/SUMB[43][4] ), .CO(
        \mult_22/CARRYB[44][3] ), .S(\mult_22/SUMB[44][3] ) );
  FA_X1 \mult_22/S2_44_2  ( .A(\mult_22/ab[44][2] ), .B(
        \mult_22/CARRYB[43][2] ), .CI(\mult_22/SUMB[43][3] ), .CO(
        \mult_22/CARRYB[44][2] ), .S(\mult_22/SUMB[44][2] ) );
  FA_X1 \mult_22/S2_44_1  ( .A(\mult_22/ab[44][1] ), .B(
        \mult_22/CARRYB[43][1] ), .CI(\mult_22/SUMB[43][2] ), .CO(
        \mult_22/CARRYB[44][1] ), .S(\mult_22/SUMB[44][1] ) );
  FA_X1 \mult_22/S1_44_0  ( .A(\mult_22/ab[44][0] ), .B(
        \mult_22/CARRYB[43][0] ), .CI(\mult_22/SUMB[43][1] ), .CO(
        \mult_22/CARRYB[44][0] ), .S(N172) );
  FA_X1 \mult_22/S3_45_62  ( .A(\mult_22/ab[45][62] ), .B(
        \mult_22/CARRYB[44][62] ), .CI(\mult_22/ab[44][63] ), .CO(
        \mult_22/CARRYB[45][62] ), .S(\mult_22/SUMB[45][62] ) );
  FA_X1 \mult_22/S2_45_61  ( .A(\mult_22/ab[45][61] ), .B(
        \mult_22/CARRYB[44][61] ), .CI(\mult_22/SUMB[44][62] ), .CO(
        \mult_22/CARRYB[45][61] ), .S(\mult_22/SUMB[45][61] ) );
  FA_X1 \mult_22/S2_45_60  ( .A(\mult_22/ab[45][60] ), .B(
        \mult_22/CARRYB[44][60] ), .CI(\mult_22/SUMB[44][61] ), .CO(
        \mult_22/CARRYB[45][60] ), .S(\mult_22/SUMB[45][60] ) );
  FA_X1 \mult_22/S2_45_59  ( .A(\mult_22/ab[45][59] ), .B(
        \mult_22/CARRYB[44][59] ), .CI(\mult_22/SUMB[44][60] ), .CO(
        \mult_22/CARRYB[45][59] ), .S(\mult_22/SUMB[45][59] ) );
  FA_X1 \mult_22/S2_45_58  ( .A(\mult_22/ab[45][58] ), .B(
        \mult_22/CARRYB[44][58] ), .CI(\mult_22/SUMB[44][59] ), .CO(
        \mult_22/CARRYB[45][58] ), .S(\mult_22/SUMB[45][58] ) );
  FA_X1 \mult_22/S2_45_57  ( .A(\mult_22/ab[45][57] ), .B(
        \mult_22/CARRYB[44][57] ), .CI(\mult_22/SUMB[44][58] ), .CO(
        \mult_22/CARRYB[45][57] ), .S(\mult_22/SUMB[45][57] ) );
  FA_X1 \mult_22/S2_45_56  ( .A(\mult_22/ab[45][56] ), .B(
        \mult_22/CARRYB[44][56] ), .CI(\mult_22/SUMB[44][57] ), .CO(
        \mult_22/CARRYB[45][56] ), .S(\mult_22/SUMB[45][56] ) );
  FA_X1 \mult_22/S2_45_55  ( .A(\mult_22/ab[45][55] ), .B(
        \mult_22/CARRYB[44][55] ), .CI(\mult_22/SUMB[44][56] ), .CO(
        \mult_22/CARRYB[45][55] ), .S(\mult_22/SUMB[45][55] ) );
  FA_X1 \mult_22/S2_45_54  ( .A(\mult_22/ab[45][54] ), .B(
        \mult_22/CARRYB[44][54] ), .CI(\mult_22/SUMB[44][55] ), .CO(
        \mult_22/CARRYB[45][54] ), .S(\mult_22/SUMB[45][54] ) );
  FA_X1 \mult_22/S2_45_53  ( .A(\mult_22/ab[45][53] ), .B(
        \mult_22/CARRYB[44][53] ), .CI(\mult_22/SUMB[44][54] ), .CO(
        \mult_22/CARRYB[45][53] ), .S(\mult_22/SUMB[45][53] ) );
  FA_X1 \mult_22/S2_45_52  ( .A(\mult_22/ab[45][52] ), .B(
        \mult_22/CARRYB[44][52] ), .CI(\mult_22/SUMB[44][53] ), .CO(
        \mult_22/CARRYB[45][52] ), .S(\mult_22/SUMB[45][52] ) );
  FA_X1 \mult_22/S2_45_51  ( .A(\mult_22/ab[45][51] ), .B(
        \mult_22/CARRYB[44][51] ), .CI(\mult_22/SUMB[44][52] ), .CO(
        \mult_22/CARRYB[45][51] ), .S(\mult_22/SUMB[45][51] ) );
  FA_X1 \mult_22/S2_45_50  ( .A(\mult_22/ab[45][50] ), .B(
        \mult_22/CARRYB[44][50] ), .CI(\mult_22/SUMB[44][51] ), .CO(
        \mult_22/CARRYB[45][50] ), .S(\mult_22/SUMB[45][50] ) );
  FA_X1 \mult_22/S2_45_49  ( .A(\mult_22/ab[45][49] ), .B(
        \mult_22/CARRYB[44][49] ), .CI(\mult_22/SUMB[44][50] ), .CO(
        \mult_22/CARRYB[45][49] ), .S(\mult_22/SUMB[45][49] ) );
  FA_X1 \mult_22/S2_45_48  ( .A(\mult_22/ab[45][48] ), .B(
        \mult_22/CARRYB[44][48] ), .CI(\mult_22/SUMB[44][49] ), .CO(
        \mult_22/CARRYB[45][48] ), .S(\mult_22/SUMB[45][48] ) );
  FA_X1 \mult_22/S2_45_47  ( .A(\mult_22/ab[45][47] ), .B(
        \mult_22/CARRYB[44][47] ), .CI(\mult_22/SUMB[44][48] ), .CO(
        \mult_22/CARRYB[45][47] ), .S(\mult_22/SUMB[45][47] ) );
  FA_X1 \mult_22/S2_45_46  ( .A(\mult_22/ab[45][46] ), .B(
        \mult_22/CARRYB[44][46] ), .CI(\mult_22/SUMB[44][47] ), .CO(
        \mult_22/CARRYB[45][46] ), .S(\mult_22/SUMB[45][46] ) );
  FA_X1 \mult_22/S2_45_45  ( .A(\mult_22/ab[45][45] ), .B(
        \mult_22/CARRYB[44][45] ), .CI(\mult_22/SUMB[44][46] ), .CO(
        \mult_22/CARRYB[45][45] ), .S(\mult_22/SUMB[45][45] ) );
  FA_X1 \mult_22/S2_45_44  ( .A(\mult_22/ab[45][44] ), .B(
        \mult_22/CARRYB[44][44] ), .CI(\mult_22/SUMB[44][45] ), .CO(
        \mult_22/CARRYB[45][44] ), .S(\mult_22/SUMB[45][44] ) );
  FA_X1 \mult_22/S2_45_43  ( .A(\mult_22/ab[45][43] ), .B(
        \mult_22/CARRYB[44][43] ), .CI(\mult_22/SUMB[44][44] ), .CO(
        \mult_22/CARRYB[45][43] ), .S(\mult_22/SUMB[45][43] ) );
  FA_X1 \mult_22/S2_45_42  ( .A(\mult_22/ab[45][42] ), .B(
        \mult_22/CARRYB[44][42] ), .CI(\mult_22/SUMB[44][43] ), .CO(
        \mult_22/CARRYB[45][42] ), .S(\mult_22/SUMB[45][42] ) );
  FA_X1 \mult_22/S2_45_41  ( .A(\mult_22/ab[45][41] ), .B(
        \mult_22/CARRYB[44][41] ), .CI(\mult_22/SUMB[44][42] ), .CO(
        \mult_22/CARRYB[45][41] ), .S(\mult_22/SUMB[45][41] ) );
  FA_X1 \mult_22/S2_45_40  ( .A(\mult_22/ab[45][40] ), .B(
        \mult_22/CARRYB[44][40] ), .CI(\mult_22/SUMB[44][41] ), .CO(
        \mult_22/CARRYB[45][40] ), .S(\mult_22/SUMB[45][40] ) );
  FA_X1 \mult_22/S2_45_39  ( .A(\mult_22/ab[45][39] ), .B(
        \mult_22/CARRYB[44][39] ), .CI(\mult_22/SUMB[44][40] ), .CO(
        \mult_22/CARRYB[45][39] ), .S(\mult_22/SUMB[45][39] ) );
  FA_X1 \mult_22/S2_45_38  ( .A(\mult_22/ab[45][38] ), .B(
        \mult_22/CARRYB[44][38] ), .CI(\mult_22/SUMB[44][39] ), .CO(
        \mult_22/CARRYB[45][38] ), .S(\mult_22/SUMB[45][38] ) );
  FA_X1 \mult_22/S2_45_37  ( .A(\mult_22/ab[45][37] ), .B(
        \mult_22/CARRYB[44][37] ), .CI(\mult_22/SUMB[44][38] ), .CO(
        \mult_22/CARRYB[45][37] ), .S(\mult_22/SUMB[45][37] ) );
  FA_X1 \mult_22/S2_45_36  ( .A(\mult_22/ab[45][36] ), .B(
        \mult_22/CARRYB[44][36] ), .CI(\mult_22/SUMB[44][37] ), .CO(
        \mult_22/CARRYB[45][36] ), .S(\mult_22/SUMB[45][36] ) );
  FA_X1 \mult_22/S2_45_35  ( .A(\mult_22/ab[45][35] ), .B(
        \mult_22/CARRYB[44][35] ), .CI(\mult_22/SUMB[44][36] ), .CO(
        \mult_22/CARRYB[45][35] ), .S(\mult_22/SUMB[45][35] ) );
  FA_X1 \mult_22/S2_45_34  ( .A(\mult_22/ab[45][34] ), .B(
        \mult_22/CARRYB[44][34] ), .CI(\mult_22/SUMB[44][35] ), .CO(
        \mult_22/CARRYB[45][34] ), .S(\mult_22/SUMB[45][34] ) );
  FA_X1 \mult_22/S2_45_33  ( .A(\mult_22/ab[45][33] ), .B(
        \mult_22/CARRYB[44][33] ), .CI(\mult_22/SUMB[44][34] ), .CO(
        \mult_22/CARRYB[45][33] ), .S(\mult_22/SUMB[45][33] ) );
  FA_X1 \mult_22/S2_45_32  ( .A(\mult_22/ab[45][32] ), .B(
        \mult_22/CARRYB[44][32] ), .CI(\mult_22/SUMB[44][33] ), .CO(
        \mult_22/CARRYB[45][32] ), .S(\mult_22/SUMB[45][32] ) );
  FA_X1 \mult_22/S2_45_31  ( .A(\mult_22/ab[45][31] ), .B(
        \mult_22/CARRYB[44][31] ), .CI(\mult_22/SUMB[44][32] ), .CO(
        \mult_22/CARRYB[45][31] ), .S(\mult_22/SUMB[45][31] ) );
  FA_X1 \mult_22/S2_45_30  ( .A(\mult_22/ab[45][30] ), .B(
        \mult_22/CARRYB[44][30] ), .CI(\mult_22/SUMB[44][31] ), .CO(
        \mult_22/CARRYB[45][30] ), .S(\mult_22/SUMB[45][30] ) );
  FA_X1 \mult_22/S2_45_29  ( .A(\mult_22/ab[45][29] ), .B(
        \mult_22/CARRYB[44][29] ), .CI(\mult_22/SUMB[44][30] ), .CO(
        \mult_22/CARRYB[45][29] ), .S(\mult_22/SUMB[45][29] ) );
  FA_X1 \mult_22/S2_45_28  ( .A(\mult_22/ab[45][28] ), .B(
        \mult_22/CARRYB[44][28] ), .CI(\mult_22/SUMB[44][29] ), .CO(
        \mult_22/CARRYB[45][28] ), .S(\mult_22/SUMB[45][28] ) );
  FA_X1 \mult_22/S2_45_27  ( .A(\mult_22/ab[45][27] ), .B(
        \mult_22/CARRYB[44][27] ), .CI(\mult_22/SUMB[44][28] ), .CO(
        \mult_22/CARRYB[45][27] ), .S(\mult_22/SUMB[45][27] ) );
  FA_X1 \mult_22/S2_45_26  ( .A(\mult_22/ab[45][26] ), .B(
        \mult_22/CARRYB[44][26] ), .CI(\mult_22/SUMB[44][27] ), .CO(
        \mult_22/CARRYB[45][26] ), .S(\mult_22/SUMB[45][26] ) );
  FA_X1 \mult_22/S2_45_25  ( .A(\mult_22/ab[45][25] ), .B(
        \mult_22/CARRYB[44][25] ), .CI(\mult_22/SUMB[44][26] ), .CO(
        \mult_22/CARRYB[45][25] ), .S(\mult_22/SUMB[45][25] ) );
  FA_X1 \mult_22/S2_45_24  ( .A(\mult_22/ab[45][24] ), .B(
        \mult_22/CARRYB[44][24] ), .CI(\mult_22/SUMB[44][25] ), .CO(
        \mult_22/CARRYB[45][24] ), .S(\mult_22/SUMB[45][24] ) );
  FA_X1 \mult_22/S2_45_23  ( .A(\mult_22/ab[45][23] ), .B(
        \mult_22/CARRYB[44][23] ), .CI(\mult_22/SUMB[44][24] ), .CO(
        \mult_22/CARRYB[45][23] ), .S(\mult_22/SUMB[45][23] ) );
  FA_X1 \mult_22/S2_45_22  ( .A(\mult_22/CARRYB[44][22] ), .B(
        \mult_22/ab[45][22] ), .CI(\mult_22/SUMB[44][23] ), .CO(
        \mult_22/CARRYB[45][22] ), .S(\mult_22/SUMB[45][22] ) );
  FA_X1 \mult_22/S2_45_21  ( .A(\mult_22/CARRYB[44][21] ), .B(
        \mult_22/ab[45][21] ), .CI(\mult_22/SUMB[44][22] ), .CO(
        \mult_22/CARRYB[45][21] ), .S(\mult_22/SUMB[45][21] ) );
  FA_X1 \mult_22/S2_45_20  ( .A(\mult_22/CARRYB[44][20] ), .B(
        \mult_22/ab[45][20] ), .CI(\mult_22/SUMB[44][21] ), .CO(
        \mult_22/CARRYB[45][20] ), .S(\mult_22/SUMB[45][20] ) );
  FA_X1 \mult_22/S2_45_19  ( .A(\mult_22/ab[45][19] ), .B(
        \mult_22/CARRYB[44][19] ), .CI(\mult_22/SUMB[44][20] ), .CO(
        \mult_22/CARRYB[45][19] ), .S(\mult_22/SUMB[45][19] ) );
  FA_X1 \mult_22/S2_45_18  ( .A(\mult_22/ab[45][18] ), .B(
        \mult_22/CARRYB[44][18] ), .CI(\mult_22/SUMB[44][19] ), .CO(
        \mult_22/CARRYB[45][18] ), .S(\mult_22/SUMB[45][18] ) );
  FA_X1 \mult_22/S2_45_17  ( .A(\mult_22/ab[45][17] ), .B(
        \mult_22/CARRYB[44][17] ), .CI(\mult_22/SUMB[44][18] ), .CO(
        \mult_22/CARRYB[45][17] ), .S(\mult_22/SUMB[45][17] ) );
  FA_X1 \mult_22/S2_45_16  ( .A(\mult_22/ab[45][16] ), .B(
        \mult_22/CARRYB[44][16] ), .CI(\mult_22/SUMB[44][17] ), .CO(
        \mult_22/CARRYB[45][16] ), .S(\mult_22/SUMB[45][16] ) );
  FA_X1 \mult_22/S2_45_15  ( .A(\mult_22/ab[45][15] ), .B(
        \mult_22/CARRYB[44][15] ), .CI(\mult_22/SUMB[44][16] ), .CO(
        \mult_22/CARRYB[45][15] ), .S(\mult_22/SUMB[45][15] ) );
  FA_X1 \mult_22/S2_45_14  ( .A(\mult_22/ab[45][14] ), .B(
        \mult_22/CARRYB[44][14] ), .CI(\mult_22/SUMB[44][15] ), .CO(
        \mult_22/CARRYB[45][14] ), .S(\mult_22/SUMB[45][14] ) );
  FA_X1 \mult_22/S2_45_13  ( .A(\mult_22/ab[45][13] ), .B(
        \mult_22/CARRYB[44][13] ), .CI(\mult_22/SUMB[44][14] ), .CO(
        \mult_22/CARRYB[45][13] ), .S(\mult_22/SUMB[45][13] ) );
  FA_X1 \mult_22/S2_45_12  ( .A(\mult_22/ab[45][12] ), .B(
        \mult_22/CARRYB[44][12] ), .CI(\mult_22/SUMB[44][13] ), .CO(
        \mult_22/CARRYB[45][12] ), .S(\mult_22/SUMB[45][12] ) );
  FA_X1 \mult_22/S2_45_11  ( .A(\mult_22/ab[45][11] ), .B(
        \mult_22/CARRYB[44][11] ), .CI(\mult_22/SUMB[44][12] ), .CO(
        \mult_22/CARRYB[45][11] ), .S(\mult_22/SUMB[45][11] ) );
  FA_X1 \mult_22/S2_45_10  ( .A(\mult_22/ab[45][10] ), .B(
        \mult_22/CARRYB[44][10] ), .CI(\mult_22/SUMB[44][11] ), .CO(
        \mult_22/CARRYB[45][10] ), .S(\mult_22/SUMB[45][10] ) );
  FA_X1 \mult_22/S2_45_9  ( .A(\mult_22/ab[45][9] ), .B(
        \mult_22/CARRYB[44][9] ), .CI(\mult_22/SUMB[44][10] ), .CO(
        \mult_22/CARRYB[45][9] ), .S(\mult_22/SUMB[45][9] ) );
  FA_X1 \mult_22/S2_45_8  ( .A(\mult_22/ab[45][8] ), .B(
        \mult_22/CARRYB[44][8] ), .CI(\mult_22/SUMB[44][9] ), .CO(
        \mult_22/CARRYB[45][8] ), .S(\mult_22/SUMB[45][8] ) );
  FA_X1 \mult_22/S2_45_7  ( .A(\mult_22/ab[45][7] ), .B(
        \mult_22/CARRYB[44][7] ), .CI(\mult_22/SUMB[44][8] ), .CO(
        \mult_22/CARRYB[45][7] ), .S(\mult_22/SUMB[45][7] ) );
  FA_X1 \mult_22/S2_45_6  ( .A(\mult_22/ab[45][6] ), .B(
        \mult_22/CARRYB[44][6] ), .CI(\mult_22/SUMB[44][7] ), .CO(
        \mult_22/CARRYB[45][6] ), .S(\mult_22/SUMB[45][6] ) );
  FA_X1 \mult_22/S2_45_5  ( .A(\mult_22/ab[45][5] ), .B(
        \mult_22/CARRYB[44][5] ), .CI(\mult_22/SUMB[44][6] ), .CO(
        \mult_22/CARRYB[45][5] ), .S(\mult_22/SUMB[45][5] ) );
  FA_X1 \mult_22/S2_45_4  ( .A(\mult_22/ab[45][4] ), .B(
        \mult_22/CARRYB[44][4] ), .CI(\mult_22/SUMB[44][5] ), .CO(
        \mult_22/CARRYB[45][4] ), .S(\mult_22/SUMB[45][4] ) );
  FA_X1 \mult_22/S2_45_3  ( .A(\mult_22/ab[45][3] ), .B(
        \mult_22/CARRYB[44][3] ), .CI(\mult_22/SUMB[44][4] ), .CO(
        \mult_22/CARRYB[45][3] ), .S(\mult_22/SUMB[45][3] ) );
  FA_X1 \mult_22/S2_45_2  ( .A(\mult_22/ab[45][2] ), .B(
        \mult_22/CARRYB[44][2] ), .CI(\mult_22/SUMB[44][3] ), .CO(
        \mult_22/CARRYB[45][2] ), .S(\mult_22/SUMB[45][2] ) );
  FA_X1 \mult_22/S2_45_1  ( .A(\mult_22/ab[45][1] ), .B(
        \mult_22/CARRYB[44][1] ), .CI(\mult_22/SUMB[44][2] ), .CO(
        \mult_22/CARRYB[45][1] ), .S(\mult_22/SUMB[45][1] ) );
  FA_X1 \mult_22/S1_45_0  ( .A(\mult_22/ab[45][0] ), .B(
        \mult_22/CARRYB[44][0] ), .CI(\mult_22/SUMB[44][1] ), .CO(
        \mult_22/CARRYB[45][0] ), .S(N173) );
  FA_X1 \mult_22/S3_46_62  ( .A(\mult_22/ab[46][62] ), .B(
        \mult_22/CARRYB[45][62] ), .CI(\mult_22/ab[45][63] ), .CO(
        \mult_22/CARRYB[46][62] ), .S(\mult_22/SUMB[46][62] ) );
  FA_X1 \mult_22/S2_46_61  ( .A(\mult_22/ab[46][61] ), .B(
        \mult_22/CARRYB[45][61] ), .CI(\mult_22/SUMB[45][62] ), .CO(
        \mult_22/CARRYB[46][61] ), .S(\mult_22/SUMB[46][61] ) );
  FA_X1 \mult_22/S2_46_60  ( .A(\mult_22/ab[46][60] ), .B(
        \mult_22/CARRYB[45][60] ), .CI(\mult_22/SUMB[45][61] ), .CO(
        \mult_22/CARRYB[46][60] ), .S(\mult_22/SUMB[46][60] ) );
  FA_X1 \mult_22/S2_46_59  ( .A(\mult_22/ab[46][59] ), .B(
        \mult_22/CARRYB[45][59] ), .CI(\mult_22/SUMB[45][60] ), .CO(
        \mult_22/CARRYB[46][59] ), .S(\mult_22/SUMB[46][59] ) );
  FA_X1 \mult_22/S2_46_58  ( .A(\mult_22/ab[46][58] ), .B(
        \mult_22/CARRYB[45][58] ), .CI(\mult_22/SUMB[45][59] ), .CO(
        \mult_22/CARRYB[46][58] ), .S(\mult_22/SUMB[46][58] ) );
  FA_X1 \mult_22/S2_46_57  ( .A(\mult_22/ab[46][57] ), .B(
        \mult_22/CARRYB[45][57] ), .CI(\mult_22/SUMB[45][58] ), .CO(
        \mult_22/CARRYB[46][57] ), .S(\mult_22/SUMB[46][57] ) );
  FA_X1 \mult_22/S2_46_56  ( .A(\mult_22/ab[46][56] ), .B(
        \mult_22/CARRYB[45][56] ), .CI(\mult_22/SUMB[45][57] ), .CO(
        \mult_22/CARRYB[46][56] ), .S(\mult_22/SUMB[46][56] ) );
  FA_X1 \mult_22/S2_46_55  ( .A(\mult_22/ab[46][55] ), .B(
        \mult_22/CARRYB[45][55] ), .CI(\mult_22/SUMB[45][56] ), .CO(
        \mult_22/CARRYB[46][55] ), .S(\mult_22/SUMB[46][55] ) );
  FA_X1 \mult_22/S2_46_54  ( .A(\mult_22/ab[46][54] ), .B(
        \mult_22/CARRYB[45][54] ), .CI(\mult_22/SUMB[45][55] ), .CO(
        \mult_22/CARRYB[46][54] ), .S(\mult_22/SUMB[46][54] ) );
  FA_X1 \mult_22/S2_46_53  ( .A(\mult_22/ab[46][53] ), .B(
        \mult_22/CARRYB[45][53] ), .CI(\mult_22/SUMB[45][54] ), .CO(
        \mult_22/CARRYB[46][53] ), .S(\mult_22/SUMB[46][53] ) );
  FA_X1 \mult_22/S2_46_52  ( .A(\mult_22/ab[46][52] ), .B(
        \mult_22/CARRYB[45][52] ), .CI(\mult_22/SUMB[45][53] ), .CO(
        \mult_22/CARRYB[46][52] ), .S(\mult_22/SUMB[46][52] ) );
  FA_X1 \mult_22/S2_46_51  ( .A(\mult_22/ab[46][51] ), .B(
        \mult_22/CARRYB[45][51] ), .CI(\mult_22/SUMB[45][52] ), .CO(
        \mult_22/CARRYB[46][51] ), .S(\mult_22/SUMB[46][51] ) );
  FA_X1 \mult_22/S2_46_50  ( .A(\mult_22/ab[46][50] ), .B(
        \mult_22/CARRYB[45][50] ), .CI(\mult_22/SUMB[45][51] ), .CO(
        \mult_22/CARRYB[46][50] ), .S(\mult_22/SUMB[46][50] ) );
  FA_X1 \mult_22/S2_46_49  ( .A(\mult_22/ab[46][49] ), .B(
        \mult_22/CARRYB[45][49] ), .CI(\mult_22/SUMB[45][50] ), .CO(
        \mult_22/CARRYB[46][49] ), .S(\mult_22/SUMB[46][49] ) );
  FA_X1 \mult_22/S2_46_48  ( .A(\mult_22/ab[46][48] ), .B(
        \mult_22/CARRYB[45][48] ), .CI(\mult_22/SUMB[45][49] ), .CO(
        \mult_22/CARRYB[46][48] ), .S(\mult_22/SUMB[46][48] ) );
  FA_X1 \mult_22/S2_46_47  ( .A(\mult_22/ab[46][47] ), .B(
        \mult_22/CARRYB[45][47] ), .CI(\mult_22/SUMB[45][48] ), .CO(
        \mult_22/CARRYB[46][47] ), .S(\mult_22/SUMB[46][47] ) );
  FA_X1 \mult_22/S2_46_46  ( .A(\mult_22/ab[46][46] ), .B(
        \mult_22/CARRYB[45][46] ), .CI(\mult_22/SUMB[45][47] ), .CO(
        \mult_22/CARRYB[46][46] ), .S(\mult_22/SUMB[46][46] ) );
  FA_X1 \mult_22/S2_46_45  ( .A(\mult_22/ab[46][45] ), .B(
        \mult_22/CARRYB[45][45] ), .CI(\mult_22/SUMB[45][46] ), .CO(
        \mult_22/CARRYB[46][45] ), .S(\mult_22/SUMB[46][45] ) );
  FA_X1 \mult_22/S2_46_44  ( .A(\mult_22/ab[46][44] ), .B(
        \mult_22/CARRYB[45][44] ), .CI(\mult_22/SUMB[45][45] ), .CO(
        \mult_22/CARRYB[46][44] ), .S(\mult_22/SUMB[46][44] ) );
  FA_X1 \mult_22/S2_46_43  ( .A(\mult_22/ab[46][43] ), .B(
        \mult_22/CARRYB[45][43] ), .CI(\mult_22/SUMB[45][44] ), .CO(
        \mult_22/CARRYB[46][43] ), .S(\mult_22/SUMB[46][43] ) );
  FA_X1 \mult_22/S2_46_42  ( .A(\mult_22/ab[46][42] ), .B(
        \mult_22/CARRYB[45][42] ), .CI(\mult_22/SUMB[45][43] ), .CO(
        \mult_22/CARRYB[46][42] ), .S(\mult_22/SUMB[46][42] ) );
  FA_X1 \mult_22/S2_46_41  ( .A(\mult_22/ab[46][41] ), .B(
        \mult_22/CARRYB[45][41] ), .CI(\mult_22/SUMB[45][42] ), .CO(
        \mult_22/CARRYB[46][41] ), .S(\mult_22/SUMB[46][41] ) );
  FA_X1 \mult_22/S2_46_40  ( .A(\mult_22/ab[46][40] ), .B(
        \mult_22/CARRYB[45][40] ), .CI(\mult_22/SUMB[45][41] ), .CO(
        \mult_22/CARRYB[46][40] ), .S(\mult_22/SUMB[46][40] ) );
  FA_X1 \mult_22/S2_46_39  ( .A(\mult_22/ab[46][39] ), .B(
        \mult_22/CARRYB[45][39] ), .CI(\mult_22/SUMB[45][40] ), .CO(
        \mult_22/CARRYB[46][39] ), .S(\mult_22/SUMB[46][39] ) );
  FA_X1 \mult_22/S2_46_38  ( .A(\mult_22/ab[46][38] ), .B(
        \mult_22/CARRYB[45][38] ), .CI(\mult_22/SUMB[45][39] ), .CO(
        \mult_22/CARRYB[46][38] ), .S(\mult_22/SUMB[46][38] ) );
  FA_X1 \mult_22/S2_46_37  ( .A(\mult_22/ab[46][37] ), .B(
        \mult_22/CARRYB[45][37] ), .CI(\mult_22/SUMB[45][38] ), .CO(
        \mult_22/CARRYB[46][37] ), .S(\mult_22/SUMB[46][37] ) );
  FA_X1 \mult_22/S2_46_36  ( .A(\mult_22/ab[46][36] ), .B(
        \mult_22/CARRYB[45][36] ), .CI(\mult_22/SUMB[45][37] ), .CO(
        \mult_22/CARRYB[46][36] ), .S(\mult_22/SUMB[46][36] ) );
  FA_X1 \mult_22/S2_46_35  ( .A(\mult_22/ab[46][35] ), .B(
        \mult_22/CARRYB[45][35] ), .CI(\mult_22/SUMB[45][36] ), .CO(
        \mult_22/CARRYB[46][35] ), .S(\mult_22/SUMB[46][35] ) );
  FA_X1 \mult_22/S2_46_34  ( .A(\mult_22/ab[46][34] ), .B(
        \mult_22/CARRYB[45][34] ), .CI(\mult_22/SUMB[45][35] ), .CO(
        \mult_22/CARRYB[46][34] ), .S(\mult_22/SUMB[46][34] ) );
  FA_X1 \mult_22/S2_46_33  ( .A(\mult_22/ab[46][33] ), .B(
        \mult_22/CARRYB[45][33] ), .CI(\mult_22/SUMB[45][34] ), .CO(
        \mult_22/CARRYB[46][33] ), .S(\mult_22/SUMB[46][33] ) );
  FA_X1 \mult_22/S2_46_32  ( .A(\mult_22/ab[46][32] ), .B(
        \mult_22/CARRYB[45][32] ), .CI(\mult_22/SUMB[45][33] ), .CO(
        \mult_22/CARRYB[46][32] ), .S(\mult_22/SUMB[46][32] ) );
  FA_X1 \mult_22/S2_46_31  ( .A(\mult_22/ab[46][31] ), .B(
        \mult_22/CARRYB[45][31] ), .CI(\mult_22/SUMB[45][32] ), .CO(
        \mult_22/CARRYB[46][31] ), .S(\mult_22/SUMB[46][31] ) );
  FA_X1 \mult_22/S2_46_30  ( .A(\mult_22/ab[46][30] ), .B(
        \mult_22/CARRYB[45][30] ), .CI(\mult_22/SUMB[45][31] ), .CO(
        \mult_22/CARRYB[46][30] ), .S(\mult_22/SUMB[46][30] ) );
  FA_X1 \mult_22/S2_46_29  ( .A(\mult_22/ab[46][29] ), .B(
        \mult_22/CARRYB[45][29] ), .CI(\mult_22/SUMB[45][30] ), .CO(
        \mult_22/CARRYB[46][29] ), .S(\mult_22/SUMB[46][29] ) );
  FA_X1 \mult_22/S2_46_28  ( .A(\mult_22/ab[46][28] ), .B(
        \mult_22/CARRYB[45][28] ), .CI(\mult_22/SUMB[45][29] ), .CO(
        \mult_22/CARRYB[46][28] ), .S(\mult_22/SUMB[46][28] ) );
  FA_X1 \mult_22/S2_46_27  ( .A(\mult_22/ab[46][27] ), .B(
        \mult_22/CARRYB[45][27] ), .CI(\mult_22/SUMB[45][28] ), .CO(
        \mult_22/CARRYB[46][27] ), .S(\mult_22/SUMB[46][27] ) );
  FA_X1 \mult_22/S2_46_26  ( .A(\mult_22/ab[46][26] ), .B(
        \mult_22/CARRYB[45][26] ), .CI(\mult_22/SUMB[45][27] ), .CO(
        \mult_22/CARRYB[46][26] ), .S(\mult_22/SUMB[46][26] ) );
  FA_X1 \mult_22/S2_46_25  ( .A(\mult_22/ab[46][25] ), .B(
        \mult_22/CARRYB[45][25] ), .CI(\mult_22/SUMB[45][26] ), .CO(
        \mult_22/CARRYB[46][25] ), .S(\mult_22/SUMB[46][25] ) );
  FA_X1 \mult_22/S2_46_24  ( .A(\mult_22/ab[46][24] ), .B(
        \mult_22/CARRYB[45][24] ), .CI(\mult_22/SUMB[45][25] ), .CO(
        \mult_22/CARRYB[46][24] ), .S(\mult_22/SUMB[46][24] ) );
  FA_X1 \mult_22/S2_46_23  ( .A(\mult_22/ab[46][23] ), .B(
        \mult_22/CARRYB[45][23] ), .CI(\mult_22/SUMB[45][24] ), .CO(
        \mult_22/CARRYB[46][23] ), .S(\mult_22/SUMB[46][23] ) );
  FA_X1 \mult_22/S2_46_22  ( .A(\mult_22/ab[46][22] ), .B(
        \mult_22/CARRYB[45][22] ), .CI(\mult_22/SUMB[45][23] ), .CO(
        \mult_22/CARRYB[46][22] ), .S(\mult_22/SUMB[46][22] ) );
  FA_X1 \mult_22/S2_46_21  ( .A(\mult_22/ab[46][21] ), .B(
        \mult_22/CARRYB[45][21] ), .CI(\mult_22/SUMB[45][22] ), .CO(
        \mult_22/CARRYB[46][21] ), .S(\mult_22/SUMB[46][21] ) );
  FA_X1 \mult_22/S2_46_20  ( .A(\mult_22/ab[46][20] ), .B(
        \mult_22/CARRYB[45][20] ), .CI(\mult_22/SUMB[45][21] ), .CO(
        \mult_22/CARRYB[46][20] ), .S(\mult_22/SUMB[46][20] ) );
  FA_X1 \mult_22/S2_46_19  ( .A(\mult_22/ab[46][19] ), .B(
        \mult_22/CARRYB[45][19] ), .CI(\mult_22/SUMB[45][20] ), .CO(
        \mult_22/CARRYB[46][19] ), .S(\mult_22/SUMB[46][19] ) );
  FA_X1 \mult_22/S2_46_18  ( .A(\mult_22/ab[46][18] ), .B(
        \mult_22/CARRYB[45][18] ), .CI(\mult_22/SUMB[45][19] ), .CO(
        \mult_22/CARRYB[46][18] ), .S(\mult_22/SUMB[46][18] ) );
  FA_X1 \mult_22/S2_46_17  ( .A(\mult_22/CARRYB[45][17] ), .B(
        \mult_22/ab[46][17] ), .CI(\mult_22/SUMB[45][18] ), .CO(
        \mult_22/CARRYB[46][17] ), .S(\mult_22/SUMB[46][17] ) );
  FA_X1 \mult_22/S2_46_16  ( .A(\mult_22/ab[46][16] ), .B(
        \mult_22/CARRYB[45][16] ), .CI(\mult_22/SUMB[45][17] ), .CO(
        \mult_22/CARRYB[46][16] ), .S(\mult_22/SUMB[46][16] ) );
  FA_X1 \mult_22/S2_46_15  ( .A(\mult_22/ab[46][15] ), .B(
        \mult_22/CARRYB[45][15] ), .CI(\mult_22/SUMB[45][16] ), .CO(
        \mult_22/CARRYB[46][15] ), .S(\mult_22/SUMB[46][15] ) );
  FA_X1 \mult_22/S2_46_14  ( .A(\mult_22/ab[46][14] ), .B(
        \mult_22/CARRYB[45][14] ), .CI(\mult_22/SUMB[45][15] ), .CO(
        \mult_22/CARRYB[46][14] ), .S(\mult_22/SUMB[46][14] ) );
  FA_X1 \mult_22/S2_46_13  ( .A(\mult_22/ab[46][13] ), .B(
        \mult_22/CARRYB[45][13] ), .CI(\mult_22/SUMB[45][14] ), .CO(
        \mult_22/CARRYB[46][13] ), .S(\mult_22/SUMB[46][13] ) );
  FA_X1 \mult_22/S2_46_12  ( .A(\mult_22/ab[46][12] ), .B(
        \mult_22/CARRYB[45][12] ), .CI(\mult_22/SUMB[45][13] ), .CO(
        \mult_22/CARRYB[46][12] ), .S(\mult_22/SUMB[46][12] ) );
  FA_X1 \mult_22/S2_46_11  ( .A(\mult_22/ab[46][11] ), .B(
        \mult_22/CARRYB[45][11] ), .CI(\mult_22/SUMB[45][12] ), .CO(
        \mult_22/CARRYB[46][11] ), .S(\mult_22/SUMB[46][11] ) );
  FA_X1 \mult_22/S2_46_10  ( .A(\mult_22/ab[46][10] ), .B(
        \mult_22/CARRYB[45][10] ), .CI(\mult_22/SUMB[45][11] ), .CO(
        \mult_22/CARRYB[46][10] ), .S(\mult_22/SUMB[46][10] ) );
  FA_X1 \mult_22/S2_46_9  ( .A(\mult_22/ab[46][9] ), .B(
        \mult_22/CARRYB[45][9] ), .CI(\mult_22/SUMB[45][10] ), .CO(
        \mult_22/CARRYB[46][9] ), .S(\mult_22/SUMB[46][9] ) );
  FA_X1 \mult_22/S2_46_8  ( .A(\mult_22/ab[46][8] ), .B(
        \mult_22/CARRYB[45][8] ), .CI(\mult_22/SUMB[45][9] ), .CO(
        \mult_22/CARRYB[46][8] ), .S(\mult_22/SUMB[46][8] ) );
  FA_X1 \mult_22/S2_46_7  ( .A(\mult_22/ab[46][7] ), .B(
        \mult_22/CARRYB[45][7] ), .CI(\mult_22/SUMB[45][8] ), .CO(
        \mult_22/CARRYB[46][7] ), .S(\mult_22/SUMB[46][7] ) );
  FA_X1 \mult_22/S2_46_6  ( .A(\mult_22/ab[46][6] ), .B(
        \mult_22/CARRYB[45][6] ), .CI(\mult_22/SUMB[45][7] ), .CO(
        \mult_22/CARRYB[46][6] ), .S(\mult_22/SUMB[46][6] ) );
  FA_X1 \mult_22/S2_46_5  ( .A(\mult_22/ab[46][5] ), .B(
        \mult_22/CARRYB[45][5] ), .CI(\mult_22/SUMB[45][6] ), .CO(
        \mult_22/CARRYB[46][5] ), .S(\mult_22/SUMB[46][5] ) );
  FA_X1 \mult_22/S2_46_4  ( .A(\mult_22/ab[46][4] ), .B(
        \mult_22/CARRYB[45][4] ), .CI(\mult_22/SUMB[45][5] ), .CO(
        \mult_22/CARRYB[46][4] ), .S(\mult_22/SUMB[46][4] ) );
  FA_X1 \mult_22/S2_46_3  ( .A(\mult_22/ab[46][3] ), .B(
        \mult_22/CARRYB[45][3] ), .CI(\mult_22/SUMB[45][4] ), .CO(
        \mult_22/CARRYB[46][3] ), .S(\mult_22/SUMB[46][3] ) );
  FA_X1 \mult_22/S2_46_2  ( .A(\mult_22/ab[46][2] ), .B(
        \mult_22/CARRYB[45][2] ), .CI(\mult_22/SUMB[45][3] ), .CO(
        \mult_22/CARRYB[46][2] ), .S(\mult_22/SUMB[46][2] ) );
  FA_X1 \mult_22/S2_46_1  ( .A(\mult_22/ab[46][1] ), .B(
        \mult_22/CARRYB[45][1] ), .CI(\mult_22/SUMB[45][2] ), .CO(
        \mult_22/CARRYB[46][1] ), .S(\mult_22/SUMB[46][1] ) );
  FA_X1 \mult_22/S1_46_0  ( .A(\mult_22/ab[46][0] ), .B(
        \mult_22/CARRYB[45][0] ), .CI(\mult_22/SUMB[45][1] ), .CO(
        \mult_22/CARRYB[46][0] ), .S(N174) );
  FA_X1 \mult_22/S3_47_62  ( .A(\mult_22/ab[47][62] ), .B(
        \mult_22/CARRYB[46][62] ), .CI(\mult_22/ab[46][63] ), .CO(
        \mult_22/CARRYB[47][62] ), .S(\mult_22/SUMB[47][62] ) );
  FA_X1 \mult_22/S2_47_61  ( .A(\mult_22/ab[47][61] ), .B(
        \mult_22/CARRYB[46][61] ), .CI(\mult_22/SUMB[46][62] ), .CO(
        \mult_22/CARRYB[47][61] ), .S(\mult_22/SUMB[47][61] ) );
  FA_X1 \mult_22/S2_47_60  ( .A(\mult_22/ab[47][60] ), .B(
        \mult_22/CARRYB[46][60] ), .CI(\mult_22/SUMB[46][61] ), .CO(
        \mult_22/CARRYB[47][60] ), .S(\mult_22/SUMB[47][60] ) );
  FA_X1 \mult_22/S2_47_59  ( .A(\mult_22/ab[47][59] ), .B(
        \mult_22/CARRYB[46][59] ), .CI(\mult_22/SUMB[46][60] ), .CO(
        \mult_22/CARRYB[47][59] ), .S(\mult_22/SUMB[47][59] ) );
  FA_X1 \mult_22/S2_47_58  ( .A(\mult_22/ab[47][58] ), .B(
        \mult_22/CARRYB[46][58] ), .CI(\mult_22/SUMB[46][59] ), .CO(
        \mult_22/CARRYB[47][58] ), .S(\mult_22/SUMB[47][58] ) );
  FA_X1 \mult_22/S2_47_57  ( .A(\mult_22/ab[47][57] ), .B(
        \mult_22/CARRYB[46][57] ), .CI(\mult_22/SUMB[46][58] ), .CO(
        \mult_22/CARRYB[47][57] ), .S(\mult_22/SUMB[47][57] ) );
  FA_X1 \mult_22/S2_47_56  ( .A(\mult_22/ab[47][56] ), .B(
        \mult_22/CARRYB[46][56] ), .CI(\mult_22/SUMB[46][57] ), .CO(
        \mult_22/CARRYB[47][56] ), .S(\mult_22/SUMB[47][56] ) );
  FA_X1 \mult_22/S2_47_55  ( .A(\mult_22/ab[47][55] ), .B(
        \mult_22/CARRYB[46][55] ), .CI(\mult_22/SUMB[46][56] ), .CO(
        \mult_22/CARRYB[47][55] ), .S(\mult_22/SUMB[47][55] ) );
  FA_X1 \mult_22/S2_47_54  ( .A(\mult_22/ab[47][54] ), .B(
        \mult_22/CARRYB[46][54] ), .CI(\mult_22/SUMB[46][55] ), .CO(
        \mult_22/CARRYB[47][54] ), .S(\mult_22/SUMB[47][54] ) );
  FA_X1 \mult_22/S2_47_53  ( .A(\mult_22/ab[47][53] ), .B(
        \mult_22/CARRYB[46][53] ), .CI(\mult_22/SUMB[46][54] ), .CO(
        \mult_22/CARRYB[47][53] ), .S(\mult_22/SUMB[47][53] ) );
  FA_X1 \mult_22/S2_47_52  ( .A(\mult_22/ab[47][52] ), .B(
        \mult_22/CARRYB[46][52] ), .CI(\mult_22/SUMB[46][53] ), .CO(
        \mult_22/CARRYB[47][52] ), .S(\mult_22/SUMB[47][52] ) );
  FA_X1 \mult_22/S2_47_51  ( .A(\mult_22/ab[47][51] ), .B(
        \mult_22/CARRYB[46][51] ), .CI(\mult_22/SUMB[46][52] ), .CO(
        \mult_22/CARRYB[47][51] ), .S(\mult_22/SUMB[47][51] ) );
  FA_X1 \mult_22/S2_47_50  ( .A(\mult_22/ab[47][50] ), .B(
        \mult_22/CARRYB[46][50] ), .CI(\mult_22/SUMB[46][51] ), .CO(
        \mult_22/CARRYB[47][50] ), .S(\mult_22/SUMB[47][50] ) );
  FA_X1 \mult_22/S2_47_49  ( .A(\mult_22/ab[47][49] ), .B(
        \mult_22/CARRYB[46][49] ), .CI(\mult_22/SUMB[46][50] ), .CO(
        \mult_22/CARRYB[47][49] ), .S(\mult_22/SUMB[47][49] ) );
  FA_X1 \mult_22/S2_47_48  ( .A(\mult_22/ab[47][48] ), .B(
        \mult_22/CARRYB[46][48] ), .CI(\mult_22/SUMB[46][49] ), .CO(
        \mult_22/CARRYB[47][48] ), .S(\mult_22/SUMB[47][48] ) );
  FA_X1 \mult_22/S2_47_47  ( .A(\mult_22/ab[47][47] ), .B(
        \mult_22/CARRYB[46][47] ), .CI(\mult_22/SUMB[46][48] ), .CO(
        \mult_22/CARRYB[47][47] ), .S(\mult_22/SUMB[47][47] ) );
  FA_X1 \mult_22/S2_47_46  ( .A(\mult_22/ab[47][46] ), .B(
        \mult_22/CARRYB[46][46] ), .CI(\mult_22/SUMB[46][47] ), .CO(
        \mult_22/CARRYB[47][46] ), .S(\mult_22/SUMB[47][46] ) );
  FA_X1 \mult_22/S2_47_45  ( .A(\mult_22/ab[47][45] ), .B(
        \mult_22/CARRYB[46][45] ), .CI(\mult_22/SUMB[46][46] ), .CO(
        \mult_22/CARRYB[47][45] ), .S(\mult_22/SUMB[47][45] ) );
  FA_X1 \mult_22/S2_47_44  ( .A(\mult_22/ab[47][44] ), .B(
        \mult_22/CARRYB[46][44] ), .CI(\mult_22/SUMB[46][45] ), .CO(
        \mult_22/CARRYB[47][44] ), .S(\mult_22/SUMB[47][44] ) );
  FA_X1 \mult_22/S2_47_43  ( .A(\mult_22/ab[47][43] ), .B(
        \mult_22/CARRYB[46][43] ), .CI(\mult_22/SUMB[46][44] ), .CO(
        \mult_22/CARRYB[47][43] ), .S(\mult_22/SUMB[47][43] ) );
  FA_X1 \mult_22/S2_47_42  ( .A(\mult_22/ab[47][42] ), .B(
        \mult_22/CARRYB[46][42] ), .CI(\mult_22/SUMB[46][43] ), .CO(
        \mult_22/CARRYB[47][42] ), .S(\mult_22/SUMB[47][42] ) );
  FA_X1 \mult_22/S2_47_41  ( .A(\mult_22/ab[47][41] ), .B(
        \mult_22/CARRYB[46][41] ), .CI(\mult_22/SUMB[46][42] ), .CO(
        \mult_22/CARRYB[47][41] ), .S(\mult_22/SUMB[47][41] ) );
  FA_X1 \mult_22/S2_47_40  ( .A(\mult_22/ab[47][40] ), .B(
        \mult_22/CARRYB[46][40] ), .CI(\mult_22/SUMB[46][41] ), .CO(
        \mult_22/CARRYB[47][40] ), .S(\mult_22/SUMB[47][40] ) );
  FA_X1 \mult_22/S2_47_39  ( .A(\mult_22/ab[47][39] ), .B(
        \mult_22/CARRYB[46][39] ), .CI(\mult_22/SUMB[46][40] ), .CO(
        \mult_22/CARRYB[47][39] ), .S(\mult_22/SUMB[47][39] ) );
  FA_X1 \mult_22/S2_47_38  ( .A(\mult_22/ab[47][38] ), .B(
        \mult_22/CARRYB[46][38] ), .CI(\mult_22/SUMB[46][39] ), .CO(
        \mult_22/CARRYB[47][38] ), .S(\mult_22/SUMB[47][38] ) );
  FA_X1 \mult_22/S2_47_37  ( .A(\mult_22/ab[47][37] ), .B(
        \mult_22/CARRYB[46][37] ), .CI(\mult_22/SUMB[46][38] ), .CO(
        \mult_22/CARRYB[47][37] ), .S(\mult_22/SUMB[47][37] ) );
  FA_X1 \mult_22/S2_47_36  ( .A(\mult_22/ab[47][36] ), .B(
        \mult_22/CARRYB[46][36] ), .CI(\mult_22/SUMB[46][37] ), .CO(
        \mult_22/CARRYB[47][36] ), .S(\mult_22/SUMB[47][36] ) );
  FA_X1 \mult_22/S2_47_35  ( .A(\mult_22/ab[47][35] ), .B(
        \mult_22/CARRYB[46][35] ), .CI(\mult_22/SUMB[46][36] ), .CO(
        \mult_22/CARRYB[47][35] ), .S(\mult_22/SUMB[47][35] ) );
  FA_X1 \mult_22/S2_47_34  ( .A(\mult_22/ab[47][34] ), .B(
        \mult_22/CARRYB[46][34] ), .CI(\mult_22/SUMB[46][35] ), .CO(
        \mult_22/CARRYB[47][34] ), .S(\mult_22/SUMB[47][34] ) );
  FA_X1 \mult_22/S2_47_33  ( .A(\mult_22/ab[47][33] ), .B(
        \mult_22/CARRYB[46][33] ), .CI(\mult_22/SUMB[46][34] ), .CO(
        \mult_22/CARRYB[47][33] ), .S(\mult_22/SUMB[47][33] ) );
  FA_X1 \mult_22/S2_47_32  ( .A(\mult_22/ab[47][32] ), .B(
        \mult_22/CARRYB[46][32] ), .CI(\mult_22/SUMB[46][33] ), .CO(
        \mult_22/CARRYB[47][32] ), .S(\mult_22/SUMB[47][32] ) );
  FA_X1 \mult_22/S2_47_31  ( .A(\mult_22/ab[47][31] ), .B(
        \mult_22/CARRYB[46][31] ), .CI(\mult_22/SUMB[46][32] ), .CO(
        \mult_22/CARRYB[47][31] ), .S(\mult_22/SUMB[47][31] ) );
  FA_X1 \mult_22/S2_47_30  ( .A(\mult_22/ab[47][30] ), .B(
        \mult_22/CARRYB[46][30] ), .CI(\mult_22/SUMB[46][31] ), .CO(
        \mult_22/CARRYB[47][30] ), .S(\mult_22/SUMB[47][30] ) );
  FA_X1 \mult_22/S2_47_29  ( .A(\mult_22/ab[47][29] ), .B(
        \mult_22/CARRYB[46][29] ), .CI(\mult_22/SUMB[46][30] ), .CO(
        \mult_22/CARRYB[47][29] ), .S(\mult_22/SUMB[47][29] ) );
  FA_X1 \mult_22/S2_47_28  ( .A(\mult_22/ab[47][28] ), .B(
        \mult_22/CARRYB[46][28] ), .CI(\mult_22/SUMB[46][29] ), .CO(
        \mult_22/CARRYB[47][28] ), .S(\mult_22/SUMB[47][28] ) );
  FA_X1 \mult_22/S2_47_27  ( .A(\mult_22/ab[47][27] ), .B(
        \mult_22/CARRYB[46][27] ), .CI(\mult_22/SUMB[46][28] ), .CO(
        \mult_22/CARRYB[47][27] ), .S(\mult_22/SUMB[47][27] ) );
  FA_X1 \mult_22/S2_47_26  ( .A(\mult_22/ab[47][26] ), .B(
        \mult_22/CARRYB[46][26] ), .CI(\mult_22/SUMB[46][27] ), .CO(
        \mult_22/CARRYB[47][26] ), .S(\mult_22/SUMB[47][26] ) );
  FA_X1 \mult_22/S2_47_25  ( .A(\mult_22/ab[47][25] ), .B(
        \mult_22/CARRYB[46][25] ), .CI(\mult_22/SUMB[46][26] ), .CO(
        \mult_22/CARRYB[47][25] ), .S(\mult_22/SUMB[47][25] ) );
  FA_X1 \mult_22/S2_47_24  ( .A(\mult_22/ab[47][24] ), .B(
        \mult_22/CARRYB[46][24] ), .CI(\mult_22/SUMB[46][25] ), .CO(
        \mult_22/CARRYB[47][24] ), .S(\mult_22/SUMB[47][24] ) );
  FA_X1 \mult_22/S2_47_23  ( .A(\mult_22/ab[47][23] ), .B(
        \mult_22/CARRYB[46][23] ), .CI(\mult_22/SUMB[46][24] ), .CO(
        \mult_22/CARRYB[47][23] ), .S(\mult_22/SUMB[47][23] ) );
  FA_X1 \mult_22/S2_47_22  ( .A(\mult_22/ab[47][22] ), .B(
        \mult_22/CARRYB[46][22] ), .CI(\mult_22/SUMB[46][23] ), .CO(
        \mult_22/CARRYB[47][22] ), .S(\mult_22/SUMB[47][22] ) );
  FA_X1 \mult_22/S2_47_21  ( .A(\mult_22/ab[47][21] ), .B(
        \mult_22/CARRYB[46][21] ), .CI(\mult_22/SUMB[46][22] ), .CO(
        \mult_22/CARRYB[47][21] ), .S(\mult_22/SUMB[47][21] ) );
  FA_X1 \mult_22/S2_47_20  ( .A(\mult_22/CARRYB[46][20] ), .B(
        \mult_22/ab[47][20] ), .CI(\mult_22/SUMB[46][21] ), .CO(
        \mult_22/CARRYB[47][20] ), .S(\mult_22/SUMB[47][20] ) );
  FA_X1 \mult_22/S2_47_19  ( .A(\mult_22/CARRYB[46][19] ), .B(
        \mult_22/ab[47][19] ), .CI(\mult_22/SUMB[46][20] ), .CO(
        \mult_22/CARRYB[47][19] ), .S(\mult_22/SUMB[47][19] ) );
  FA_X1 \mult_22/S2_47_18  ( .A(\mult_22/ab[47][18] ), .B(
        \mult_22/CARRYB[46][18] ), .CI(\mult_22/SUMB[46][19] ), .CO(
        \mult_22/CARRYB[47][18] ), .S(\mult_22/SUMB[47][18] ) );
  FA_X1 \mult_22/S2_47_17  ( .A(\mult_22/ab[47][17] ), .B(
        \mult_22/CARRYB[46][17] ), .CI(\mult_22/SUMB[46][18] ), .CO(
        \mult_22/CARRYB[47][17] ), .S(\mult_22/SUMB[47][17] ) );
  FA_X1 \mult_22/S2_47_16  ( .A(\mult_22/ab[47][16] ), .B(
        \mult_22/CARRYB[46][16] ), .CI(\mult_22/SUMB[46][17] ), .CO(
        \mult_22/CARRYB[47][16] ), .S(\mult_22/SUMB[47][16] ) );
  FA_X1 \mult_22/S2_47_15  ( .A(\mult_22/ab[47][15] ), .B(
        \mult_22/CARRYB[46][15] ), .CI(\mult_22/SUMB[46][16] ), .CO(
        \mult_22/CARRYB[47][15] ), .S(\mult_22/SUMB[47][15] ) );
  FA_X1 \mult_22/S2_47_14  ( .A(\mult_22/ab[47][14] ), .B(
        \mult_22/CARRYB[46][14] ), .CI(\mult_22/SUMB[46][15] ), .CO(
        \mult_22/CARRYB[47][14] ), .S(\mult_22/SUMB[47][14] ) );
  FA_X1 \mult_22/S2_47_13  ( .A(\mult_22/ab[47][13] ), .B(
        \mult_22/CARRYB[46][13] ), .CI(\mult_22/SUMB[46][14] ), .CO(
        \mult_22/CARRYB[47][13] ), .S(\mult_22/SUMB[47][13] ) );
  FA_X1 \mult_22/S2_47_12  ( .A(\mult_22/ab[47][12] ), .B(
        \mult_22/CARRYB[46][12] ), .CI(\mult_22/SUMB[46][13] ), .CO(
        \mult_22/CARRYB[47][12] ), .S(\mult_22/SUMB[47][12] ) );
  FA_X1 \mult_22/S2_47_11  ( .A(\mult_22/ab[47][11] ), .B(
        \mult_22/CARRYB[46][11] ), .CI(\mult_22/SUMB[46][12] ), .CO(
        \mult_22/CARRYB[47][11] ), .S(\mult_22/SUMB[47][11] ) );
  FA_X1 \mult_22/S2_47_10  ( .A(\mult_22/ab[47][10] ), .B(
        \mult_22/CARRYB[46][10] ), .CI(\mult_22/SUMB[46][11] ), .CO(
        \mult_22/CARRYB[47][10] ), .S(\mult_22/SUMB[47][10] ) );
  FA_X1 \mult_22/S2_47_9  ( .A(\mult_22/ab[47][9] ), .B(
        \mult_22/CARRYB[46][9] ), .CI(\mult_22/SUMB[46][10] ), .CO(
        \mult_22/CARRYB[47][9] ), .S(\mult_22/SUMB[47][9] ) );
  FA_X1 \mult_22/S2_47_8  ( .A(\mult_22/ab[47][8] ), .B(
        \mult_22/CARRYB[46][8] ), .CI(\mult_22/SUMB[46][9] ), .CO(
        \mult_22/CARRYB[47][8] ), .S(\mult_22/SUMB[47][8] ) );
  FA_X1 \mult_22/S2_47_7  ( .A(\mult_22/ab[47][7] ), .B(
        \mult_22/CARRYB[46][7] ), .CI(\mult_22/SUMB[46][8] ), .CO(
        \mult_22/CARRYB[47][7] ), .S(\mult_22/SUMB[47][7] ) );
  FA_X1 \mult_22/S2_47_6  ( .A(\mult_22/ab[47][6] ), .B(
        \mult_22/CARRYB[46][6] ), .CI(\mult_22/SUMB[46][7] ), .CO(
        \mult_22/CARRYB[47][6] ), .S(\mult_22/SUMB[47][6] ) );
  FA_X1 \mult_22/S2_47_5  ( .A(\mult_22/ab[47][5] ), .B(
        \mult_22/CARRYB[46][5] ), .CI(\mult_22/SUMB[46][6] ), .CO(
        \mult_22/CARRYB[47][5] ), .S(\mult_22/SUMB[47][5] ) );
  FA_X1 \mult_22/S2_47_4  ( .A(\mult_22/ab[47][4] ), .B(
        \mult_22/CARRYB[46][4] ), .CI(\mult_22/SUMB[46][5] ), .CO(
        \mult_22/CARRYB[47][4] ), .S(\mult_22/SUMB[47][4] ) );
  FA_X1 \mult_22/S2_47_3  ( .A(\mult_22/ab[47][3] ), .B(
        \mult_22/CARRYB[46][3] ), .CI(\mult_22/SUMB[46][4] ), .CO(
        \mult_22/CARRYB[47][3] ), .S(\mult_22/SUMB[47][3] ) );
  FA_X1 \mult_22/S2_47_2  ( .A(\mult_22/ab[47][2] ), .B(
        \mult_22/CARRYB[46][2] ), .CI(\mult_22/SUMB[46][3] ), .CO(
        \mult_22/CARRYB[47][2] ), .S(\mult_22/SUMB[47][2] ) );
  FA_X1 \mult_22/S2_47_1  ( .A(\mult_22/ab[47][1] ), .B(
        \mult_22/CARRYB[46][1] ), .CI(\mult_22/SUMB[46][2] ), .CO(
        \mult_22/CARRYB[47][1] ), .S(\mult_22/SUMB[47][1] ) );
  FA_X1 \mult_22/S1_47_0  ( .A(\mult_22/ab[47][0] ), .B(
        \mult_22/CARRYB[46][0] ), .CI(\mult_22/SUMB[46][1] ), .CO(
        \mult_22/CARRYB[47][0] ), .S(N175) );
  FA_X1 \mult_22/S3_48_62  ( .A(\mult_22/ab[48][62] ), .B(
        \mult_22/CARRYB[47][62] ), .CI(\mult_22/ab[47][63] ), .CO(
        \mult_22/CARRYB[48][62] ), .S(\mult_22/SUMB[48][62] ) );
  FA_X1 \mult_22/S2_48_61  ( .A(\mult_22/ab[48][61] ), .B(
        \mult_22/CARRYB[47][61] ), .CI(\mult_22/SUMB[47][62] ), .CO(
        \mult_22/CARRYB[48][61] ), .S(\mult_22/SUMB[48][61] ) );
  FA_X1 \mult_22/S2_48_60  ( .A(\mult_22/ab[48][60] ), .B(
        \mult_22/CARRYB[47][60] ), .CI(\mult_22/SUMB[47][61] ), .CO(
        \mult_22/CARRYB[48][60] ), .S(\mult_22/SUMB[48][60] ) );
  FA_X1 \mult_22/S2_48_59  ( .A(\mult_22/ab[48][59] ), .B(
        \mult_22/CARRYB[47][59] ), .CI(\mult_22/SUMB[47][60] ), .CO(
        \mult_22/CARRYB[48][59] ), .S(\mult_22/SUMB[48][59] ) );
  FA_X1 \mult_22/S2_48_58  ( .A(\mult_22/ab[48][58] ), .B(
        \mult_22/CARRYB[47][58] ), .CI(\mult_22/SUMB[47][59] ), .CO(
        \mult_22/CARRYB[48][58] ), .S(\mult_22/SUMB[48][58] ) );
  FA_X1 \mult_22/S2_48_57  ( .A(\mult_22/ab[48][57] ), .B(
        \mult_22/CARRYB[47][57] ), .CI(\mult_22/SUMB[47][58] ), .CO(
        \mult_22/CARRYB[48][57] ), .S(\mult_22/SUMB[48][57] ) );
  FA_X1 \mult_22/S2_48_56  ( .A(\mult_22/ab[48][56] ), .B(
        \mult_22/CARRYB[47][56] ), .CI(\mult_22/SUMB[47][57] ), .CO(
        \mult_22/CARRYB[48][56] ), .S(\mult_22/SUMB[48][56] ) );
  FA_X1 \mult_22/S2_48_55  ( .A(\mult_22/ab[48][55] ), .B(
        \mult_22/CARRYB[47][55] ), .CI(\mult_22/SUMB[47][56] ), .CO(
        \mult_22/CARRYB[48][55] ), .S(\mult_22/SUMB[48][55] ) );
  FA_X1 \mult_22/S2_48_54  ( .A(\mult_22/ab[48][54] ), .B(
        \mult_22/CARRYB[47][54] ), .CI(\mult_22/SUMB[47][55] ), .CO(
        \mult_22/CARRYB[48][54] ), .S(\mult_22/SUMB[48][54] ) );
  FA_X1 \mult_22/S2_48_53  ( .A(\mult_22/ab[48][53] ), .B(
        \mult_22/CARRYB[47][53] ), .CI(\mult_22/SUMB[47][54] ), .CO(
        \mult_22/CARRYB[48][53] ), .S(\mult_22/SUMB[48][53] ) );
  FA_X1 \mult_22/S2_48_52  ( .A(\mult_22/ab[48][52] ), .B(
        \mult_22/CARRYB[47][52] ), .CI(\mult_22/SUMB[47][53] ), .CO(
        \mult_22/CARRYB[48][52] ), .S(\mult_22/SUMB[48][52] ) );
  FA_X1 \mult_22/S2_48_51  ( .A(\mult_22/ab[48][51] ), .B(
        \mult_22/CARRYB[47][51] ), .CI(\mult_22/SUMB[47][52] ), .CO(
        \mult_22/CARRYB[48][51] ), .S(\mult_22/SUMB[48][51] ) );
  FA_X1 \mult_22/S2_48_50  ( .A(\mult_22/ab[48][50] ), .B(
        \mult_22/CARRYB[47][50] ), .CI(\mult_22/SUMB[47][51] ), .CO(
        \mult_22/CARRYB[48][50] ), .S(\mult_22/SUMB[48][50] ) );
  FA_X1 \mult_22/S2_48_49  ( .A(\mult_22/ab[48][49] ), .B(
        \mult_22/CARRYB[47][49] ), .CI(\mult_22/SUMB[47][50] ), .CO(
        \mult_22/CARRYB[48][49] ), .S(\mult_22/SUMB[48][49] ) );
  FA_X1 \mult_22/S2_48_48  ( .A(\mult_22/ab[48][48] ), .B(
        \mult_22/CARRYB[47][48] ), .CI(\mult_22/SUMB[47][49] ), .CO(
        \mult_22/CARRYB[48][48] ), .S(\mult_22/SUMB[48][48] ) );
  FA_X1 \mult_22/S2_48_47  ( .A(\mult_22/ab[48][47] ), .B(
        \mult_22/CARRYB[47][47] ), .CI(\mult_22/SUMB[47][48] ), .CO(
        \mult_22/CARRYB[48][47] ), .S(\mult_22/SUMB[48][47] ) );
  FA_X1 \mult_22/S2_48_46  ( .A(\mult_22/ab[48][46] ), .B(
        \mult_22/CARRYB[47][46] ), .CI(\mult_22/SUMB[47][47] ), .CO(
        \mult_22/CARRYB[48][46] ), .S(\mult_22/SUMB[48][46] ) );
  FA_X1 \mult_22/S2_48_45  ( .A(\mult_22/ab[48][45] ), .B(
        \mult_22/CARRYB[47][45] ), .CI(\mult_22/SUMB[47][46] ), .CO(
        \mult_22/CARRYB[48][45] ), .S(\mult_22/SUMB[48][45] ) );
  FA_X1 \mult_22/S2_48_44  ( .A(\mult_22/ab[48][44] ), .B(
        \mult_22/CARRYB[47][44] ), .CI(\mult_22/SUMB[47][45] ), .CO(
        \mult_22/CARRYB[48][44] ), .S(\mult_22/SUMB[48][44] ) );
  FA_X1 \mult_22/S2_48_43  ( .A(\mult_22/ab[48][43] ), .B(
        \mult_22/CARRYB[47][43] ), .CI(\mult_22/SUMB[47][44] ), .CO(
        \mult_22/CARRYB[48][43] ), .S(\mult_22/SUMB[48][43] ) );
  FA_X1 \mult_22/S2_48_42  ( .A(\mult_22/ab[48][42] ), .B(
        \mult_22/CARRYB[47][42] ), .CI(\mult_22/SUMB[47][43] ), .CO(
        \mult_22/CARRYB[48][42] ), .S(\mult_22/SUMB[48][42] ) );
  FA_X1 \mult_22/S2_48_41  ( .A(\mult_22/ab[48][41] ), .B(
        \mult_22/CARRYB[47][41] ), .CI(\mult_22/SUMB[47][42] ), .CO(
        \mult_22/CARRYB[48][41] ), .S(\mult_22/SUMB[48][41] ) );
  FA_X1 \mult_22/S2_48_40  ( .A(\mult_22/ab[48][40] ), .B(
        \mult_22/CARRYB[47][40] ), .CI(\mult_22/SUMB[47][41] ), .CO(
        \mult_22/CARRYB[48][40] ), .S(\mult_22/SUMB[48][40] ) );
  FA_X1 \mult_22/S2_48_39  ( .A(\mult_22/ab[48][39] ), .B(
        \mult_22/CARRYB[47][39] ), .CI(\mult_22/SUMB[47][40] ), .CO(
        \mult_22/CARRYB[48][39] ), .S(\mult_22/SUMB[48][39] ) );
  FA_X1 \mult_22/S2_48_38  ( .A(\mult_22/ab[48][38] ), .B(
        \mult_22/CARRYB[47][38] ), .CI(\mult_22/SUMB[47][39] ), .CO(
        \mult_22/CARRYB[48][38] ), .S(\mult_22/SUMB[48][38] ) );
  FA_X1 \mult_22/S2_48_37  ( .A(\mult_22/ab[48][37] ), .B(
        \mult_22/CARRYB[47][37] ), .CI(\mult_22/SUMB[47][38] ), .CO(
        \mult_22/CARRYB[48][37] ), .S(\mult_22/SUMB[48][37] ) );
  FA_X1 \mult_22/S2_48_36  ( .A(\mult_22/ab[48][36] ), .B(
        \mult_22/CARRYB[47][36] ), .CI(\mult_22/SUMB[47][37] ), .CO(
        \mult_22/CARRYB[48][36] ), .S(\mult_22/SUMB[48][36] ) );
  FA_X1 \mult_22/S2_48_35  ( .A(\mult_22/ab[48][35] ), .B(
        \mult_22/CARRYB[47][35] ), .CI(\mult_22/SUMB[47][36] ), .CO(
        \mult_22/CARRYB[48][35] ), .S(\mult_22/SUMB[48][35] ) );
  FA_X1 \mult_22/S2_48_34  ( .A(\mult_22/ab[48][34] ), .B(
        \mult_22/CARRYB[47][34] ), .CI(\mult_22/SUMB[47][35] ), .CO(
        \mult_22/CARRYB[48][34] ), .S(\mult_22/SUMB[48][34] ) );
  FA_X1 \mult_22/S2_48_33  ( .A(\mult_22/ab[48][33] ), .B(
        \mult_22/CARRYB[47][33] ), .CI(\mult_22/SUMB[47][34] ), .CO(
        \mult_22/CARRYB[48][33] ), .S(\mult_22/SUMB[48][33] ) );
  FA_X1 \mult_22/S2_48_32  ( .A(\mult_22/ab[48][32] ), .B(
        \mult_22/CARRYB[47][32] ), .CI(\mult_22/SUMB[47][33] ), .CO(
        \mult_22/CARRYB[48][32] ), .S(\mult_22/SUMB[48][32] ) );
  FA_X1 \mult_22/S2_48_31  ( .A(\mult_22/ab[48][31] ), .B(
        \mult_22/CARRYB[47][31] ), .CI(\mult_22/SUMB[47][32] ), .CO(
        \mult_22/CARRYB[48][31] ), .S(\mult_22/SUMB[48][31] ) );
  FA_X1 \mult_22/S2_48_30  ( .A(\mult_22/ab[48][30] ), .B(
        \mult_22/CARRYB[47][30] ), .CI(\mult_22/SUMB[47][31] ), .CO(
        \mult_22/CARRYB[48][30] ), .S(\mult_22/SUMB[48][30] ) );
  FA_X1 \mult_22/S2_48_29  ( .A(\mult_22/ab[48][29] ), .B(
        \mult_22/CARRYB[47][29] ), .CI(\mult_22/SUMB[47][30] ), .CO(
        \mult_22/CARRYB[48][29] ), .S(\mult_22/SUMB[48][29] ) );
  FA_X1 \mult_22/S2_48_28  ( .A(\mult_22/ab[48][28] ), .B(
        \mult_22/CARRYB[47][28] ), .CI(\mult_22/SUMB[47][29] ), .CO(
        \mult_22/CARRYB[48][28] ), .S(\mult_22/SUMB[48][28] ) );
  FA_X1 \mult_22/S2_48_27  ( .A(\mult_22/ab[48][27] ), .B(
        \mult_22/CARRYB[47][27] ), .CI(\mult_22/SUMB[47][28] ), .CO(
        \mult_22/CARRYB[48][27] ), .S(\mult_22/SUMB[48][27] ) );
  FA_X1 \mult_22/S2_48_26  ( .A(\mult_22/ab[48][26] ), .B(
        \mult_22/CARRYB[47][26] ), .CI(\mult_22/SUMB[47][27] ), .CO(
        \mult_22/CARRYB[48][26] ), .S(\mult_22/SUMB[48][26] ) );
  FA_X1 \mult_22/S2_48_25  ( .A(\mult_22/ab[48][25] ), .B(
        \mult_22/CARRYB[47][25] ), .CI(\mult_22/SUMB[47][26] ), .CO(
        \mult_22/CARRYB[48][25] ), .S(\mult_22/SUMB[48][25] ) );
  FA_X1 \mult_22/S2_48_24  ( .A(\mult_22/ab[48][24] ), .B(
        \mult_22/CARRYB[47][24] ), .CI(\mult_22/SUMB[47][25] ), .CO(
        \mult_22/CARRYB[48][24] ), .S(\mult_22/SUMB[48][24] ) );
  FA_X1 \mult_22/S2_48_23  ( .A(\mult_22/ab[48][23] ), .B(
        \mult_22/CARRYB[47][23] ), .CI(\mult_22/SUMB[47][24] ), .CO(
        \mult_22/CARRYB[48][23] ), .S(\mult_22/SUMB[48][23] ) );
  FA_X1 \mult_22/S2_48_22  ( .A(\mult_22/ab[48][22] ), .B(
        \mult_22/CARRYB[47][22] ), .CI(\mult_22/SUMB[47][23] ), .CO(
        \mult_22/CARRYB[48][22] ), .S(\mult_22/SUMB[48][22] ) );
  FA_X1 \mult_22/S2_48_21  ( .A(\mult_22/ab[48][21] ), .B(
        \mult_22/CARRYB[47][21] ), .CI(\mult_22/SUMB[47][22] ), .CO(
        \mult_22/CARRYB[48][21] ), .S(\mult_22/SUMB[48][21] ) );
  FA_X1 \mult_22/S2_48_20  ( .A(\mult_22/ab[48][20] ), .B(
        \mult_22/CARRYB[47][20] ), .CI(\mult_22/SUMB[47][21] ), .CO(
        \mult_22/CARRYB[48][20] ), .S(\mult_22/SUMB[48][20] ) );
  FA_X1 \mult_22/S2_48_19  ( .A(\mult_22/ab[48][19] ), .B(
        \mult_22/CARRYB[47][19] ), .CI(\mult_22/SUMB[47][20] ), .CO(
        \mult_22/CARRYB[48][19] ), .S(\mult_22/SUMB[48][19] ) );
  FA_X1 \mult_22/S2_48_18  ( .A(\mult_22/ab[48][18] ), .B(
        \mult_22/CARRYB[47][18] ), .CI(\mult_22/SUMB[47][19] ), .CO(
        \mult_22/CARRYB[48][18] ), .S(\mult_22/SUMB[48][18] ) );
  FA_X1 \mult_22/S2_48_17  ( .A(\mult_22/ab[48][17] ), .B(
        \mult_22/CARRYB[47][17] ), .CI(\mult_22/SUMB[47][18] ), .CO(
        \mult_22/CARRYB[48][17] ), .S(\mult_22/SUMB[48][17] ) );
  FA_X1 \mult_22/S2_48_16  ( .A(\mult_22/ab[48][16] ), .B(
        \mult_22/CARRYB[47][16] ), .CI(\mult_22/SUMB[47][17] ), .CO(
        \mult_22/CARRYB[48][16] ), .S(\mult_22/SUMB[48][16] ) );
  FA_X1 \mult_22/S2_48_15  ( .A(\mult_22/CARRYB[47][15] ), .B(
        \mult_22/ab[48][15] ), .CI(\mult_22/SUMB[47][16] ), .CO(
        \mult_22/CARRYB[48][15] ), .S(\mult_22/SUMB[48][15] ) );
  FA_X1 \mult_22/S2_48_14  ( .A(\mult_22/ab[48][14] ), .B(
        \mult_22/CARRYB[47][14] ), .CI(\mult_22/SUMB[47][15] ), .CO(
        \mult_22/CARRYB[48][14] ), .S(\mult_22/SUMB[48][14] ) );
  FA_X1 \mult_22/S2_48_13  ( .A(\mult_22/ab[48][13] ), .B(
        \mult_22/CARRYB[47][13] ), .CI(\mult_22/SUMB[47][14] ), .CO(
        \mult_22/CARRYB[48][13] ), .S(\mult_22/SUMB[48][13] ) );
  FA_X1 \mult_22/S2_48_12  ( .A(\mult_22/ab[48][12] ), .B(
        \mult_22/CARRYB[47][12] ), .CI(\mult_22/SUMB[47][13] ), .CO(
        \mult_22/CARRYB[48][12] ), .S(\mult_22/SUMB[48][12] ) );
  FA_X1 \mult_22/S2_48_11  ( .A(\mult_22/ab[48][11] ), .B(
        \mult_22/CARRYB[47][11] ), .CI(\mult_22/SUMB[47][12] ), .CO(
        \mult_22/CARRYB[48][11] ), .S(\mult_22/SUMB[48][11] ) );
  FA_X1 \mult_22/S2_48_10  ( .A(\mult_22/ab[48][10] ), .B(
        \mult_22/CARRYB[47][10] ), .CI(\mult_22/SUMB[47][11] ), .CO(
        \mult_22/CARRYB[48][10] ), .S(\mult_22/SUMB[48][10] ) );
  FA_X1 \mult_22/S2_48_9  ( .A(\mult_22/ab[48][9] ), .B(
        \mult_22/CARRYB[47][9] ), .CI(\mult_22/SUMB[47][10] ), .CO(
        \mult_22/CARRYB[48][9] ), .S(\mult_22/SUMB[48][9] ) );
  FA_X1 \mult_22/S2_48_8  ( .A(\mult_22/ab[48][8] ), .B(
        \mult_22/CARRYB[47][8] ), .CI(\mult_22/SUMB[47][9] ), .CO(
        \mult_22/CARRYB[48][8] ), .S(\mult_22/SUMB[48][8] ) );
  FA_X1 \mult_22/S2_48_7  ( .A(\mult_22/ab[48][7] ), .B(
        \mult_22/CARRYB[47][7] ), .CI(\mult_22/SUMB[47][8] ), .CO(
        \mult_22/CARRYB[48][7] ), .S(\mult_22/SUMB[48][7] ) );
  FA_X1 \mult_22/S2_48_6  ( .A(\mult_22/ab[48][6] ), .B(
        \mult_22/CARRYB[47][6] ), .CI(\mult_22/SUMB[47][7] ), .CO(
        \mult_22/CARRYB[48][6] ), .S(\mult_22/SUMB[48][6] ) );
  FA_X1 \mult_22/S2_48_5  ( .A(\mult_22/ab[48][5] ), .B(
        \mult_22/CARRYB[47][5] ), .CI(\mult_22/SUMB[47][6] ), .CO(
        \mult_22/CARRYB[48][5] ), .S(\mult_22/SUMB[48][5] ) );
  FA_X1 \mult_22/S2_48_4  ( .A(\mult_22/ab[48][4] ), .B(
        \mult_22/CARRYB[47][4] ), .CI(\mult_22/SUMB[47][5] ), .CO(
        \mult_22/CARRYB[48][4] ), .S(\mult_22/SUMB[48][4] ) );
  FA_X1 \mult_22/S2_48_3  ( .A(\mult_22/ab[48][3] ), .B(
        \mult_22/CARRYB[47][3] ), .CI(\mult_22/SUMB[47][4] ), .CO(
        \mult_22/CARRYB[48][3] ), .S(\mult_22/SUMB[48][3] ) );
  FA_X1 \mult_22/S2_48_2  ( .A(\mult_22/ab[48][2] ), .B(
        \mult_22/CARRYB[47][2] ), .CI(\mult_22/SUMB[47][3] ), .CO(
        \mult_22/CARRYB[48][2] ), .S(\mult_22/SUMB[48][2] ) );
  FA_X1 \mult_22/S2_48_1  ( .A(\mult_22/ab[48][1] ), .B(
        \mult_22/CARRYB[47][1] ), .CI(\mult_22/SUMB[47][2] ), .CO(
        \mult_22/CARRYB[48][1] ), .S(\mult_22/SUMB[48][1] ) );
  FA_X1 \mult_22/S1_48_0  ( .A(\mult_22/ab[48][0] ), .B(
        \mult_22/CARRYB[47][0] ), .CI(\mult_22/SUMB[47][1] ), .CO(
        \mult_22/CARRYB[48][0] ), .S(N176) );
  FA_X1 \mult_22/S3_49_62  ( .A(\mult_22/ab[49][62] ), .B(
        \mult_22/CARRYB[48][62] ), .CI(\mult_22/ab[48][63] ), .CO(
        \mult_22/CARRYB[49][62] ), .S(\mult_22/SUMB[49][62] ) );
  FA_X1 \mult_22/S2_49_61  ( .A(\mult_22/ab[49][61] ), .B(
        \mult_22/CARRYB[48][61] ), .CI(\mult_22/SUMB[48][62] ), .CO(
        \mult_22/CARRYB[49][61] ), .S(\mult_22/SUMB[49][61] ) );
  FA_X1 \mult_22/S2_49_60  ( .A(\mult_22/ab[49][60] ), .B(
        \mult_22/CARRYB[48][60] ), .CI(\mult_22/SUMB[48][61] ), .CO(
        \mult_22/CARRYB[49][60] ), .S(\mult_22/SUMB[49][60] ) );
  FA_X1 \mult_22/S2_49_59  ( .A(\mult_22/ab[49][59] ), .B(
        \mult_22/CARRYB[48][59] ), .CI(\mult_22/SUMB[48][60] ), .CO(
        \mult_22/CARRYB[49][59] ), .S(\mult_22/SUMB[49][59] ) );
  FA_X1 \mult_22/S2_49_58  ( .A(\mult_22/ab[49][58] ), .B(
        \mult_22/CARRYB[48][58] ), .CI(\mult_22/SUMB[48][59] ), .CO(
        \mult_22/CARRYB[49][58] ), .S(\mult_22/SUMB[49][58] ) );
  FA_X1 \mult_22/S2_49_57  ( .A(\mult_22/ab[49][57] ), .B(
        \mult_22/CARRYB[48][57] ), .CI(\mult_22/SUMB[48][58] ), .CO(
        \mult_22/CARRYB[49][57] ), .S(\mult_22/SUMB[49][57] ) );
  FA_X1 \mult_22/S2_49_56  ( .A(\mult_22/ab[49][56] ), .B(
        \mult_22/CARRYB[48][56] ), .CI(\mult_22/SUMB[48][57] ), .CO(
        \mult_22/CARRYB[49][56] ), .S(\mult_22/SUMB[49][56] ) );
  FA_X1 \mult_22/S2_49_55  ( .A(\mult_22/ab[49][55] ), .B(
        \mult_22/CARRYB[48][55] ), .CI(\mult_22/SUMB[48][56] ), .CO(
        \mult_22/CARRYB[49][55] ), .S(\mult_22/SUMB[49][55] ) );
  FA_X1 \mult_22/S2_49_54  ( .A(\mult_22/ab[49][54] ), .B(
        \mult_22/CARRYB[48][54] ), .CI(\mult_22/SUMB[48][55] ), .CO(
        \mult_22/CARRYB[49][54] ), .S(\mult_22/SUMB[49][54] ) );
  FA_X1 \mult_22/S2_49_53  ( .A(\mult_22/ab[49][53] ), .B(
        \mult_22/CARRYB[48][53] ), .CI(\mult_22/SUMB[48][54] ), .CO(
        \mult_22/CARRYB[49][53] ), .S(\mult_22/SUMB[49][53] ) );
  FA_X1 \mult_22/S2_49_52  ( .A(\mult_22/ab[49][52] ), .B(
        \mult_22/CARRYB[48][52] ), .CI(\mult_22/SUMB[48][53] ), .CO(
        \mult_22/CARRYB[49][52] ), .S(\mult_22/SUMB[49][52] ) );
  FA_X1 \mult_22/S2_49_51  ( .A(\mult_22/ab[49][51] ), .B(
        \mult_22/CARRYB[48][51] ), .CI(\mult_22/SUMB[48][52] ), .CO(
        \mult_22/CARRYB[49][51] ), .S(\mult_22/SUMB[49][51] ) );
  FA_X1 \mult_22/S2_49_50  ( .A(\mult_22/ab[49][50] ), .B(
        \mult_22/CARRYB[48][50] ), .CI(\mult_22/SUMB[48][51] ), .CO(
        \mult_22/CARRYB[49][50] ), .S(\mult_22/SUMB[49][50] ) );
  FA_X1 \mult_22/S2_49_49  ( .A(\mult_22/ab[49][49] ), .B(
        \mult_22/CARRYB[48][49] ), .CI(\mult_22/SUMB[48][50] ), .CO(
        \mult_22/CARRYB[49][49] ), .S(\mult_22/SUMB[49][49] ) );
  FA_X1 \mult_22/S2_49_48  ( .A(\mult_22/ab[49][48] ), .B(
        \mult_22/CARRYB[48][48] ), .CI(\mult_22/SUMB[48][49] ), .CO(
        \mult_22/CARRYB[49][48] ), .S(\mult_22/SUMB[49][48] ) );
  FA_X1 \mult_22/S2_49_47  ( .A(\mult_22/ab[49][47] ), .B(
        \mult_22/CARRYB[48][47] ), .CI(\mult_22/SUMB[48][48] ), .CO(
        \mult_22/CARRYB[49][47] ), .S(\mult_22/SUMB[49][47] ) );
  FA_X1 \mult_22/S2_49_46  ( .A(\mult_22/ab[49][46] ), .B(
        \mult_22/CARRYB[48][46] ), .CI(\mult_22/SUMB[48][47] ), .CO(
        \mult_22/CARRYB[49][46] ), .S(\mult_22/SUMB[49][46] ) );
  FA_X1 \mult_22/S2_49_45  ( .A(\mult_22/ab[49][45] ), .B(
        \mult_22/CARRYB[48][45] ), .CI(\mult_22/SUMB[48][46] ), .CO(
        \mult_22/CARRYB[49][45] ), .S(\mult_22/SUMB[49][45] ) );
  FA_X1 \mult_22/S2_49_44  ( .A(\mult_22/ab[49][44] ), .B(
        \mult_22/CARRYB[48][44] ), .CI(\mult_22/SUMB[48][45] ), .CO(
        \mult_22/CARRYB[49][44] ), .S(\mult_22/SUMB[49][44] ) );
  FA_X1 \mult_22/S2_49_43  ( .A(\mult_22/ab[49][43] ), .B(
        \mult_22/CARRYB[48][43] ), .CI(\mult_22/SUMB[48][44] ), .CO(
        \mult_22/CARRYB[49][43] ), .S(\mult_22/SUMB[49][43] ) );
  FA_X1 \mult_22/S2_49_42  ( .A(\mult_22/ab[49][42] ), .B(
        \mult_22/CARRYB[48][42] ), .CI(\mult_22/SUMB[48][43] ), .CO(
        \mult_22/CARRYB[49][42] ), .S(\mult_22/SUMB[49][42] ) );
  FA_X1 \mult_22/S2_49_41  ( .A(\mult_22/ab[49][41] ), .B(
        \mult_22/CARRYB[48][41] ), .CI(\mult_22/SUMB[48][42] ), .CO(
        \mult_22/CARRYB[49][41] ), .S(\mult_22/SUMB[49][41] ) );
  FA_X1 \mult_22/S2_49_40  ( .A(\mult_22/ab[49][40] ), .B(
        \mult_22/CARRYB[48][40] ), .CI(\mult_22/SUMB[48][41] ), .CO(
        \mult_22/CARRYB[49][40] ), .S(\mult_22/SUMB[49][40] ) );
  FA_X1 \mult_22/S2_49_39  ( .A(\mult_22/ab[49][39] ), .B(
        \mult_22/CARRYB[48][39] ), .CI(\mult_22/SUMB[48][40] ), .CO(
        \mult_22/CARRYB[49][39] ), .S(\mult_22/SUMB[49][39] ) );
  FA_X1 \mult_22/S2_49_38  ( .A(\mult_22/ab[49][38] ), .B(
        \mult_22/CARRYB[48][38] ), .CI(\mult_22/SUMB[48][39] ), .CO(
        \mult_22/CARRYB[49][38] ), .S(\mult_22/SUMB[49][38] ) );
  FA_X1 \mult_22/S2_49_37  ( .A(\mult_22/ab[49][37] ), .B(
        \mult_22/CARRYB[48][37] ), .CI(\mult_22/SUMB[48][38] ), .CO(
        \mult_22/CARRYB[49][37] ), .S(\mult_22/SUMB[49][37] ) );
  FA_X1 \mult_22/S2_49_36  ( .A(\mult_22/ab[49][36] ), .B(
        \mult_22/CARRYB[48][36] ), .CI(\mult_22/SUMB[48][37] ), .CO(
        \mult_22/CARRYB[49][36] ), .S(\mult_22/SUMB[49][36] ) );
  FA_X1 \mult_22/S2_49_35  ( .A(\mult_22/ab[49][35] ), .B(
        \mult_22/CARRYB[48][35] ), .CI(\mult_22/SUMB[48][36] ), .CO(
        \mult_22/CARRYB[49][35] ), .S(\mult_22/SUMB[49][35] ) );
  FA_X1 \mult_22/S2_49_34  ( .A(\mult_22/ab[49][34] ), .B(
        \mult_22/CARRYB[48][34] ), .CI(\mult_22/SUMB[48][35] ), .CO(
        \mult_22/CARRYB[49][34] ), .S(\mult_22/SUMB[49][34] ) );
  FA_X1 \mult_22/S2_49_33  ( .A(\mult_22/ab[49][33] ), .B(
        \mult_22/CARRYB[48][33] ), .CI(\mult_22/SUMB[48][34] ), .CO(
        \mult_22/CARRYB[49][33] ), .S(\mult_22/SUMB[49][33] ) );
  FA_X1 \mult_22/S2_49_32  ( .A(\mult_22/ab[49][32] ), .B(
        \mult_22/CARRYB[48][32] ), .CI(\mult_22/SUMB[48][33] ), .CO(
        \mult_22/CARRYB[49][32] ), .S(\mult_22/SUMB[49][32] ) );
  FA_X1 \mult_22/S2_49_31  ( .A(\mult_22/ab[49][31] ), .B(
        \mult_22/CARRYB[48][31] ), .CI(\mult_22/SUMB[48][32] ), .CO(
        \mult_22/CARRYB[49][31] ), .S(\mult_22/SUMB[49][31] ) );
  FA_X1 \mult_22/S2_49_30  ( .A(\mult_22/ab[49][30] ), .B(
        \mult_22/CARRYB[48][30] ), .CI(\mult_22/SUMB[48][31] ), .CO(
        \mult_22/CARRYB[49][30] ), .S(\mult_22/SUMB[49][30] ) );
  FA_X1 \mult_22/S2_49_29  ( .A(\mult_22/ab[49][29] ), .B(
        \mult_22/CARRYB[48][29] ), .CI(\mult_22/SUMB[48][30] ), .CO(
        \mult_22/CARRYB[49][29] ), .S(\mult_22/SUMB[49][29] ) );
  FA_X1 \mult_22/S2_49_28  ( .A(\mult_22/ab[49][28] ), .B(
        \mult_22/CARRYB[48][28] ), .CI(\mult_22/SUMB[48][29] ), .CO(
        \mult_22/CARRYB[49][28] ), .S(\mult_22/SUMB[49][28] ) );
  FA_X1 \mult_22/S2_49_27  ( .A(\mult_22/ab[49][27] ), .B(
        \mult_22/CARRYB[48][27] ), .CI(\mult_22/SUMB[48][28] ), .CO(
        \mult_22/CARRYB[49][27] ), .S(\mult_22/SUMB[49][27] ) );
  FA_X1 \mult_22/S2_49_26  ( .A(\mult_22/ab[49][26] ), .B(
        \mult_22/CARRYB[48][26] ), .CI(\mult_22/SUMB[48][27] ), .CO(
        \mult_22/CARRYB[49][26] ), .S(\mult_22/SUMB[49][26] ) );
  FA_X1 \mult_22/S2_49_25  ( .A(\mult_22/ab[49][25] ), .B(
        \mult_22/CARRYB[48][25] ), .CI(\mult_22/SUMB[48][26] ), .CO(
        \mult_22/CARRYB[49][25] ), .S(\mult_22/SUMB[49][25] ) );
  FA_X1 \mult_22/S2_49_24  ( .A(\mult_22/ab[49][24] ), .B(
        \mult_22/CARRYB[48][24] ), .CI(\mult_22/SUMB[48][25] ), .CO(
        \mult_22/CARRYB[49][24] ), .S(\mult_22/SUMB[49][24] ) );
  FA_X1 \mult_22/S2_49_23  ( .A(\mult_22/ab[49][23] ), .B(
        \mult_22/CARRYB[48][23] ), .CI(\mult_22/SUMB[48][24] ), .CO(
        \mult_22/CARRYB[49][23] ), .S(\mult_22/SUMB[49][23] ) );
  FA_X1 \mult_22/S2_49_22  ( .A(\mult_22/ab[49][22] ), .B(
        \mult_22/CARRYB[48][22] ), .CI(\mult_22/SUMB[48][23] ), .CO(
        \mult_22/CARRYB[49][22] ), .S(\mult_22/SUMB[49][22] ) );
  FA_X1 \mult_22/S2_49_21  ( .A(\mult_22/ab[49][21] ), .B(
        \mult_22/CARRYB[48][21] ), .CI(\mult_22/SUMB[48][22] ), .CO(
        \mult_22/CARRYB[49][21] ), .S(\mult_22/SUMB[49][21] ) );
  FA_X1 \mult_22/S2_49_20  ( .A(\mult_22/ab[49][20] ), .B(
        \mult_22/CARRYB[48][20] ), .CI(\mult_22/SUMB[48][21] ), .CO(
        \mult_22/CARRYB[49][20] ), .S(\mult_22/SUMB[49][20] ) );
  FA_X1 \mult_22/S2_49_19  ( .A(\mult_22/ab[49][19] ), .B(
        \mult_22/CARRYB[48][19] ), .CI(\mult_22/SUMB[48][20] ), .CO(
        \mult_22/CARRYB[49][19] ), .S(\mult_22/SUMB[49][19] ) );
  FA_X1 \mult_22/S2_49_18  ( .A(\mult_22/CARRYB[48][18] ), .B(
        \mult_22/ab[49][18] ), .CI(\mult_22/SUMB[48][19] ), .CO(
        \mult_22/CARRYB[49][18] ), .S(\mult_22/SUMB[49][18] ) );
  FA_X1 \mult_22/S2_49_17  ( .A(\mult_22/CARRYB[48][17] ), .B(
        \mult_22/ab[49][17] ), .CI(\mult_22/SUMB[48][18] ), .CO(
        \mult_22/CARRYB[49][17] ), .S(\mult_22/SUMB[49][17] ) );
  FA_X1 \mult_22/S2_49_16  ( .A(\mult_22/CARRYB[48][16] ), .B(
        \mult_22/ab[49][16] ), .CI(\mult_22/SUMB[48][17] ), .CO(
        \mult_22/CARRYB[49][16] ), .S(\mult_22/SUMB[49][16] ) );
  FA_X1 \mult_22/S2_49_15  ( .A(\mult_22/ab[49][15] ), .B(
        \mult_22/CARRYB[48][15] ), .CI(\mult_22/SUMB[48][16] ), .CO(
        \mult_22/CARRYB[49][15] ), .S(\mult_22/SUMB[49][15] ) );
  FA_X1 \mult_22/S2_49_14  ( .A(\mult_22/ab[49][14] ), .B(
        \mult_22/CARRYB[48][14] ), .CI(\mult_22/SUMB[48][15] ), .CO(
        \mult_22/CARRYB[49][14] ), .S(\mult_22/SUMB[49][14] ) );
  FA_X1 \mult_22/S2_49_13  ( .A(\mult_22/CARRYB[48][13] ), .B(
        \mult_22/ab[49][13] ), .CI(\mult_22/SUMB[48][14] ), .CO(
        \mult_22/CARRYB[49][13] ), .S(\mult_22/SUMB[49][13] ) );
  FA_X1 \mult_22/S2_49_12  ( .A(\mult_22/ab[49][12] ), .B(
        \mult_22/CARRYB[48][12] ), .CI(\mult_22/SUMB[48][13] ), .CO(
        \mult_22/CARRYB[49][12] ), .S(\mult_22/SUMB[49][12] ) );
  FA_X1 \mult_22/S2_49_11  ( .A(\mult_22/ab[49][11] ), .B(
        \mult_22/CARRYB[48][11] ), .CI(\mult_22/SUMB[48][12] ), .CO(
        \mult_22/CARRYB[49][11] ), .S(\mult_22/SUMB[49][11] ) );
  FA_X1 \mult_22/S2_49_10  ( .A(\mult_22/ab[49][10] ), .B(
        \mult_22/CARRYB[48][10] ), .CI(\mult_22/SUMB[48][11] ), .CO(
        \mult_22/CARRYB[49][10] ), .S(\mult_22/SUMB[49][10] ) );
  FA_X1 \mult_22/S2_49_9  ( .A(\mult_22/ab[49][9] ), .B(
        \mult_22/CARRYB[48][9] ), .CI(\mult_22/SUMB[48][10] ), .CO(
        \mult_22/CARRYB[49][9] ), .S(\mult_22/SUMB[49][9] ) );
  FA_X1 \mult_22/S2_49_8  ( .A(\mult_22/ab[49][8] ), .B(
        \mult_22/CARRYB[48][8] ), .CI(\mult_22/SUMB[48][9] ), .CO(
        \mult_22/CARRYB[49][8] ), .S(\mult_22/SUMB[49][8] ) );
  FA_X1 \mult_22/S2_49_7  ( .A(\mult_22/ab[49][7] ), .B(
        \mult_22/CARRYB[48][7] ), .CI(\mult_22/SUMB[48][8] ), .CO(
        \mult_22/CARRYB[49][7] ), .S(\mult_22/SUMB[49][7] ) );
  FA_X1 \mult_22/S2_49_6  ( .A(\mult_22/ab[49][6] ), .B(
        \mult_22/CARRYB[48][6] ), .CI(\mult_22/SUMB[48][7] ), .CO(
        \mult_22/CARRYB[49][6] ), .S(\mult_22/SUMB[49][6] ) );
  FA_X1 \mult_22/S2_49_5  ( .A(\mult_22/ab[49][5] ), .B(
        \mult_22/CARRYB[48][5] ), .CI(\mult_22/SUMB[48][6] ), .CO(
        \mult_22/CARRYB[49][5] ), .S(\mult_22/SUMB[49][5] ) );
  FA_X1 \mult_22/S2_49_4  ( .A(\mult_22/ab[49][4] ), .B(
        \mult_22/CARRYB[48][4] ), .CI(\mult_22/SUMB[48][5] ), .CO(
        \mult_22/CARRYB[49][4] ), .S(\mult_22/SUMB[49][4] ) );
  FA_X1 \mult_22/S2_49_3  ( .A(\mult_22/ab[49][3] ), .B(
        \mult_22/CARRYB[48][3] ), .CI(\mult_22/SUMB[48][4] ), .CO(
        \mult_22/CARRYB[49][3] ), .S(\mult_22/SUMB[49][3] ) );
  FA_X1 \mult_22/S2_49_2  ( .A(\mult_22/ab[49][2] ), .B(
        \mult_22/CARRYB[48][2] ), .CI(\mult_22/SUMB[48][3] ), .CO(
        \mult_22/CARRYB[49][2] ), .S(\mult_22/SUMB[49][2] ) );
  FA_X1 \mult_22/S2_49_1  ( .A(\mult_22/ab[49][1] ), .B(
        \mult_22/CARRYB[48][1] ), .CI(\mult_22/SUMB[48][2] ), .CO(
        \mult_22/CARRYB[49][1] ), .S(\mult_22/SUMB[49][1] ) );
  FA_X1 \mult_22/S1_49_0  ( .A(\mult_22/ab[49][0] ), .B(
        \mult_22/CARRYB[48][0] ), .CI(\mult_22/SUMB[48][1] ), .CO(
        \mult_22/CARRYB[49][0] ), .S(N177) );
  FA_X1 \mult_22/S3_50_62  ( .A(\mult_22/ab[50][62] ), .B(
        \mult_22/CARRYB[49][62] ), .CI(\mult_22/ab[49][63] ), .CO(
        \mult_22/CARRYB[50][62] ), .S(\mult_22/SUMB[50][62] ) );
  FA_X1 \mult_22/S2_50_61  ( .A(\mult_22/ab[50][61] ), .B(
        \mult_22/CARRYB[49][61] ), .CI(\mult_22/SUMB[49][62] ), .CO(
        \mult_22/CARRYB[50][61] ), .S(\mult_22/SUMB[50][61] ) );
  FA_X1 \mult_22/S2_50_60  ( .A(\mult_22/ab[50][60] ), .B(
        \mult_22/CARRYB[49][60] ), .CI(\mult_22/SUMB[49][61] ), .CO(
        \mult_22/CARRYB[50][60] ), .S(\mult_22/SUMB[50][60] ) );
  FA_X1 \mult_22/S2_50_59  ( .A(\mult_22/ab[50][59] ), .B(
        \mult_22/CARRYB[49][59] ), .CI(\mult_22/SUMB[49][60] ), .CO(
        \mult_22/CARRYB[50][59] ), .S(\mult_22/SUMB[50][59] ) );
  FA_X1 \mult_22/S2_50_58  ( .A(\mult_22/ab[50][58] ), .B(
        \mult_22/CARRYB[49][58] ), .CI(\mult_22/SUMB[49][59] ), .CO(
        \mult_22/CARRYB[50][58] ), .S(\mult_22/SUMB[50][58] ) );
  FA_X1 \mult_22/S2_50_57  ( .A(\mult_22/ab[50][57] ), .B(
        \mult_22/CARRYB[49][57] ), .CI(\mult_22/SUMB[49][58] ), .CO(
        \mult_22/CARRYB[50][57] ), .S(\mult_22/SUMB[50][57] ) );
  FA_X1 \mult_22/S2_50_56  ( .A(\mult_22/ab[50][56] ), .B(
        \mult_22/CARRYB[49][56] ), .CI(\mult_22/SUMB[49][57] ), .CO(
        \mult_22/CARRYB[50][56] ), .S(\mult_22/SUMB[50][56] ) );
  FA_X1 \mult_22/S2_50_55  ( .A(\mult_22/ab[50][55] ), .B(
        \mult_22/CARRYB[49][55] ), .CI(\mult_22/SUMB[49][56] ), .CO(
        \mult_22/CARRYB[50][55] ), .S(\mult_22/SUMB[50][55] ) );
  FA_X1 \mult_22/S2_50_54  ( .A(\mult_22/ab[50][54] ), .B(
        \mult_22/CARRYB[49][54] ), .CI(\mult_22/SUMB[49][55] ), .CO(
        \mult_22/CARRYB[50][54] ), .S(\mult_22/SUMB[50][54] ) );
  FA_X1 \mult_22/S2_50_53  ( .A(\mult_22/ab[50][53] ), .B(
        \mult_22/CARRYB[49][53] ), .CI(\mult_22/SUMB[49][54] ), .CO(
        \mult_22/CARRYB[50][53] ), .S(\mult_22/SUMB[50][53] ) );
  FA_X1 \mult_22/S2_50_52  ( .A(\mult_22/ab[50][52] ), .B(
        \mult_22/CARRYB[49][52] ), .CI(\mult_22/SUMB[49][53] ), .CO(
        \mult_22/CARRYB[50][52] ), .S(\mult_22/SUMB[50][52] ) );
  FA_X1 \mult_22/S2_50_51  ( .A(\mult_22/ab[50][51] ), .B(
        \mult_22/CARRYB[49][51] ), .CI(\mult_22/SUMB[49][52] ), .CO(
        \mult_22/CARRYB[50][51] ), .S(\mult_22/SUMB[50][51] ) );
  FA_X1 \mult_22/S2_50_50  ( .A(\mult_22/ab[50][50] ), .B(
        \mult_22/CARRYB[49][50] ), .CI(\mult_22/SUMB[49][51] ), .CO(
        \mult_22/CARRYB[50][50] ), .S(\mult_22/SUMB[50][50] ) );
  FA_X1 \mult_22/S2_50_49  ( .A(\mult_22/ab[50][49] ), .B(
        \mult_22/CARRYB[49][49] ), .CI(\mult_22/SUMB[49][50] ), .CO(
        \mult_22/CARRYB[50][49] ), .S(\mult_22/SUMB[50][49] ) );
  FA_X1 \mult_22/S2_50_48  ( .A(\mult_22/ab[50][48] ), .B(
        \mult_22/CARRYB[49][48] ), .CI(\mult_22/SUMB[49][49] ), .CO(
        \mult_22/CARRYB[50][48] ), .S(\mult_22/SUMB[50][48] ) );
  FA_X1 \mult_22/S2_50_47  ( .A(\mult_22/ab[50][47] ), .B(
        \mult_22/CARRYB[49][47] ), .CI(\mult_22/SUMB[49][48] ), .CO(
        \mult_22/CARRYB[50][47] ), .S(\mult_22/SUMB[50][47] ) );
  FA_X1 \mult_22/S2_50_46  ( .A(\mult_22/ab[50][46] ), .B(
        \mult_22/CARRYB[49][46] ), .CI(\mult_22/SUMB[49][47] ), .CO(
        \mult_22/CARRYB[50][46] ), .S(\mult_22/SUMB[50][46] ) );
  FA_X1 \mult_22/S2_50_45  ( .A(\mult_22/ab[50][45] ), .B(
        \mult_22/CARRYB[49][45] ), .CI(\mult_22/SUMB[49][46] ), .CO(
        \mult_22/CARRYB[50][45] ), .S(\mult_22/SUMB[50][45] ) );
  FA_X1 \mult_22/S2_50_44  ( .A(\mult_22/ab[50][44] ), .B(
        \mult_22/CARRYB[49][44] ), .CI(\mult_22/SUMB[49][45] ), .CO(
        \mult_22/CARRYB[50][44] ), .S(\mult_22/SUMB[50][44] ) );
  FA_X1 \mult_22/S2_50_43  ( .A(\mult_22/ab[50][43] ), .B(
        \mult_22/CARRYB[49][43] ), .CI(\mult_22/SUMB[49][44] ), .CO(
        \mult_22/CARRYB[50][43] ), .S(\mult_22/SUMB[50][43] ) );
  FA_X1 \mult_22/S2_50_42  ( .A(\mult_22/ab[50][42] ), .B(
        \mult_22/CARRYB[49][42] ), .CI(\mult_22/SUMB[49][43] ), .CO(
        \mult_22/CARRYB[50][42] ), .S(\mult_22/SUMB[50][42] ) );
  FA_X1 \mult_22/S2_50_41  ( .A(\mult_22/ab[50][41] ), .B(
        \mult_22/CARRYB[49][41] ), .CI(\mult_22/SUMB[49][42] ), .CO(
        \mult_22/CARRYB[50][41] ), .S(\mult_22/SUMB[50][41] ) );
  FA_X1 \mult_22/S2_50_40  ( .A(\mult_22/ab[50][40] ), .B(
        \mult_22/CARRYB[49][40] ), .CI(\mult_22/SUMB[49][41] ), .CO(
        \mult_22/CARRYB[50][40] ), .S(\mult_22/SUMB[50][40] ) );
  FA_X1 \mult_22/S2_50_39  ( .A(\mult_22/ab[50][39] ), .B(
        \mult_22/CARRYB[49][39] ), .CI(\mult_22/SUMB[49][40] ), .CO(
        \mult_22/CARRYB[50][39] ), .S(\mult_22/SUMB[50][39] ) );
  FA_X1 \mult_22/S2_50_38  ( .A(\mult_22/ab[50][38] ), .B(
        \mult_22/CARRYB[49][38] ), .CI(\mult_22/SUMB[49][39] ), .CO(
        \mult_22/CARRYB[50][38] ), .S(\mult_22/SUMB[50][38] ) );
  FA_X1 \mult_22/S2_50_37  ( .A(\mult_22/ab[50][37] ), .B(
        \mult_22/CARRYB[49][37] ), .CI(\mult_22/SUMB[49][38] ), .CO(
        \mult_22/CARRYB[50][37] ), .S(\mult_22/SUMB[50][37] ) );
  FA_X1 \mult_22/S2_50_36  ( .A(\mult_22/ab[50][36] ), .B(
        \mult_22/CARRYB[49][36] ), .CI(\mult_22/SUMB[49][37] ), .CO(
        \mult_22/CARRYB[50][36] ), .S(\mult_22/SUMB[50][36] ) );
  FA_X1 \mult_22/S2_50_35  ( .A(\mult_22/ab[50][35] ), .B(
        \mult_22/CARRYB[49][35] ), .CI(\mult_22/SUMB[49][36] ), .CO(
        \mult_22/CARRYB[50][35] ), .S(\mult_22/SUMB[50][35] ) );
  FA_X1 \mult_22/S2_50_34  ( .A(\mult_22/ab[50][34] ), .B(
        \mult_22/CARRYB[49][34] ), .CI(\mult_22/SUMB[49][35] ), .CO(
        \mult_22/CARRYB[50][34] ), .S(\mult_22/SUMB[50][34] ) );
  FA_X1 \mult_22/S2_50_33  ( .A(\mult_22/ab[50][33] ), .B(
        \mult_22/CARRYB[49][33] ), .CI(\mult_22/SUMB[49][34] ), .CO(
        \mult_22/CARRYB[50][33] ), .S(\mult_22/SUMB[50][33] ) );
  FA_X1 \mult_22/S2_50_32  ( .A(\mult_22/ab[50][32] ), .B(
        \mult_22/CARRYB[49][32] ), .CI(\mult_22/SUMB[49][33] ), .CO(
        \mult_22/CARRYB[50][32] ), .S(\mult_22/SUMB[50][32] ) );
  FA_X1 \mult_22/S2_50_31  ( .A(\mult_22/ab[50][31] ), .B(
        \mult_22/CARRYB[49][31] ), .CI(\mult_22/SUMB[49][32] ), .CO(
        \mult_22/CARRYB[50][31] ), .S(\mult_22/SUMB[50][31] ) );
  FA_X1 \mult_22/S2_50_30  ( .A(\mult_22/ab[50][30] ), .B(
        \mult_22/CARRYB[49][30] ), .CI(\mult_22/SUMB[49][31] ), .CO(
        \mult_22/CARRYB[50][30] ), .S(\mult_22/SUMB[50][30] ) );
  FA_X1 \mult_22/S2_50_29  ( .A(\mult_22/ab[50][29] ), .B(
        \mult_22/CARRYB[49][29] ), .CI(\mult_22/SUMB[49][30] ), .CO(
        \mult_22/CARRYB[50][29] ), .S(\mult_22/SUMB[50][29] ) );
  FA_X1 \mult_22/S2_50_28  ( .A(\mult_22/ab[50][28] ), .B(
        \mult_22/CARRYB[49][28] ), .CI(\mult_22/SUMB[49][29] ), .CO(
        \mult_22/CARRYB[50][28] ), .S(\mult_22/SUMB[50][28] ) );
  FA_X1 \mult_22/S2_50_27  ( .A(\mult_22/ab[50][27] ), .B(
        \mult_22/CARRYB[49][27] ), .CI(\mult_22/SUMB[49][28] ), .CO(
        \mult_22/CARRYB[50][27] ), .S(\mult_22/SUMB[50][27] ) );
  FA_X1 \mult_22/S2_50_26  ( .A(\mult_22/ab[50][26] ), .B(
        \mult_22/CARRYB[49][26] ), .CI(\mult_22/SUMB[49][27] ), .CO(
        \mult_22/CARRYB[50][26] ), .S(\mult_22/SUMB[50][26] ) );
  FA_X1 \mult_22/S2_50_25  ( .A(\mult_22/ab[50][25] ), .B(
        \mult_22/CARRYB[49][25] ), .CI(\mult_22/SUMB[49][26] ), .CO(
        \mult_22/CARRYB[50][25] ), .S(\mult_22/SUMB[50][25] ) );
  FA_X1 \mult_22/S2_50_24  ( .A(\mult_22/ab[50][24] ), .B(
        \mult_22/CARRYB[49][24] ), .CI(\mult_22/SUMB[49][25] ), .CO(
        \mult_22/CARRYB[50][24] ), .S(\mult_22/SUMB[50][24] ) );
  FA_X1 \mult_22/S2_50_23  ( .A(\mult_22/ab[50][23] ), .B(
        \mult_22/CARRYB[49][23] ), .CI(\mult_22/SUMB[49][24] ), .CO(
        \mult_22/CARRYB[50][23] ), .S(\mult_22/SUMB[50][23] ) );
  FA_X1 \mult_22/S2_50_22  ( .A(\mult_22/ab[50][22] ), .B(
        \mult_22/CARRYB[49][22] ), .CI(\mult_22/SUMB[49][23] ), .CO(
        \mult_22/CARRYB[50][22] ), .S(\mult_22/SUMB[50][22] ) );
  FA_X1 \mult_22/S2_50_21  ( .A(\mult_22/ab[50][21] ), .B(
        \mult_22/CARRYB[49][21] ), .CI(\mult_22/SUMB[49][22] ), .CO(
        \mult_22/CARRYB[50][21] ), .S(\mult_22/SUMB[50][21] ) );
  FA_X1 \mult_22/S2_50_20  ( .A(\mult_22/ab[50][20] ), .B(
        \mult_22/CARRYB[49][20] ), .CI(\mult_22/SUMB[49][21] ), .CO(
        \mult_22/CARRYB[50][20] ), .S(\mult_22/SUMB[50][20] ) );
  FA_X1 \mult_22/S2_50_19  ( .A(\mult_22/ab[50][19] ), .B(
        \mult_22/CARRYB[49][19] ), .CI(\mult_22/SUMB[49][20] ), .CO(
        \mult_22/CARRYB[50][19] ), .S(\mult_22/SUMB[50][19] ) );
  FA_X1 \mult_22/S2_50_18  ( .A(\mult_22/ab[50][18] ), .B(
        \mult_22/CARRYB[49][18] ), .CI(\mult_22/SUMB[49][19] ), .CO(
        \mult_22/CARRYB[50][18] ), .S(\mult_22/SUMB[50][18] ) );
  FA_X1 \mult_22/S2_50_17  ( .A(\mult_22/ab[50][17] ), .B(
        \mult_22/CARRYB[49][17] ), .CI(\mult_22/SUMB[49][18] ), .CO(
        \mult_22/CARRYB[50][17] ), .S(\mult_22/SUMB[50][17] ) );
  FA_X1 \mult_22/S2_50_16  ( .A(\mult_22/ab[50][16] ), .B(
        \mult_22/CARRYB[49][16] ), .CI(\mult_22/SUMB[49][17] ), .CO(
        \mult_22/CARRYB[50][16] ), .S(\mult_22/SUMB[50][16] ) );
  FA_X1 \mult_22/S2_50_15  ( .A(\mult_22/CARRYB[49][15] ), .B(
        \mult_22/ab[50][15] ), .CI(\mult_22/SUMB[49][16] ), .CO(
        \mult_22/CARRYB[50][15] ), .S(\mult_22/SUMB[50][15] ) );
  FA_X1 \mult_22/S2_50_14  ( .A(\mult_22/CARRYB[49][14] ), .B(
        \mult_22/ab[50][14] ), .CI(\mult_22/SUMB[49][15] ), .CO(
        \mult_22/CARRYB[50][14] ), .S(\mult_22/SUMB[50][14] ) );
  FA_X1 \mult_22/S2_50_13  ( .A(\mult_22/ab[50][13] ), .B(
        \mult_22/CARRYB[49][13] ), .CI(\mult_22/SUMB[49][14] ), .CO(
        \mult_22/CARRYB[50][13] ), .S(\mult_22/SUMB[50][13] ) );
  FA_X1 \mult_22/S2_50_12  ( .A(\mult_22/ab[50][12] ), .B(
        \mult_22/CARRYB[49][12] ), .CI(\mult_22/SUMB[49][13] ), .CO(
        \mult_22/CARRYB[50][12] ), .S(\mult_22/SUMB[50][12] ) );
  FA_X1 \mult_22/S2_50_11  ( .A(\mult_22/ab[50][11] ), .B(
        \mult_22/CARRYB[49][11] ), .CI(\mult_22/SUMB[49][12] ), .CO(
        \mult_22/CARRYB[50][11] ), .S(\mult_22/SUMB[50][11] ) );
  FA_X1 \mult_22/S2_50_10  ( .A(\mult_22/ab[50][10] ), .B(
        \mult_22/CARRYB[49][10] ), .CI(\mult_22/SUMB[49][11] ), .CO(
        \mult_22/CARRYB[50][10] ), .S(\mult_22/SUMB[50][10] ) );
  FA_X1 \mult_22/S2_50_9  ( .A(\mult_22/ab[50][9] ), .B(
        \mult_22/CARRYB[49][9] ), .CI(\mult_22/SUMB[49][10] ), .CO(
        \mult_22/CARRYB[50][9] ), .S(\mult_22/SUMB[50][9] ) );
  FA_X1 \mult_22/S2_50_8  ( .A(\mult_22/ab[50][8] ), .B(
        \mult_22/CARRYB[49][8] ), .CI(\mult_22/SUMB[49][9] ), .CO(
        \mult_22/CARRYB[50][8] ), .S(\mult_22/SUMB[50][8] ) );
  FA_X1 \mult_22/S2_50_7  ( .A(\mult_22/ab[50][7] ), .B(
        \mult_22/CARRYB[49][7] ), .CI(\mult_22/SUMB[49][8] ), .CO(
        \mult_22/CARRYB[50][7] ), .S(\mult_22/SUMB[50][7] ) );
  FA_X1 \mult_22/S2_50_6  ( .A(\mult_22/ab[50][6] ), .B(
        \mult_22/CARRYB[49][6] ), .CI(\mult_22/SUMB[49][7] ), .CO(
        \mult_22/CARRYB[50][6] ), .S(\mult_22/SUMB[50][6] ) );
  FA_X1 \mult_22/S2_50_5  ( .A(\mult_22/ab[50][5] ), .B(
        \mult_22/CARRYB[49][5] ), .CI(\mult_22/SUMB[49][6] ), .CO(
        \mult_22/CARRYB[50][5] ), .S(\mult_22/SUMB[50][5] ) );
  FA_X1 \mult_22/S2_50_4  ( .A(\mult_22/ab[50][4] ), .B(
        \mult_22/CARRYB[49][4] ), .CI(\mult_22/SUMB[49][5] ), .CO(
        \mult_22/CARRYB[50][4] ), .S(\mult_22/SUMB[50][4] ) );
  FA_X1 \mult_22/S2_50_3  ( .A(\mult_22/ab[50][3] ), .B(
        \mult_22/CARRYB[49][3] ), .CI(\mult_22/SUMB[49][4] ), .CO(
        \mult_22/CARRYB[50][3] ), .S(\mult_22/SUMB[50][3] ) );
  FA_X1 \mult_22/S2_50_2  ( .A(\mult_22/ab[50][2] ), .B(
        \mult_22/CARRYB[49][2] ), .CI(\mult_22/SUMB[49][3] ), .CO(
        \mult_22/CARRYB[50][2] ), .S(\mult_22/SUMB[50][2] ) );
  FA_X1 \mult_22/S2_50_1  ( .A(\mult_22/ab[50][1] ), .B(
        \mult_22/CARRYB[49][1] ), .CI(\mult_22/SUMB[49][2] ), .CO(
        \mult_22/CARRYB[50][1] ), .S(\mult_22/SUMB[50][1] ) );
  FA_X1 \mult_22/S1_50_0  ( .A(\mult_22/ab[50][0] ), .B(
        \mult_22/CARRYB[49][0] ), .CI(\mult_22/SUMB[49][1] ), .CO(
        \mult_22/CARRYB[50][0] ), .S(N178) );
  FA_X1 \mult_22/S3_51_62  ( .A(\mult_22/ab[51][62] ), .B(
        \mult_22/CARRYB[50][62] ), .CI(\mult_22/ab[50][63] ), .CO(
        \mult_22/CARRYB[51][62] ), .S(\mult_22/SUMB[51][62] ) );
  FA_X1 \mult_22/S2_51_61  ( .A(\mult_22/ab[51][61] ), .B(
        \mult_22/CARRYB[50][61] ), .CI(\mult_22/SUMB[50][62] ), .CO(
        \mult_22/CARRYB[51][61] ), .S(\mult_22/SUMB[51][61] ) );
  FA_X1 \mult_22/S2_51_60  ( .A(\mult_22/ab[51][60] ), .B(
        \mult_22/CARRYB[50][60] ), .CI(\mult_22/SUMB[50][61] ), .CO(
        \mult_22/CARRYB[51][60] ), .S(\mult_22/SUMB[51][60] ) );
  FA_X1 \mult_22/S2_51_59  ( .A(\mult_22/ab[51][59] ), .B(
        \mult_22/CARRYB[50][59] ), .CI(\mult_22/SUMB[50][60] ), .CO(
        \mult_22/CARRYB[51][59] ), .S(\mult_22/SUMB[51][59] ) );
  FA_X1 \mult_22/S2_51_58  ( .A(\mult_22/ab[51][58] ), .B(
        \mult_22/CARRYB[50][58] ), .CI(\mult_22/SUMB[50][59] ), .CO(
        \mult_22/CARRYB[51][58] ), .S(\mult_22/SUMB[51][58] ) );
  FA_X1 \mult_22/S2_51_57  ( .A(\mult_22/ab[51][57] ), .B(
        \mult_22/CARRYB[50][57] ), .CI(\mult_22/SUMB[50][58] ), .CO(
        \mult_22/CARRYB[51][57] ), .S(\mult_22/SUMB[51][57] ) );
  FA_X1 \mult_22/S2_51_56  ( .A(\mult_22/ab[51][56] ), .B(
        \mult_22/CARRYB[50][56] ), .CI(\mult_22/SUMB[50][57] ), .CO(
        \mult_22/CARRYB[51][56] ), .S(\mult_22/SUMB[51][56] ) );
  FA_X1 \mult_22/S2_51_55  ( .A(\mult_22/ab[51][55] ), .B(
        \mult_22/CARRYB[50][55] ), .CI(\mult_22/SUMB[50][56] ), .CO(
        \mult_22/CARRYB[51][55] ), .S(\mult_22/SUMB[51][55] ) );
  FA_X1 \mult_22/S2_51_54  ( .A(\mult_22/ab[51][54] ), .B(
        \mult_22/CARRYB[50][54] ), .CI(\mult_22/SUMB[50][55] ), .CO(
        \mult_22/CARRYB[51][54] ), .S(\mult_22/SUMB[51][54] ) );
  FA_X1 \mult_22/S2_51_53  ( .A(\mult_22/ab[51][53] ), .B(
        \mult_22/CARRYB[50][53] ), .CI(\mult_22/SUMB[50][54] ), .CO(
        \mult_22/CARRYB[51][53] ), .S(\mult_22/SUMB[51][53] ) );
  FA_X1 \mult_22/S2_51_52  ( .A(\mult_22/ab[51][52] ), .B(
        \mult_22/CARRYB[50][52] ), .CI(\mult_22/SUMB[50][53] ), .CO(
        \mult_22/CARRYB[51][52] ), .S(\mult_22/SUMB[51][52] ) );
  FA_X1 \mult_22/S2_51_51  ( .A(\mult_22/ab[51][51] ), .B(
        \mult_22/CARRYB[50][51] ), .CI(\mult_22/SUMB[50][52] ), .CO(
        \mult_22/CARRYB[51][51] ), .S(\mult_22/SUMB[51][51] ) );
  FA_X1 \mult_22/S2_51_50  ( .A(\mult_22/ab[51][50] ), .B(
        \mult_22/CARRYB[50][50] ), .CI(\mult_22/SUMB[50][51] ), .CO(
        \mult_22/CARRYB[51][50] ), .S(\mult_22/SUMB[51][50] ) );
  FA_X1 \mult_22/S2_51_49  ( .A(\mult_22/ab[51][49] ), .B(
        \mult_22/CARRYB[50][49] ), .CI(\mult_22/SUMB[50][50] ), .CO(
        \mult_22/CARRYB[51][49] ), .S(\mult_22/SUMB[51][49] ) );
  FA_X1 \mult_22/S2_51_48  ( .A(\mult_22/ab[51][48] ), .B(
        \mult_22/CARRYB[50][48] ), .CI(\mult_22/SUMB[50][49] ), .CO(
        \mult_22/CARRYB[51][48] ), .S(\mult_22/SUMB[51][48] ) );
  FA_X1 \mult_22/S2_51_47  ( .A(\mult_22/ab[51][47] ), .B(
        \mult_22/CARRYB[50][47] ), .CI(\mult_22/SUMB[50][48] ), .CO(
        \mult_22/CARRYB[51][47] ), .S(\mult_22/SUMB[51][47] ) );
  FA_X1 \mult_22/S2_51_46  ( .A(\mult_22/ab[51][46] ), .B(
        \mult_22/CARRYB[50][46] ), .CI(\mult_22/SUMB[50][47] ), .CO(
        \mult_22/CARRYB[51][46] ), .S(\mult_22/SUMB[51][46] ) );
  FA_X1 \mult_22/S2_51_45  ( .A(\mult_22/ab[51][45] ), .B(
        \mult_22/CARRYB[50][45] ), .CI(\mult_22/SUMB[50][46] ), .CO(
        \mult_22/CARRYB[51][45] ), .S(\mult_22/SUMB[51][45] ) );
  FA_X1 \mult_22/S2_51_44  ( .A(\mult_22/ab[51][44] ), .B(
        \mult_22/CARRYB[50][44] ), .CI(\mult_22/SUMB[50][45] ), .CO(
        \mult_22/CARRYB[51][44] ), .S(\mult_22/SUMB[51][44] ) );
  FA_X1 \mult_22/S2_51_43  ( .A(\mult_22/ab[51][43] ), .B(
        \mult_22/CARRYB[50][43] ), .CI(\mult_22/SUMB[50][44] ), .CO(
        \mult_22/CARRYB[51][43] ), .S(\mult_22/SUMB[51][43] ) );
  FA_X1 \mult_22/S2_51_42  ( .A(\mult_22/ab[51][42] ), .B(
        \mult_22/CARRYB[50][42] ), .CI(\mult_22/SUMB[50][43] ), .CO(
        \mult_22/CARRYB[51][42] ), .S(\mult_22/SUMB[51][42] ) );
  FA_X1 \mult_22/S2_51_41  ( .A(\mult_22/ab[51][41] ), .B(
        \mult_22/CARRYB[50][41] ), .CI(\mult_22/SUMB[50][42] ), .CO(
        \mult_22/CARRYB[51][41] ), .S(\mult_22/SUMB[51][41] ) );
  FA_X1 \mult_22/S2_51_40  ( .A(\mult_22/ab[51][40] ), .B(
        \mult_22/CARRYB[50][40] ), .CI(\mult_22/SUMB[50][41] ), .CO(
        \mult_22/CARRYB[51][40] ), .S(\mult_22/SUMB[51][40] ) );
  FA_X1 \mult_22/S2_51_39  ( .A(\mult_22/ab[51][39] ), .B(
        \mult_22/CARRYB[50][39] ), .CI(\mult_22/SUMB[50][40] ), .CO(
        \mult_22/CARRYB[51][39] ), .S(\mult_22/SUMB[51][39] ) );
  FA_X1 \mult_22/S2_51_38  ( .A(\mult_22/ab[51][38] ), .B(
        \mult_22/CARRYB[50][38] ), .CI(\mult_22/SUMB[50][39] ), .CO(
        \mult_22/CARRYB[51][38] ), .S(\mult_22/SUMB[51][38] ) );
  FA_X1 \mult_22/S2_51_37  ( .A(\mult_22/ab[51][37] ), .B(
        \mult_22/CARRYB[50][37] ), .CI(\mult_22/SUMB[50][38] ), .CO(
        \mult_22/CARRYB[51][37] ), .S(\mult_22/SUMB[51][37] ) );
  FA_X1 \mult_22/S2_51_36  ( .A(\mult_22/ab[51][36] ), .B(
        \mult_22/CARRYB[50][36] ), .CI(\mult_22/SUMB[50][37] ), .CO(
        \mult_22/CARRYB[51][36] ), .S(\mult_22/SUMB[51][36] ) );
  FA_X1 \mult_22/S2_51_35  ( .A(\mult_22/ab[51][35] ), .B(
        \mult_22/CARRYB[50][35] ), .CI(\mult_22/SUMB[50][36] ), .CO(
        \mult_22/CARRYB[51][35] ), .S(\mult_22/SUMB[51][35] ) );
  FA_X1 \mult_22/S2_51_34  ( .A(\mult_22/ab[51][34] ), .B(
        \mult_22/CARRYB[50][34] ), .CI(\mult_22/SUMB[50][35] ), .CO(
        \mult_22/CARRYB[51][34] ), .S(\mult_22/SUMB[51][34] ) );
  FA_X1 \mult_22/S2_51_33  ( .A(\mult_22/ab[51][33] ), .B(
        \mult_22/CARRYB[50][33] ), .CI(\mult_22/SUMB[50][34] ), .CO(
        \mult_22/CARRYB[51][33] ), .S(\mult_22/SUMB[51][33] ) );
  FA_X1 \mult_22/S2_51_32  ( .A(\mult_22/ab[51][32] ), .B(
        \mult_22/CARRYB[50][32] ), .CI(\mult_22/SUMB[50][33] ), .CO(
        \mult_22/CARRYB[51][32] ), .S(\mult_22/SUMB[51][32] ) );
  FA_X1 \mult_22/S2_51_31  ( .A(\mult_22/ab[51][31] ), .B(
        \mult_22/CARRYB[50][31] ), .CI(\mult_22/SUMB[50][32] ), .CO(
        \mult_22/CARRYB[51][31] ), .S(\mult_22/SUMB[51][31] ) );
  FA_X1 \mult_22/S2_51_30  ( .A(\mult_22/ab[51][30] ), .B(
        \mult_22/CARRYB[50][30] ), .CI(\mult_22/SUMB[50][31] ), .CO(
        \mult_22/CARRYB[51][30] ), .S(\mult_22/SUMB[51][30] ) );
  FA_X1 \mult_22/S2_51_29  ( .A(\mult_22/ab[51][29] ), .B(
        \mult_22/CARRYB[50][29] ), .CI(\mult_22/SUMB[50][30] ), .CO(
        \mult_22/CARRYB[51][29] ), .S(\mult_22/SUMB[51][29] ) );
  FA_X1 \mult_22/S2_51_28  ( .A(\mult_22/ab[51][28] ), .B(
        \mult_22/CARRYB[50][28] ), .CI(\mult_22/SUMB[50][29] ), .CO(
        \mult_22/CARRYB[51][28] ), .S(\mult_22/SUMB[51][28] ) );
  FA_X1 \mult_22/S2_51_27  ( .A(\mult_22/ab[51][27] ), .B(
        \mult_22/CARRYB[50][27] ), .CI(\mult_22/SUMB[50][28] ), .CO(
        \mult_22/CARRYB[51][27] ), .S(\mult_22/SUMB[51][27] ) );
  FA_X1 \mult_22/S2_51_26  ( .A(\mult_22/ab[51][26] ), .B(
        \mult_22/CARRYB[50][26] ), .CI(\mult_22/SUMB[50][27] ), .CO(
        \mult_22/CARRYB[51][26] ), .S(\mult_22/SUMB[51][26] ) );
  FA_X1 \mult_22/S2_51_25  ( .A(\mult_22/ab[51][25] ), .B(
        \mult_22/CARRYB[50][25] ), .CI(\mult_22/SUMB[50][26] ), .CO(
        \mult_22/CARRYB[51][25] ), .S(\mult_22/SUMB[51][25] ) );
  FA_X1 \mult_22/S2_51_24  ( .A(\mult_22/ab[51][24] ), .B(
        \mult_22/CARRYB[50][24] ), .CI(\mult_22/SUMB[50][25] ), .CO(
        \mult_22/CARRYB[51][24] ), .S(\mult_22/SUMB[51][24] ) );
  FA_X1 \mult_22/S2_51_23  ( .A(\mult_22/ab[51][23] ), .B(
        \mult_22/CARRYB[50][23] ), .CI(\mult_22/SUMB[50][24] ), .CO(
        \mult_22/CARRYB[51][23] ), .S(\mult_22/SUMB[51][23] ) );
  FA_X1 \mult_22/S2_51_22  ( .A(\mult_22/ab[51][22] ), .B(
        \mult_22/CARRYB[50][22] ), .CI(\mult_22/SUMB[50][23] ), .CO(
        \mult_22/CARRYB[51][22] ), .S(\mult_22/SUMB[51][22] ) );
  FA_X1 \mult_22/S2_51_21  ( .A(\mult_22/ab[51][21] ), .B(
        \mult_22/CARRYB[50][21] ), .CI(\mult_22/SUMB[50][22] ), .CO(
        \mult_22/CARRYB[51][21] ), .S(\mult_22/SUMB[51][21] ) );
  FA_X1 \mult_22/S2_51_20  ( .A(\mult_22/ab[51][20] ), .B(
        \mult_22/CARRYB[50][20] ), .CI(\mult_22/SUMB[50][21] ), .CO(
        \mult_22/CARRYB[51][20] ), .S(\mult_22/SUMB[51][20] ) );
  FA_X1 \mult_22/S2_51_19  ( .A(\mult_22/ab[51][19] ), .B(
        \mult_22/CARRYB[50][19] ), .CI(\mult_22/SUMB[50][20] ), .CO(
        \mult_22/CARRYB[51][19] ), .S(\mult_22/SUMB[51][19] ) );
  FA_X1 \mult_22/S2_51_18  ( .A(\mult_22/ab[51][18] ), .B(
        \mult_22/CARRYB[50][18] ), .CI(\mult_22/SUMB[50][19] ), .CO(
        \mult_22/CARRYB[51][18] ), .S(\mult_22/SUMB[51][18] ) );
  FA_X1 \mult_22/S2_51_17  ( .A(\mult_22/ab[51][17] ), .B(
        \mult_22/CARRYB[50][17] ), .CI(\mult_22/SUMB[50][18] ), .CO(
        \mult_22/CARRYB[51][17] ), .S(\mult_22/SUMB[51][17] ) );
  FA_X1 \mult_22/S2_51_16  ( .A(\mult_22/CARRYB[50][16] ), .B(
        \mult_22/ab[51][16] ), .CI(\mult_22/SUMB[50][17] ), .CO(
        \mult_22/CARRYB[51][16] ), .S(\mult_22/SUMB[51][16] ) );
  FA_X1 \mult_22/S2_51_15  ( .A(\mult_22/CARRYB[50][15] ), .B(
        \mult_22/ab[51][15] ), .CI(\mult_22/SUMB[50][16] ), .CO(
        \mult_22/CARRYB[51][15] ), .S(\mult_22/SUMB[51][15] ) );
  FA_X1 \mult_22/S2_51_14  ( .A(\mult_22/ab[51][14] ), .B(
        \mult_22/CARRYB[50][14] ), .CI(\mult_22/SUMB[50][15] ), .CO(
        \mult_22/CARRYB[51][14] ), .S(\mult_22/SUMB[51][14] ) );
  FA_X1 \mult_22/S2_51_13  ( .A(\mult_22/ab[51][13] ), .B(
        \mult_22/CARRYB[50][13] ), .CI(\mult_22/SUMB[50][14] ), .CO(
        \mult_22/CARRYB[51][13] ), .S(\mult_22/SUMB[51][13] ) );
  FA_X1 \mult_22/S2_51_12  ( .A(\mult_22/ab[51][12] ), .B(
        \mult_22/CARRYB[50][12] ), .CI(\mult_22/SUMB[50][13] ), .CO(
        \mult_22/CARRYB[51][12] ), .S(\mult_22/SUMB[51][12] ) );
  FA_X1 \mult_22/S2_51_11  ( .A(\mult_22/ab[51][11] ), .B(
        \mult_22/CARRYB[50][11] ), .CI(\mult_22/SUMB[50][12] ), .CO(
        \mult_22/CARRYB[51][11] ), .S(\mult_22/SUMB[51][11] ) );
  FA_X1 \mult_22/S2_51_10  ( .A(\mult_22/ab[51][10] ), .B(
        \mult_22/CARRYB[50][10] ), .CI(\mult_22/SUMB[50][11] ), .CO(
        \mult_22/CARRYB[51][10] ), .S(\mult_22/SUMB[51][10] ) );
  FA_X1 \mult_22/S2_51_9  ( .A(\mult_22/ab[51][9] ), .B(
        \mult_22/CARRYB[50][9] ), .CI(\mult_22/SUMB[50][10] ), .CO(
        \mult_22/CARRYB[51][9] ), .S(\mult_22/SUMB[51][9] ) );
  FA_X1 \mult_22/S2_51_8  ( .A(\mult_22/ab[51][8] ), .B(
        \mult_22/CARRYB[50][8] ), .CI(\mult_22/SUMB[50][9] ), .CO(
        \mult_22/CARRYB[51][8] ), .S(\mult_22/SUMB[51][8] ) );
  FA_X1 \mult_22/S2_51_7  ( .A(\mult_22/ab[51][7] ), .B(
        \mult_22/CARRYB[50][7] ), .CI(\mult_22/SUMB[50][8] ), .CO(
        \mult_22/CARRYB[51][7] ), .S(\mult_22/SUMB[51][7] ) );
  FA_X1 \mult_22/S2_51_6  ( .A(\mult_22/ab[51][6] ), .B(
        \mult_22/CARRYB[50][6] ), .CI(\mult_22/SUMB[50][7] ), .CO(
        \mult_22/CARRYB[51][6] ), .S(\mult_22/SUMB[51][6] ) );
  FA_X1 \mult_22/S2_51_5  ( .A(\mult_22/ab[51][5] ), .B(
        \mult_22/CARRYB[50][5] ), .CI(\mult_22/SUMB[50][6] ), .CO(
        \mult_22/CARRYB[51][5] ), .S(\mult_22/SUMB[51][5] ) );
  FA_X1 \mult_22/S2_51_4  ( .A(\mult_22/ab[51][4] ), .B(
        \mult_22/CARRYB[50][4] ), .CI(\mult_22/SUMB[50][5] ), .CO(
        \mult_22/CARRYB[51][4] ), .S(\mult_22/SUMB[51][4] ) );
  FA_X1 \mult_22/S2_51_3  ( .A(\mult_22/ab[51][3] ), .B(
        \mult_22/CARRYB[50][3] ), .CI(\mult_22/SUMB[50][4] ), .CO(
        \mult_22/CARRYB[51][3] ), .S(\mult_22/SUMB[51][3] ) );
  FA_X1 \mult_22/S2_51_2  ( .A(\mult_22/ab[51][2] ), .B(
        \mult_22/CARRYB[50][2] ), .CI(\mult_22/SUMB[50][3] ), .CO(
        \mult_22/CARRYB[51][2] ), .S(\mult_22/SUMB[51][2] ) );
  FA_X1 \mult_22/S2_51_1  ( .A(\mult_22/ab[51][1] ), .B(
        \mult_22/CARRYB[50][1] ), .CI(\mult_22/SUMB[50][2] ), .CO(
        \mult_22/CARRYB[51][1] ), .S(\mult_22/SUMB[51][1] ) );
  FA_X1 \mult_22/S1_51_0  ( .A(\mult_22/ab[51][0] ), .B(
        \mult_22/CARRYB[50][0] ), .CI(\mult_22/SUMB[50][1] ), .CO(
        \mult_22/CARRYB[51][0] ), .S(N179) );
  FA_X1 \mult_22/S3_52_62  ( .A(\mult_22/ab[52][62] ), .B(
        \mult_22/CARRYB[51][62] ), .CI(\mult_22/ab[51][63] ), .CO(
        \mult_22/CARRYB[52][62] ), .S(\mult_22/SUMB[52][62] ) );
  FA_X1 \mult_22/S2_52_61  ( .A(\mult_22/ab[52][61] ), .B(
        \mult_22/CARRYB[51][61] ), .CI(\mult_22/SUMB[51][62] ), .CO(
        \mult_22/CARRYB[52][61] ), .S(\mult_22/SUMB[52][61] ) );
  FA_X1 \mult_22/S2_52_60  ( .A(\mult_22/ab[52][60] ), .B(
        \mult_22/CARRYB[51][60] ), .CI(\mult_22/SUMB[51][61] ), .CO(
        \mult_22/CARRYB[52][60] ), .S(\mult_22/SUMB[52][60] ) );
  FA_X1 \mult_22/S2_52_59  ( .A(\mult_22/ab[52][59] ), .B(
        \mult_22/CARRYB[51][59] ), .CI(\mult_22/SUMB[51][60] ), .CO(
        \mult_22/CARRYB[52][59] ), .S(\mult_22/SUMB[52][59] ) );
  FA_X1 \mult_22/S2_52_58  ( .A(\mult_22/ab[52][58] ), .B(
        \mult_22/CARRYB[51][58] ), .CI(\mult_22/SUMB[51][59] ), .CO(
        \mult_22/CARRYB[52][58] ), .S(\mult_22/SUMB[52][58] ) );
  FA_X1 \mult_22/S2_52_57  ( .A(\mult_22/ab[52][57] ), .B(
        \mult_22/CARRYB[51][57] ), .CI(\mult_22/SUMB[51][58] ), .CO(
        \mult_22/CARRYB[52][57] ), .S(\mult_22/SUMB[52][57] ) );
  FA_X1 \mult_22/S2_52_56  ( .A(\mult_22/ab[52][56] ), .B(
        \mult_22/CARRYB[51][56] ), .CI(\mult_22/SUMB[51][57] ), .CO(
        \mult_22/CARRYB[52][56] ), .S(\mult_22/SUMB[52][56] ) );
  FA_X1 \mult_22/S2_52_55  ( .A(\mult_22/ab[52][55] ), .B(
        \mult_22/CARRYB[51][55] ), .CI(\mult_22/SUMB[51][56] ), .CO(
        \mult_22/CARRYB[52][55] ), .S(\mult_22/SUMB[52][55] ) );
  FA_X1 \mult_22/S2_52_54  ( .A(\mult_22/ab[52][54] ), .B(
        \mult_22/CARRYB[51][54] ), .CI(\mult_22/SUMB[51][55] ), .CO(
        \mult_22/CARRYB[52][54] ), .S(\mult_22/SUMB[52][54] ) );
  FA_X1 \mult_22/S2_52_53  ( .A(\mult_22/ab[52][53] ), .B(
        \mult_22/CARRYB[51][53] ), .CI(\mult_22/SUMB[51][54] ), .CO(
        \mult_22/CARRYB[52][53] ), .S(\mult_22/SUMB[52][53] ) );
  FA_X1 \mult_22/S2_52_52  ( .A(\mult_22/ab[52][52] ), .B(
        \mult_22/CARRYB[51][52] ), .CI(\mult_22/SUMB[51][53] ), .CO(
        \mult_22/CARRYB[52][52] ), .S(\mult_22/SUMB[52][52] ) );
  FA_X1 \mult_22/S2_52_51  ( .A(\mult_22/ab[52][51] ), .B(
        \mult_22/CARRYB[51][51] ), .CI(\mult_22/SUMB[51][52] ), .CO(
        \mult_22/CARRYB[52][51] ), .S(\mult_22/SUMB[52][51] ) );
  FA_X1 \mult_22/S2_52_50  ( .A(\mult_22/ab[52][50] ), .B(
        \mult_22/CARRYB[51][50] ), .CI(\mult_22/SUMB[51][51] ), .CO(
        \mult_22/CARRYB[52][50] ), .S(\mult_22/SUMB[52][50] ) );
  FA_X1 \mult_22/S2_52_49  ( .A(\mult_22/ab[52][49] ), .B(
        \mult_22/CARRYB[51][49] ), .CI(\mult_22/SUMB[51][50] ), .CO(
        \mult_22/CARRYB[52][49] ), .S(\mult_22/SUMB[52][49] ) );
  FA_X1 \mult_22/S2_52_48  ( .A(\mult_22/ab[52][48] ), .B(
        \mult_22/CARRYB[51][48] ), .CI(\mult_22/SUMB[51][49] ), .CO(
        \mult_22/CARRYB[52][48] ), .S(\mult_22/SUMB[52][48] ) );
  FA_X1 \mult_22/S2_52_47  ( .A(\mult_22/ab[52][47] ), .B(
        \mult_22/CARRYB[51][47] ), .CI(\mult_22/SUMB[51][48] ), .CO(
        \mult_22/CARRYB[52][47] ), .S(\mult_22/SUMB[52][47] ) );
  FA_X1 \mult_22/S2_52_46  ( .A(\mult_22/ab[52][46] ), .B(
        \mult_22/CARRYB[51][46] ), .CI(\mult_22/SUMB[51][47] ), .CO(
        \mult_22/CARRYB[52][46] ), .S(\mult_22/SUMB[52][46] ) );
  FA_X1 \mult_22/S2_52_45  ( .A(\mult_22/ab[52][45] ), .B(
        \mult_22/CARRYB[51][45] ), .CI(\mult_22/SUMB[51][46] ), .CO(
        \mult_22/CARRYB[52][45] ), .S(\mult_22/SUMB[52][45] ) );
  FA_X1 \mult_22/S2_52_44  ( .A(\mult_22/ab[52][44] ), .B(
        \mult_22/CARRYB[51][44] ), .CI(\mult_22/SUMB[51][45] ), .CO(
        \mult_22/CARRYB[52][44] ), .S(\mult_22/SUMB[52][44] ) );
  FA_X1 \mult_22/S2_52_43  ( .A(\mult_22/ab[52][43] ), .B(
        \mult_22/CARRYB[51][43] ), .CI(\mult_22/SUMB[51][44] ), .CO(
        \mult_22/CARRYB[52][43] ), .S(\mult_22/SUMB[52][43] ) );
  FA_X1 \mult_22/S2_52_42  ( .A(\mult_22/ab[52][42] ), .B(
        \mult_22/CARRYB[51][42] ), .CI(\mult_22/SUMB[51][43] ), .CO(
        \mult_22/CARRYB[52][42] ), .S(\mult_22/SUMB[52][42] ) );
  FA_X1 \mult_22/S2_52_41  ( .A(\mult_22/ab[52][41] ), .B(
        \mult_22/CARRYB[51][41] ), .CI(\mult_22/SUMB[51][42] ), .CO(
        \mult_22/CARRYB[52][41] ), .S(\mult_22/SUMB[52][41] ) );
  FA_X1 \mult_22/S2_52_40  ( .A(\mult_22/ab[52][40] ), .B(
        \mult_22/CARRYB[51][40] ), .CI(\mult_22/SUMB[51][41] ), .CO(
        \mult_22/CARRYB[52][40] ), .S(\mult_22/SUMB[52][40] ) );
  FA_X1 \mult_22/S2_52_39  ( .A(\mult_22/ab[52][39] ), .B(
        \mult_22/CARRYB[51][39] ), .CI(\mult_22/SUMB[51][40] ), .CO(
        \mult_22/CARRYB[52][39] ), .S(\mult_22/SUMB[52][39] ) );
  FA_X1 \mult_22/S2_52_38  ( .A(\mult_22/ab[52][38] ), .B(
        \mult_22/CARRYB[51][38] ), .CI(\mult_22/SUMB[51][39] ), .CO(
        \mult_22/CARRYB[52][38] ), .S(\mult_22/SUMB[52][38] ) );
  FA_X1 \mult_22/S2_52_37  ( .A(\mult_22/ab[52][37] ), .B(
        \mult_22/CARRYB[51][37] ), .CI(\mult_22/SUMB[51][38] ), .CO(
        \mult_22/CARRYB[52][37] ), .S(\mult_22/SUMB[52][37] ) );
  FA_X1 \mult_22/S2_52_36  ( .A(\mult_22/ab[52][36] ), .B(
        \mult_22/CARRYB[51][36] ), .CI(\mult_22/SUMB[51][37] ), .CO(
        \mult_22/CARRYB[52][36] ), .S(\mult_22/SUMB[52][36] ) );
  FA_X1 \mult_22/S2_52_35  ( .A(\mult_22/ab[52][35] ), .B(
        \mult_22/CARRYB[51][35] ), .CI(\mult_22/SUMB[51][36] ), .CO(
        \mult_22/CARRYB[52][35] ), .S(\mult_22/SUMB[52][35] ) );
  FA_X1 \mult_22/S2_52_34  ( .A(\mult_22/ab[52][34] ), .B(
        \mult_22/CARRYB[51][34] ), .CI(\mult_22/SUMB[51][35] ), .CO(
        \mult_22/CARRYB[52][34] ), .S(\mult_22/SUMB[52][34] ) );
  FA_X1 \mult_22/S2_52_33  ( .A(\mult_22/ab[52][33] ), .B(
        \mult_22/CARRYB[51][33] ), .CI(\mult_22/SUMB[51][34] ), .CO(
        \mult_22/CARRYB[52][33] ), .S(\mult_22/SUMB[52][33] ) );
  FA_X1 \mult_22/S2_52_32  ( .A(\mult_22/ab[52][32] ), .B(
        \mult_22/CARRYB[51][32] ), .CI(\mult_22/SUMB[51][33] ), .CO(
        \mult_22/CARRYB[52][32] ), .S(\mult_22/SUMB[52][32] ) );
  FA_X1 \mult_22/S2_52_31  ( .A(\mult_22/ab[52][31] ), .B(
        \mult_22/CARRYB[51][31] ), .CI(\mult_22/SUMB[51][32] ), .CO(
        \mult_22/CARRYB[52][31] ), .S(\mult_22/SUMB[52][31] ) );
  FA_X1 \mult_22/S2_52_30  ( .A(\mult_22/ab[52][30] ), .B(
        \mult_22/CARRYB[51][30] ), .CI(\mult_22/SUMB[51][31] ), .CO(
        \mult_22/CARRYB[52][30] ), .S(\mult_22/SUMB[52][30] ) );
  FA_X1 \mult_22/S2_52_29  ( .A(\mult_22/ab[52][29] ), .B(
        \mult_22/CARRYB[51][29] ), .CI(\mult_22/SUMB[51][30] ), .CO(
        \mult_22/CARRYB[52][29] ), .S(\mult_22/SUMB[52][29] ) );
  FA_X1 \mult_22/S2_52_28  ( .A(\mult_22/ab[52][28] ), .B(
        \mult_22/CARRYB[51][28] ), .CI(\mult_22/SUMB[51][29] ), .CO(
        \mult_22/CARRYB[52][28] ), .S(\mult_22/SUMB[52][28] ) );
  FA_X1 \mult_22/S2_52_27  ( .A(\mult_22/ab[52][27] ), .B(
        \mult_22/CARRYB[51][27] ), .CI(\mult_22/SUMB[51][28] ), .CO(
        \mult_22/CARRYB[52][27] ), .S(\mult_22/SUMB[52][27] ) );
  FA_X1 \mult_22/S2_52_26  ( .A(\mult_22/ab[52][26] ), .B(
        \mult_22/CARRYB[51][26] ), .CI(\mult_22/SUMB[51][27] ), .CO(
        \mult_22/CARRYB[52][26] ), .S(\mult_22/SUMB[52][26] ) );
  FA_X1 \mult_22/S2_52_25  ( .A(\mult_22/ab[52][25] ), .B(
        \mult_22/CARRYB[51][25] ), .CI(\mult_22/SUMB[51][26] ), .CO(
        \mult_22/CARRYB[52][25] ), .S(\mult_22/SUMB[52][25] ) );
  FA_X1 \mult_22/S2_52_24  ( .A(\mult_22/ab[52][24] ), .B(
        \mult_22/CARRYB[51][24] ), .CI(\mult_22/SUMB[51][25] ), .CO(
        \mult_22/CARRYB[52][24] ), .S(\mult_22/SUMB[52][24] ) );
  FA_X1 \mult_22/S2_52_23  ( .A(\mult_22/ab[52][23] ), .B(
        \mult_22/CARRYB[51][23] ), .CI(\mult_22/SUMB[51][24] ), .CO(
        \mult_22/CARRYB[52][23] ), .S(\mult_22/SUMB[52][23] ) );
  FA_X1 \mult_22/S2_52_22  ( .A(\mult_22/ab[52][22] ), .B(
        \mult_22/CARRYB[51][22] ), .CI(\mult_22/SUMB[51][23] ), .CO(
        \mult_22/CARRYB[52][22] ), .S(\mult_22/SUMB[52][22] ) );
  FA_X1 \mult_22/S2_52_21  ( .A(\mult_22/ab[52][21] ), .B(
        \mult_22/CARRYB[51][21] ), .CI(\mult_22/SUMB[51][22] ), .CO(
        \mult_22/CARRYB[52][21] ), .S(\mult_22/SUMB[52][21] ) );
  FA_X1 \mult_22/S2_52_20  ( .A(\mult_22/ab[52][20] ), .B(
        \mult_22/CARRYB[51][20] ), .CI(\mult_22/SUMB[51][21] ), .CO(
        \mult_22/CARRYB[52][20] ), .S(\mult_22/SUMB[52][20] ) );
  FA_X1 \mult_22/S2_52_19  ( .A(\mult_22/ab[52][19] ), .B(
        \mult_22/CARRYB[51][19] ), .CI(\mult_22/SUMB[51][20] ), .CO(
        \mult_22/CARRYB[52][19] ), .S(\mult_22/SUMB[52][19] ) );
  FA_X1 \mult_22/S2_52_18  ( .A(\mult_22/ab[52][18] ), .B(
        \mult_22/CARRYB[51][18] ), .CI(\mult_22/SUMB[51][19] ), .CO(
        \mult_22/CARRYB[52][18] ), .S(\mult_22/SUMB[52][18] ) );
  FA_X1 \mult_22/S2_52_17  ( .A(\mult_22/ab[52][17] ), .B(
        \mult_22/CARRYB[51][17] ), .CI(\mult_22/SUMB[51][18] ), .CO(
        \mult_22/CARRYB[52][17] ), .S(\mult_22/SUMB[52][17] ) );
  FA_X1 \mult_22/S2_52_16  ( .A(\mult_22/ab[52][16] ), .B(
        \mult_22/CARRYB[51][16] ), .CI(\mult_22/SUMB[51][17] ), .CO(
        \mult_22/CARRYB[52][16] ), .S(\mult_22/SUMB[52][16] ) );
  FA_X1 \mult_22/S2_52_15  ( .A(\mult_22/ab[52][15] ), .B(
        \mult_22/CARRYB[51][15] ), .CI(\mult_22/SUMB[51][16] ), .CO(
        \mult_22/CARRYB[52][15] ), .S(\mult_22/SUMB[52][15] ) );
  FA_X1 \mult_22/S2_52_14  ( .A(\mult_22/ab[52][14] ), .B(
        \mult_22/CARRYB[51][14] ), .CI(\mult_22/SUMB[51][15] ), .CO(
        \mult_22/CARRYB[52][14] ), .S(\mult_22/SUMB[52][14] ) );
  FA_X1 \mult_22/S2_52_13  ( .A(\mult_22/ab[52][13] ), .B(
        \mult_22/CARRYB[51][13] ), .CI(\mult_22/SUMB[51][14] ), .CO(
        \mult_22/CARRYB[52][13] ), .S(\mult_22/SUMB[52][13] ) );
  FA_X1 \mult_22/S2_52_12  ( .A(\mult_22/ab[52][12] ), .B(
        \mult_22/CARRYB[51][12] ), .CI(\mult_22/SUMB[51][13] ), .CO(
        \mult_22/CARRYB[52][12] ), .S(\mult_22/SUMB[52][12] ) );
  FA_X1 \mult_22/S2_52_11  ( .A(\mult_22/ab[52][11] ), .B(
        \mult_22/CARRYB[51][11] ), .CI(\mult_22/SUMB[51][12] ), .CO(
        \mult_22/CARRYB[52][11] ), .S(\mult_22/SUMB[52][11] ) );
  FA_X1 \mult_22/S2_52_10  ( .A(\mult_22/ab[52][10] ), .B(
        \mult_22/CARRYB[51][10] ), .CI(\mult_22/SUMB[51][11] ), .CO(
        \mult_22/CARRYB[52][10] ), .S(\mult_22/SUMB[52][10] ) );
  FA_X1 \mult_22/S2_52_9  ( .A(\mult_22/ab[52][9] ), .B(
        \mult_22/CARRYB[51][9] ), .CI(\mult_22/SUMB[51][10] ), .CO(
        \mult_22/CARRYB[52][9] ), .S(\mult_22/SUMB[52][9] ) );
  FA_X1 \mult_22/S2_52_8  ( .A(\mult_22/ab[52][8] ), .B(
        \mult_22/CARRYB[51][8] ), .CI(\mult_22/SUMB[51][9] ), .CO(
        \mult_22/CARRYB[52][8] ), .S(\mult_22/SUMB[52][8] ) );
  FA_X1 \mult_22/S2_52_7  ( .A(\mult_22/ab[52][7] ), .B(
        \mult_22/CARRYB[51][7] ), .CI(\mult_22/SUMB[51][8] ), .CO(
        \mult_22/CARRYB[52][7] ), .S(\mult_22/SUMB[52][7] ) );
  FA_X1 \mult_22/S2_52_6  ( .A(\mult_22/ab[52][6] ), .B(
        \mult_22/CARRYB[51][6] ), .CI(\mult_22/SUMB[51][7] ), .CO(
        \mult_22/CARRYB[52][6] ), .S(\mult_22/SUMB[52][6] ) );
  FA_X1 \mult_22/S2_52_5  ( .A(\mult_22/ab[52][5] ), .B(
        \mult_22/CARRYB[51][5] ), .CI(\mult_22/SUMB[51][6] ), .CO(
        \mult_22/CARRYB[52][5] ), .S(\mult_22/SUMB[52][5] ) );
  FA_X1 \mult_22/S2_52_4  ( .A(\mult_22/ab[52][4] ), .B(
        \mult_22/CARRYB[51][4] ), .CI(\mult_22/SUMB[51][5] ), .CO(
        \mult_22/CARRYB[52][4] ), .S(\mult_22/SUMB[52][4] ) );
  FA_X1 \mult_22/S2_52_3  ( .A(\mult_22/ab[52][3] ), .B(
        \mult_22/CARRYB[51][3] ), .CI(\mult_22/SUMB[51][4] ), .CO(
        \mult_22/CARRYB[52][3] ), .S(\mult_22/SUMB[52][3] ) );
  FA_X1 \mult_22/S2_52_2  ( .A(\mult_22/ab[52][2] ), .B(
        \mult_22/CARRYB[51][2] ), .CI(\mult_22/SUMB[51][3] ), .CO(
        \mult_22/CARRYB[52][2] ), .S(\mult_22/SUMB[52][2] ) );
  FA_X1 \mult_22/S2_52_1  ( .A(\mult_22/ab[52][1] ), .B(
        \mult_22/CARRYB[51][1] ), .CI(\mult_22/SUMB[51][2] ), .CO(
        \mult_22/CARRYB[52][1] ), .S(\mult_22/SUMB[52][1] ) );
  FA_X1 \mult_22/S1_52_0  ( .A(\mult_22/ab[52][0] ), .B(
        \mult_22/CARRYB[51][0] ), .CI(\mult_22/SUMB[51][1] ), .CO(
        \mult_22/CARRYB[52][0] ), .S(N180) );
  FA_X1 \mult_22/S3_53_62  ( .A(\mult_22/ab[53][62] ), .B(
        \mult_22/CARRYB[52][62] ), .CI(\mult_22/ab[52][63] ), .CO(
        \mult_22/CARRYB[53][62] ), .S(\mult_22/SUMB[53][62] ) );
  FA_X1 \mult_22/S2_53_61  ( .A(\mult_22/ab[53][61] ), .B(
        \mult_22/CARRYB[52][61] ), .CI(\mult_22/SUMB[52][62] ), .CO(
        \mult_22/CARRYB[53][61] ), .S(\mult_22/SUMB[53][61] ) );
  FA_X1 \mult_22/S2_53_60  ( .A(\mult_22/ab[53][60] ), .B(
        \mult_22/CARRYB[52][60] ), .CI(\mult_22/SUMB[52][61] ), .CO(
        \mult_22/CARRYB[53][60] ), .S(\mult_22/SUMB[53][60] ) );
  FA_X1 \mult_22/S2_53_59  ( .A(\mult_22/ab[53][59] ), .B(
        \mult_22/CARRYB[52][59] ), .CI(\mult_22/SUMB[52][60] ), .CO(
        \mult_22/CARRYB[53][59] ), .S(\mult_22/SUMB[53][59] ) );
  FA_X1 \mult_22/S2_53_58  ( .A(\mult_22/ab[53][58] ), .B(
        \mult_22/CARRYB[52][58] ), .CI(\mult_22/SUMB[52][59] ), .CO(
        \mult_22/CARRYB[53][58] ), .S(\mult_22/SUMB[53][58] ) );
  FA_X1 \mult_22/S2_53_57  ( .A(\mult_22/ab[53][57] ), .B(
        \mult_22/CARRYB[52][57] ), .CI(\mult_22/SUMB[52][58] ), .CO(
        \mult_22/CARRYB[53][57] ), .S(\mult_22/SUMB[53][57] ) );
  FA_X1 \mult_22/S2_53_56  ( .A(\mult_22/ab[53][56] ), .B(
        \mult_22/CARRYB[52][56] ), .CI(\mult_22/SUMB[52][57] ), .CO(
        \mult_22/CARRYB[53][56] ), .S(\mult_22/SUMB[53][56] ) );
  FA_X1 \mult_22/S2_53_55  ( .A(\mult_22/ab[53][55] ), .B(
        \mult_22/CARRYB[52][55] ), .CI(\mult_22/SUMB[52][56] ), .CO(
        \mult_22/CARRYB[53][55] ), .S(\mult_22/SUMB[53][55] ) );
  FA_X1 \mult_22/S2_53_54  ( .A(\mult_22/ab[53][54] ), .B(
        \mult_22/CARRYB[52][54] ), .CI(\mult_22/SUMB[52][55] ), .CO(
        \mult_22/CARRYB[53][54] ), .S(\mult_22/SUMB[53][54] ) );
  FA_X1 \mult_22/S2_53_53  ( .A(\mult_22/ab[53][53] ), .B(
        \mult_22/CARRYB[52][53] ), .CI(\mult_22/SUMB[52][54] ), .CO(
        \mult_22/CARRYB[53][53] ), .S(\mult_22/SUMB[53][53] ) );
  FA_X1 \mult_22/S2_53_52  ( .A(\mult_22/ab[53][52] ), .B(
        \mult_22/CARRYB[52][52] ), .CI(\mult_22/SUMB[52][53] ), .CO(
        \mult_22/CARRYB[53][52] ), .S(\mult_22/SUMB[53][52] ) );
  FA_X1 \mult_22/S2_53_51  ( .A(\mult_22/ab[53][51] ), .B(
        \mult_22/CARRYB[52][51] ), .CI(\mult_22/SUMB[52][52] ), .CO(
        \mult_22/CARRYB[53][51] ), .S(\mult_22/SUMB[53][51] ) );
  FA_X1 \mult_22/S2_53_50  ( .A(\mult_22/ab[53][50] ), .B(
        \mult_22/CARRYB[52][50] ), .CI(\mult_22/SUMB[52][51] ), .CO(
        \mult_22/CARRYB[53][50] ), .S(\mult_22/SUMB[53][50] ) );
  FA_X1 \mult_22/S2_53_49  ( .A(\mult_22/ab[53][49] ), .B(
        \mult_22/CARRYB[52][49] ), .CI(\mult_22/SUMB[52][50] ), .CO(
        \mult_22/CARRYB[53][49] ), .S(\mult_22/SUMB[53][49] ) );
  FA_X1 \mult_22/S2_53_48  ( .A(\mult_22/ab[53][48] ), .B(
        \mult_22/CARRYB[52][48] ), .CI(\mult_22/SUMB[52][49] ), .CO(
        \mult_22/CARRYB[53][48] ), .S(\mult_22/SUMB[53][48] ) );
  FA_X1 \mult_22/S2_53_47  ( .A(\mult_22/ab[53][47] ), .B(
        \mult_22/CARRYB[52][47] ), .CI(\mult_22/SUMB[52][48] ), .CO(
        \mult_22/CARRYB[53][47] ), .S(\mult_22/SUMB[53][47] ) );
  FA_X1 \mult_22/S2_53_46  ( .A(\mult_22/ab[53][46] ), .B(
        \mult_22/CARRYB[52][46] ), .CI(\mult_22/SUMB[52][47] ), .CO(
        \mult_22/CARRYB[53][46] ), .S(\mult_22/SUMB[53][46] ) );
  FA_X1 \mult_22/S2_53_45  ( .A(\mult_22/ab[53][45] ), .B(
        \mult_22/CARRYB[52][45] ), .CI(\mult_22/SUMB[52][46] ), .CO(
        \mult_22/CARRYB[53][45] ), .S(\mult_22/SUMB[53][45] ) );
  FA_X1 \mult_22/S2_53_44  ( .A(\mult_22/ab[53][44] ), .B(
        \mult_22/CARRYB[52][44] ), .CI(\mult_22/SUMB[52][45] ), .CO(
        \mult_22/CARRYB[53][44] ), .S(\mult_22/SUMB[53][44] ) );
  FA_X1 \mult_22/S2_53_43  ( .A(\mult_22/ab[53][43] ), .B(
        \mult_22/CARRYB[52][43] ), .CI(\mult_22/SUMB[52][44] ), .CO(
        \mult_22/CARRYB[53][43] ), .S(\mult_22/SUMB[53][43] ) );
  FA_X1 \mult_22/S2_53_42  ( .A(\mult_22/ab[53][42] ), .B(
        \mult_22/CARRYB[52][42] ), .CI(\mult_22/SUMB[52][43] ), .CO(
        \mult_22/CARRYB[53][42] ), .S(\mult_22/SUMB[53][42] ) );
  FA_X1 \mult_22/S2_53_41  ( .A(\mult_22/ab[53][41] ), .B(
        \mult_22/CARRYB[52][41] ), .CI(\mult_22/SUMB[52][42] ), .CO(
        \mult_22/CARRYB[53][41] ), .S(\mult_22/SUMB[53][41] ) );
  FA_X1 \mult_22/S2_53_40  ( .A(\mult_22/ab[53][40] ), .B(
        \mult_22/CARRYB[52][40] ), .CI(\mult_22/SUMB[52][41] ), .CO(
        \mult_22/CARRYB[53][40] ), .S(\mult_22/SUMB[53][40] ) );
  FA_X1 \mult_22/S2_53_39  ( .A(\mult_22/ab[53][39] ), .B(
        \mult_22/CARRYB[52][39] ), .CI(\mult_22/SUMB[52][40] ), .CO(
        \mult_22/CARRYB[53][39] ), .S(\mult_22/SUMB[53][39] ) );
  FA_X1 \mult_22/S2_53_38  ( .A(\mult_22/ab[53][38] ), .B(
        \mult_22/CARRYB[52][38] ), .CI(\mult_22/SUMB[52][39] ), .CO(
        \mult_22/CARRYB[53][38] ), .S(\mult_22/SUMB[53][38] ) );
  FA_X1 \mult_22/S2_53_37  ( .A(\mult_22/ab[53][37] ), .B(
        \mult_22/CARRYB[52][37] ), .CI(\mult_22/SUMB[52][38] ), .CO(
        \mult_22/CARRYB[53][37] ), .S(\mult_22/SUMB[53][37] ) );
  FA_X1 \mult_22/S2_53_36  ( .A(\mult_22/ab[53][36] ), .B(
        \mult_22/CARRYB[52][36] ), .CI(\mult_22/SUMB[52][37] ), .CO(
        \mult_22/CARRYB[53][36] ), .S(\mult_22/SUMB[53][36] ) );
  FA_X1 \mult_22/S2_53_35  ( .A(\mult_22/ab[53][35] ), .B(
        \mult_22/CARRYB[52][35] ), .CI(\mult_22/SUMB[52][36] ), .CO(
        \mult_22/CARRYB[53][35] ), .S(\mult_22/SUMB[53][35] ) );
  FA_X1 \mult_22/S2_53_34  ( .A(\mult_22/ab[53][34] ), .B(
        \mult_22/CARRYB[52][34] ), .CI(\mult_22/SUMB[52][35] ), .CO(
        \mult_22/CARRYB[53][34] ), .S(\mult_22/SUMB[53][34] ) );
  FA_X1 \mult_22/S2_53_33  ( .A(\mult_22/ab[53][33] ), .B(
        \mult_22/CARRYB[52][33] ), .CI(\mult_22/SUMB[52][34] ), .CO(
        \mult_22/CARRYB[53][33] ), .S(\mult_22/SUMB[53][33] ) );
  FA_X1 \mult_22/S2_53_32  ( .A(\mult_22/ab[53][32] ), .B(
        \mult_22/CARRYB[52][32] ), .CI(\mult_22/SUMB[52][33] ), .CO(
        \mult_22/CARRYB[53][32] ), .S(\mult_22/SUMB[53][32] ) );
  FA_X1 \mult_22/S2_53_31  ( .A(\mult_22/ab[53][31] ), .B(
        \mult_22/CARRYB[52][31] ), .CI(\mult_22/SUMB[52][32] ), .CO(
        \mult_22/CARRYB[53][31] ), .S(\mult_22/SUMB[53][31] ) );
  FA_X1 \mult_22/S2_53_30  ( .A(\mult_22/ab[53][30] ), .B(
        \mult_22/CARRYB[52][30] ), .CI(\mult_22/SUMB[52][31] ), .CO(
        \mult_22/CARRYB[53][30] ), .S(\mult_22/SUMB[53][30] ) );
  FA_X1 \mult_22/S2_53_29  ( .A(\mult_22/ab[53][29] ), .B(
        \mult_22/CARRYB[52][29] ), .CI(\mult_22/SUMB[52][30] ), .CO(
        \mult_22/CARRYB[53][29] ), .S(\mult_22/SUMB[53][29] ) );
  FA_X1 \mult_22/S2_53_28  ( .A(\mult_22/ab[53][28] ), .B(
        \mult_22/CARRYB[52][28] ), .CI(\mult_22/SUMB[52][29] ), .CO(
        \mult_22/CARRYB[53][28] ), .S(\mult_22/SUMB[53][28] ) );
  FA_X1 \mult_22/S2_53_27  ( .A(\mult_22/ab[53][27] ), .B(
        \mult_22/CARRYB[52][27] ), .CI(\mult_22/SUMB[52][28] ), .CO(
        \mult_22/CARRYB[53][27] ), .S(\mult_22/SUMB[53][27] ) );
  FA_X1 \mult_22/S2_53_26  ( .A(\mult_22/ab[53][26] ), .B(
        \mult_22/CARRYB[52][26] ), .CI(\mult_22/SUMB[52][27] ), .CO(
        \mult_22/CARRYB[53][26] ), .S(\mult_22/SUMB[53][26] ) );
  FA_X1 \mult_22/S2_53_25  ( .A(\mult_22/ab[53][25] ), .B(
        \mult_22/CARRYB[52][25] ), .CI(\mult_22/SUMB[52][26] ), .CO(
        \mult_22/CARRYB[53][25] ), .S(\mult_22/SUMB[53][25] ) );
  FA_X1 \mult_22/S2_53_24  ( .A(\mult_22/ab[53][24] ), .B(
        \mult_22/CARRYB[52][24] ), .CI(\mult_22/SUMB[52][25] ), .CO(
        \mult_22/CARRYB[53][24] ), .S(\mult_22/SUMB[53][24] ) );
  FA_X1 \mult_22/S2_53_23  ( .A(\mult_22/ab[53][23] ), .B(
        \mult_22/CARRYB[52][23] ), .CI(\mult_22/SUMB[52][24] ), .CO(
        \mult_22/CARRYB[53][23] ), .S(\mult_22/SUMB[53][23] ) );
  FA_X1 \mult_22/S2_53_22  ( .A(\mult_22/ab[53][22] ), .B(
        \mult_22/CARRYB[52][22] ), .CI(\mult_22/SUMB[52][23] ), .CO(
        \mult_22/CARRYB[53][22] ), .S(\mult_22/SUMB[53][22] ) );
  FA_X1 \mult_22/S2_53_21  ( .A(\mult_22/ab[53][21] ), .B(
        \mult_22/CARRYB[52][21] ), .CI(\mult_22/SUMB[52][22] ), .CO(
        \mult_22/CARRYB[53][21] ), .S(\mult_22/SUMB[53][21] ) );
  FA_X1 \mult_22/S2_53_20  ( .A(\mult_22/ab[53][20] ), .B(
        \mult_22/CARRYB[52][20] ), .CI(\mult_22/SUMB[52][21] ), .CO(
        \mult_22/CARRYB[53][20] ), .S(\mult_22/SUMB[53][20] ) );
  FA_X1 \mult_22/S2_53_19  ( .A(\mult_22/ab[53][19] ), .B(
        \mult_22/CARRYB[52][19] ), .CI(\mult_22/SUMB[52][20] ), .CO(
        \mult_22/CARRYB[53][19] ), .S(\mult_22/SUMB[53][19] ) );
  FA_X1 \mult_22/S2_53_18  ( .A(\mult_22/ab[53][18] ), .B(
        \mult_22/CARRYB[52][18] ), .CI(\mult_22/SUMB[52][19] ), .CO(
        \mult_22/CARRYB[53][18] ), .S(\mult_22/SUMB[53][18] ) );
  FA_X1 \mult_22/S2_53_17  ( .A(\mult_22/ab[53][17] ), .B(
        \mult_22/CARRYB[52][17] ), .CI(\mult_22/SUMB[52][18] ), .CO(
        \mult_22/CARRYB[53][17] ), .S(\mult_22/SUMB[53][17] ) );
  FA_X1 \mult_22/S2_53_16  ( .A(\mult_22/ab[53][16] ), .B(
        \mult_22/CARRYB[52][16] ), .CI(\mult_22/SUMB[52][17] ), .CO(
        \mult_22/CARRYB[53][16] ), .S(\mult_22/SUMB[53][16] ) );
  FA_X1 \mult_22/S2_53_15  ( .A(\mult_22/ab[53][15] ), .B(
        \mult_22/CARRYB[52][15] ), .CI(\mult_22/SUMB[52][16] ), .CO(
        \mult_22/CARRYB[53][15] ), .S(\mult_22/SUMB[53][15] ) );
  FA_X1 \mult_22/S2_53_14  ( .A(\mult_22/CARRYB[52][14] ), .B(
        \mult_22/ab[53][14] ), .CI(\mult_22/SUMB[52][15] ), .CO(
        \mult_22/CARRYB[53][14] ), .S(\mult_22/SUMB[53][14] ) );
  FA_X1 \mult_22/S2_53_13  ( .A(\mult_22/CARRYB[52][13] ), .B(
        \mult_22/ab[53][13] ), .CI(\mult_22/SUMB[52][14] ), .CO(
        \mult_22/CARRYB[53][13] ), .S(\mult_22/SUMB[53][13] ) );
  FA_X1 \mult_22/S2_53_12  ( .A(\mult_22/CARRYB[52][12] ), .B(
        \mult_22/ab[53][12] ), .CI(\mult_22/SUMB[52][13] ), .CO(
        \mult_22/CARRYB[53][12] ), .S(\mult_22/SUMB[53][12] ) );
  FA_X1 \mult_22/S2_53_11  ( .A(\mult_22/ab[53][11] ), .B(
        \mult_22/CARRYB[52][11] ), .CI(\mult_22/SUMB[52][12] ), .CO(
        \mult_22/CARRYB[53][11] ), .S(\mult_22/SUMB[53][11] ) );
  FA_X1 \mult_22/S2_53_10  ( .A(\mult_22/ab[53][10] ), .B(
        \mult_22/CARRYB[52][10] ), .CI(\mult_22/SUMB[52][11] ), .CO(
        \mult_22/CARRYB[53][10] ), .S(\mult_22/SUMB[53][10] ) );
  FA_X1 \mult_22/S2_53_9  ( .A(\mult_22/ab[53][9] ), .B(
        \mult_22/CARRYB[52][9] ), .CI(\mult_22/SUMB[52][10] ), .CO(
        \mult_22/CARRYB[53][9] ), .S(\mult_22/SUMB[53][9] ) );
  FA_X1 \mult_22/S2_53_8  ( .A(\mult_22/ab[53][8] ), .B(
        \mult_22/CARRYB[52][8] ), .CI(\mult_22/SUMB[52][9] ), .CO(
        \mult_22/CARRYB[53][8] ), .S(\mult_22/SUMB[53][8] ) );
  FA_X1 \mult_22/S2_53_7  ( .A(\mult_22/ab[53][7] ), .B(
        \mult_22/CARRYB[52][7] ), .CI(\mult_22/SUMB[52][8] ), .CO(
        \mult_22/CARRYB[53][7] ), .S(\mult_22/SUMB[53][7] ) );
  FA_X1 \mult_22/S2_53_6  ( .A(\mult_22/ab[53][6] ), .B(
        \mult_22/CARRYB[52][6] ), .CI(\mult_22/SUMB[52][7] ), .CO(
        \mult_22/CARRYB[53][6] ), .S(\mult_22/SUMB[53][6] ) );
  FA_X1 \mult_22/S2_53_5  ( .A(\mult_22/ab[53][5] ), .B(
        \mult_22/CARRYB[52][5] ), .CI(\mult_22/SUMB[52][6] ), .CO(
        \mult_22/CARRYB[53][5] ), .S(\mult_22/SUMB[53][5] ) );
  FA_X1 \mult_22/S2_53_4  ( .A(\mult_22/ab[53][4] ), .B(
        \mult_22/CARRYB[52][4] ), .CI(\mult_22/SUMB[52][5] ), .CO(
        \mult_22/CARRYB[53][4] ), .S(\mult_22/SUMB[53][4] ) );
  FA_X1 \mult_22/S2_53_3  ( .A(\mult_22/ab[53][3] ), .B(
        \mult_22/CARRYB[52][3] ), .CI(\mult_22/SUMB[52][4] ), .CO(
        \mult_22/CARRYB[53][3] ), .S(\mult_22/SUMB[53][3] ) );
  FA_X1 \mult_22/S2_53_2  ( .A(\mult_22/ab[53][2] ), .B(
        \mult_22/CARRYB[52][2] ), .CI(\mult_22/SUMB[52][3] ), .CO(
        \mult_22/CARRYB[53][2] ), .S(\mult_22/SUMB[53][2] ) );
  FA_X1 \mult_22/S2_53_1  ( .A(\mult_22/ab[53][1] ), .B(
        \mult_22/CARRYB[52][1] ), .CI(\mult_22/SUMB[52][2] ), .CO(
        \mult_22/CARRYB[53][1] ), .S(\mult_22/SUMB[53][1] ) );
  FA_X1 \mult_22/S1_53_0  ( .A(\mult_22/ab[53][0] ), .B(
        \mult_22/CARRYB[52][0] ), .CI(\mult_22/SUMB[52][1] ), .CO(
        \mult_22/CARRYB[53][0] ), .S(N181) );
  FA_X1 \mult_22/S3_54_62  ( .A(\mult_22/ab[54][62] ), .B(
        \mult_22/CARRYB[53][62] ), .CI(\mult_22/ab[53][63] ), .CO(
        \mult_22/CARRYB[54][62] ), .S(\mult_22/SUMB[54][62] ) );
  FA_X1 \mult_22/S2_54_61  ( .A(\mult_22/ab[54][61] ), .B(
        \mult_22/CARRYB[53][61] ), .CI(\mult_22/SUMB[53][62] ), .CO(
        \mult_22/CARRYB[54][61] ), .S(\mult_22/SUMB[54][61] ) );
  FA_X1 \mult_22/S2_54_60  ( .A(\mult_22/ab[54][60] ), .B(
        \mult_22/CARRYB[53][60] ), .CI(\mult_22/SUMB[53][61] ), .CO(
        \mult_22/CARRYB[54][60] ), .S(\mult_22/SUMB[54][60] ) );
  FA_X1 \mult_22/S2_54_59  ( .A(\mult_22/ab[54][59] ), .B(
        \mult_22/CARRYB[53][59] ), .CI(\mult_22/SUMB[53][60] ), .CO(
        \mult_22/CARRYB[54][59] ), .S(\mult_22/SUMB[54][59] ) );
  FA_X1 \mult_22/S2_54_58  ( .A(\mult_22/ab[54][58] ), .B(
        \mult_22/CARRYB[53][58] ), .CI(\mult_22/SUMB[53][59] ), .CO(
        \mult_22/CARRYB[54][58] ), .S(\mult_22/SUMB[54][58] ) );
  FA_X1 \mult_22/S2_54_57  ( .A(\mult_22/ab[54][57] ), .B(
        \mult_22/CARRYB[53][57] ), .CI(\mult_22/SUMB[53][58] ), .CO(
        \mult_22/CARRYB[54][57] ), .S(\mult_22/SUMB[54][57] ) );
  FA_X1 \mult_22/S2_54_56  ( .A(\mult_22/ab[54][56] ), .B(
        \mult_22/CARRYB[53][56] ), .CI(\mult_22/SUMB[53][57] ), .CO(
        \mult_22/CARRYB[54][56] ), .S(\mult_22/SUMB[54][56] ) );
  FA_X1 \mult_22/S2_54_55  ( .A(\mult_22/ab[54][55] ), .B(
        \mult_22/CARRYB[53][55] ), .CI(\mult_22/SUMB[53][56] ), .CO(
        \mult_22/CARRYB[54][55] ), .S(\mult_22/SUMB[54][55] ) );
  FA_X1 \mult_22/S2_54_54  ( .A(\mult_22/ab[54][54] ), .B(
        \mult_22/CARRYB[53][54] ), .CI(\mult_22/SUMB[53][55] ), .CO(
        \mult_22/CARRYB[54][54] ), .S(\mult_22/SUMB[54][54] ) );
  FA_X1 \mult_22/S2_54_53  ( .A(\mult_22/ab[54][53] ), .B(
        \mult_22/CARRYB[53][53] ), .CI(\mult_22/SUMB[53][54] ), .CO(
        \mult_22/CARRYB[54][53] ), .S(\mult_22/SUMB[54][53] ) );
  FA_X1 \mult_22/S2_54_52  ( .A(\mult_22/ab[54][52] ), .B(
        \mult_22/CARRYB[53][52] ), .CI(\mult_22/SUMB[53][53] ), .CO(
        \mult_22/CARRYB[54][52] ), .S(\mult_22/SUMB[54][52] ) );
  FA_X1 \mult_22/S2_54_51  ( .A(\mult_22/ab[54][51] ), .B(
        \mult_22/CARRYB[53][51] ), .CI(\mult_22/SUMB[53][52] ), .CO(
        \mult_22/CARRYB[54][51] ), .S(\mult_22/SUMB[54][51] ) );
  FA_X1 \mult_22/S2_54_50  ( .A(\mult_22/ab[54][50] ), .B(
        \mult_22/CARRYB[53][50] ), .CI(\mult_22/SUMB[53][51] ), .CO(
        \mult_22/CARRYB[54][50] ), .S(\mult_22/SUMB[54][50] ) );
  FA_X1 \mult_22/S2_54_49  ( .A(\mult_22/ab[54][49] ), .B(
        \mult_22/CARRYB[53][49] ), .CI(\mult_22/SUMB[53][50] ), .CO(
        \mult_22/CARRYB[54][49] ), .S(\mult_22/SUMB[54][49] ) );
  FA_X1 \mult_22/S2_54_48  ( .A(\mult_22/ab[54][48] ), .B(
        \mult_22/CARRYB[53][48] ), .CI(\mult_22/SUMB[53][49] ), .CO(
        \mult_22/CARRYB[54][48] ), .S(\mult_22/SUMB[54][48] ) );
  FA_X1 \mult_22/S2_54_47  ( .A(\mult_22/ab[54][47] ), .B(
        \mult_22/CARRYB[53][47] ), .CI(\mult_22/SUMB[53][48] ), .CO(
        \mult_22/CARRYB[54][47] ), .S(\mult_22/SUMB[54][47] ) );
  FA_X1 \mult_22/S2_54_46  ( .A(\mult_22/ab[54][46] ), .B(
        \mult_22/CARRYB[53][46] ), .CI(\mult_22/SUMB[53][47] ), .CO(
        \mult_22/CARRYB[54][46] ), .S(\mult_22/SUMB[54][46] ) );
  FA_X1 \mult_22/S2_54_45  ( .A(\mult_22/ab[54][45] ), .B(
        \mult_22/CARRYB[53][45] ), .CI(\mult_22/SUMB[53][46] ), .CO(
        \mult_22/CARRYB[54][45] ), .S(\mult_22/SUMB[54][45] ) );
  FA_X1 \mult_22/S2_54_44  ( .A(\mult_22/ab[54][44] ), .B(
        \mult_22/CARRYB[53][44] ), .CI(\mult_22/SUMB[53][45] ), .CO(
        \mult_22/CARRYB[54][44] ), .S(\mult_22/SUMB[54][44] ) );
  FA_X1 \mult_22/S2_54_43  ( .A(\mult_22/ab[54][43] ), .B(
        \mult_22/CARRYB[53][43] ), .CI(\mult_22/SUMB[53][44] ), .CO(
        \mult_22/CARRYB[54][43] ), .S(\mult_22/SUMB[54][43] ) );
  FA_X1 \mult_22/S2_54_42  ( .A(\mult_22/ab[54][42] ), .B(
        \mult_22/CARRYB[53][42] ), .CI(\mult_22/SUMB[53][43] ), .CO(
        \mult_22/CARRYB[54][42] ), .S(\mult_22/SUMB[54][42] ) );
  FA_X1 \mult_22/S2_54_41  ( .A(\mult_22/ab[54][41] ), .B(
        \mult_22/CARRYB[53][41] ), .CI(\mult_22/SUMB[53][42] ), .CO(
        \mult_22/CARRYB[54][41] ), .S(\mult_22/SUMB[54][41] ) );
  FA_X1 \mult_22/S2_54_40  ( .A(\mult_22/ab[54][40] ), .B(
        \mult_22/CARRYB[53][40] ), .CI(\mult_22/SUMB[53][41] ), .CO(
        \mult_22/CARRYB[54][40] ), .S(\mult_22/SUMB[54][40] ) );
  FA_X1 \mult_22/S2_54_39  ( .A(\mult_22/ab[54][39] ), .B(
        \mult_22/CARRYB[53][39] ), .CI(\mult_22/SUMB[53][40] ), .CO(
        \mult_22/CARRYB[54][39] ), .S(\mult_22/SUMB[54][39] ) );
  FA_X1 \mult_22/S2_54_38  ( .A(\mult_22/ab[54][38] ), .B(
        \mult_22/CARRYB[53][38] ), .CI(\mult_22/SUMB[53][39] ), .CO(
        \mult_22/CARRYB[54][38] ), .S(\mult_22/SUMB[54][38] ) );
  FA_X1 \mult_22/S2_54_37  ( .A(\mult_22/ab[54][37] ), .B(
        \mult_22/CARRYB[53][37] ), .CI(\mult_22/SUMB[53][38] ), .CO(
        \mult_22/CARRYB[54][37] ), .S(\mult_22/SUMB[54][37] ) );
  FA_X1 \mult_22/S2_54_36  ( .A(\mult_22/ab[54][36] ), .B(
        \mult_22/CARRYB[53][36] ), .CI(\mult_22/SUMB[53][37] ), .CO(
        \mult_22/CARRYB[54][36] ), .S(\mult_22/SUMB[54][36] ) );
  FA_X1 \mult_22/S2_54_35  ( .A(\mult_22/ab[54][35] ), .B(
        \mult_22/CARRYB[53][35] ), .CI(\mult_22/SUMB[53][36] ), .CO(
        \mult_22/CARRYB[54][35] ), .S(\mult_22/SUMB[54][35] ) );
  FA_X1 \mult_22/S2_54_34  ( .A(\mult_22/ab[54][34] ), .B(
        \mult_22/CARRYB[53][34] ), .CI(\mult_22/SUMB[53][35] ), .CO(
        \mult_22/CARRYB[54][34] ), .S(\mult_22/SUMB[54][34] ) );
  FA_X1 \mult_22/S2_54_33  ( .A(\mult_22/ab[54][33] ), .B(
        \mult_22/CARRYB[53][33] ), .CI(\mult_22/SUMB[53][34] ), .CO(
        \mult_22/CARRYB[54][33] ), .S(\mult_22/SUMB[54][33] ) );
  FA_X1 \mult_22/S2_54_32  ( .A(\mult_22/ab[54][32] ), .B(
        \mult_22/CARRYB[53][32] ), .CI(\mult_22/SUMB[53][33] ), .CO(
        \mult_22/CARRYB[54][32] ), .S(\mult_22/SUMB[54][32] ) );
  FA_X1 \mult_22/S2_54_31  ( .A(\mult_22/ab[54][31] ), .B(
        \mult_22/CARRYB[53][31] ), .CI(\mult_22/SUMB[53][32] ), .CO(
        \mult_22/CARRYB[54][31] ), .S(\mult_22/SUMB[54][31] ) );
  FA_X1 \mult_22/S2_54_30  ( .A(\mult_22/ab[54][30] ), .B(
        \mult_22/CARRYB[53][30] ), .CI(\mult_22/SUMB[53][31] ), .CO(
        \mult_22/CARRYB[54][30] ), .S(\mult_22/SUMB[54][30] ) );
  FA_X1 \mult_22/S2_54_29  ( .A(\mult_22/ab[54][29] ), .B(
        \mult_22/CARRYB[53][29] ), .CI(\mult_22/SUMB[53][30] ), .CO(
        \mult_22/CARRYB[54][29] ), .S(\mult_22/SUMB[54][29] ) );
  FA_X1 \mult_22/S2_54_28  ( .A(\mult_22/ab[54][28] ), .B(
        \mult_22/CARRYB[53][28] ), .CI(\mult_22/SUMB[53][29] ), .CO(
        \mult_22/CARRYB[54][28] ), .S(\mult_22/SUMB[54][28] ) );
  FA_X1 \mult_22/S2_54_27  ( .A(\mult_22/ab[54][27] ), .B(
        \mult_22/CARRYB[53][27] ), .CI(\mult_22/SUMB[53][28] ), .CO(
        \mult_22/CARRYB[54][27] ), .S(\mult_22/SUMB[54][27] ) );
  FA_X1 \mult_22/S2_54_26  ( .A(\mult_22/ab[54][26] ), .B(
        \mult_22/CARRYB[53][26] ), .CI(\mult_22/SUMB[53][27] ), .CO(
        \mult_22/CARRYB[54][26] ), .S(\mult_22/SUMB[54][26] ) );
  FA_X1 \mult_22/S2_54_25  ( .A(\mult_22/ab[54][25] ), .B(
        \mult_22/CARRYB[53][25] ), .CI(\mult_22/SUMB[53][26] ), .CO(
        \mult_22/CARRYB[54][25] ), .S(\mult_22/SUMB[54][25] ) );
  FA_X1 \mult_22/S2_54_24  ( .A(\mult_22/ab[54][24] ), .B(
        \mult_22/CARRYB[53][24] ), .CI(\mult_22/SUMB[53][25] ), .CO(
        \mult_22/CARRYB[54][24] ), .S(\mult_22/SUMB[54][24] ) );
  FA_X1 \mult_22/S2_54_23  ( .A(\mult_22/ab[54][23] ), .B(
        \mult_22/CARRYB[53][23] ), .CI(\mult_22/SUMB[53][24] ), .CO(
        \mult_22/CARRYB[54][23] ), .S(\mult_22/SUMB[54][23] ) );
  FA_X1 \mult_22/S2_54_22  ( .A(\mult_22/ab[54][22] ), .B(
        \mult_22/CARRYB[53][22] ), .CI(\mult_22/SUMB[53][23] ), .CO(
        \mult_22/CARRYB[54][22] ), .S(\mult_22/SUMB[54][22] ) );
  FA_X1 \mult_22/S2_54_21  ( .A(\mult_22/ab[54][21] ), .B(
        \mult_22/CARRYB[53][21] ), .CI(\mult_22/SUMB[53][22] ), .CO(
        \mult_22/CARRYB[54][21] ), .S(\mult_22/SUMB[54][21] ) );
  FA_X1 \mult_22/S2_54_20  ( .A(\mult_22/ab[54][20] ), .B(
        \mult_22/CARRYB[53][20] ), .CI(\mult_22/SUMB[53][21] ), .CO(
        \mult_22/CARRYB[54][20] ), .S(\mult_22/SUMB[54][20] ) );
  FA_X1 \mult_22/S2_54_19  ( .A(\mult_22/ab[54][19] ), .B(
        \mult_22/CARRYB[53][19] ), .CI(\mult_22/SUMB[53][20] ), .CO(
        \mult_22/CARRYB[54][19] ), .S(\mult_22/SUMB[54][19] ) );
  FA_X1 \mult_22/S2_54_18  ( .A(\mult_22/ab[54][18] ), .B(
        \mult_22/CARRYB[53][18] ), .CI(\mult_22/SUMB[53][19] ), .CO(
        \mult_22/CARRYB[54][18] ), .S(\mult_22/SUMB[54][18] ) );
  FA_X1 \mult_22/S2_54_17  ( .A(\mult_22/ab[54][17] ), .B(
        \mult_22/CARRYB[53][17] ), .CI(\mult_22/SUMB[53][18] ), .CO(
        \mult_22/CARRYB[54][17] ), .S(\mult_22/SUMB[54][17] ) );
  FA_X1 \mult_22/S2_54_16  ( .A(\mult_22/ab[54][16] ), .B(
        \mult_22/CARRYB[53][16] ), .CI(\mult_22/SUMB[53][17] ), .CO(
        \mult_22/CARRYB[54][16] ), .S(\mult_22/SUMB[54][16] ) );
  FA_X1 \mult_22/S2_54_15  ( .A(\mult_22/ab[54][15] ), .B(
        \mult_22/CARRYB[53][15] ), .CI(\mult_22/SUMB[53][16] ), .CO(
        \mult_22/CARRYB[54][15] ), .S(\mult_22/SUMB[54][15] ) );
  FA_X1 \mult_22/S2_54_14  ( .A(\mult_22/ab[54][14] ), .B(
        \mult_22/CARRYB[53][14] ), .CI(\mult_22/SUMB[53][15] ), .CO(
        \mult_22/CARRYB[54][14] ), .S(\mult_22/SUMB[54][14] ) );
  FA_X1 \mult_22/S2_54_13  ( .A(\mult_22/ab[54][13] ), .B(
        \mult_22/CARRYB[53][13] ), .CI(\mult_22/SUMB[53][14] ), .CO(
        \mult_22/CARRYB[54][13] ), .S(\mult_22/SUMB[54][13] ) );
  FA_X1 \mult_22/S2_54_12  ( .A(\mult_22/CARRYB[53][12] ), .B(
        \mult_22/ab[54][12] ), .CI(\mult_22/SUMB[53][13] ), .CO(
        \mult_22/CARRYB[54][12] ), .S(\mult_22/SUMB[54][12] ) );
  FA_X1 \mult_22/S2_54_11  ( .A(\mult_22/ab[54][11] ), .B(
        \mult_22/CARRYB[53][11] ), .CI(\mult_22/SUMB[53][12] ), .CO(
        \mult_22/CARRYB[54][11] ), .S(\mult_22/SUMB[54][11] ) );
  FA_X1 \mult_22/S2_54_10  ( .A(\mult_22/ab[54][10] ), .B(
        \mult_22/CARRYB[53][10] ), .CI(\mult_22/SUMB[53][11] ), .CO(
        \mult_22/CARRYB[54][10] ), .S(\mult_22/SUMB[54][10] ) );
  FA_X1 \mult_22/S2_54_9  ( .A(\mult_22/ab[54][9] ), .B(
        \mult_22/CARRYB[53][9] ), .CI(\mult_22/SUMB[53][10] ), .CO(
        \mult_22/CARRYB[54][9] ), .S(\mult_22/SUMB[54][9] ) );
  FA_X1 \mult_22/S2_54_8  ( .A(\mult_22/ab[54][8] ), .B(
        \mult_22/CARRYB[53][8] ), .CI(\mult_22/SUMB[53][9] ), .CO(
        \mult_22/CARRYB[54][8] ), .S(\mult_22/SUMB[54][8] ) );
  FA_X1 \mult_22/S2_54_7  ( .A(\mult_22/ab[54][7] ), .B(
        \mult_22/CARRYB[53][7] ), .CI(\mult_22/SUMB[53][8] ), .CO(
        \mult_22/CARRYB[54][7] ), .S(\mult_22/SUMB[54][7] ) );
  FA_X1 \mult_22/S2_54_6  ( .A(\mult_22/ab[54][6] ), .B(
        \mult_22/CARRYB[53][6] ), .CI(\mult_22/SUMB[53][7] ), .CO(
        \mult_22/CARRYB[54][6] ), .S(\mult_22/SUMB[54][6] ) );
  FA_X1 \mult_22/S2_54_5  ( .A(\mult_22/ab[54][5] ), .B(
        \mult_22/CARRYB[53][5] ), .CI(\mult_22/SUMB[53][6] ), .CO(
        \mult_22/CARRYB[54][5] ), .S(\mult_22/SUMB[54][5] ) );
  FA_X1 \mult_22/S2_54_4  ( .A(\mult_22/ab[54][4] ), .B(
        \mult_22/CARRYB[53][4] ), .CI(\mult_22/SUMB[53][5] ), .CO(
        \mult_22/CARRYB[54][4] ), .S(\mult_22/SUMB[54][4] ) );
  FA_X1 \mult_22/S2_54_3  ( .A(\mult_22/ab[54][3] ), .B(
        \mult_22/CARRYB[53][3] ), .CI(\mult_22/SUMB[53][4] ), .CO(
        \mult_22/CARRYB[54][3] ), .S(\mult_22/SUMB[54][3] ) );
  FA_X1 \mult_22/S2_54_2  ( .A(\mult_22/ab[54][2] ), .B(
        \mult_22/CARRYB[53][2] ), .CI(\mult_22/SUMB[53][3] ), .CO(
        \mult_22/CARRYB[54][2] ), .S(\mult_22/SUMB[54][2] ) );
  FA_X1 \mult_22/S2_54_1  ( .A(\mult_22/ab[54][1] ), .B(
        \mult_22/CARRYB[53][1] ), .CI(\mult_22/SUMB[53][2] ), .CO(
        \mult_22/CARRYB[54][1] ), .S(\mult_22/SUMB[54][1] ) );
  FA_X1 \mult_22/S1_54_0  ( .A(\mult_22/ab[54][0] ), .B(
        \mult_22/CARRYB[53][0] ), .CI(\mult_22/SUMB[53][1] ), .CO(
        \mult_22/CARRYB[54][0] ), .S(N182) );
  FA_X1 \mult_22/S3_55_62  ( .A(\mult_22/ab[55][62] ), .B(
        \mult_22/CARRYB[54][62] ), .CI(\mult_22/ab[54][63] ), .CO(
        \mult_22/CARRYB[55][62] ), .S(\mult_22/SUMB[55][62] ) );
  FA_X1 \mult_22/S2_55_61  ( .A(\mult_22/ab[55][61] ), .B(
        \mult_22/CARRYB[54][61] ), .CI(\mult_22/SUMB[54][62] ), .CO(
        \mult_22/CARRYB[55][61] ), .S(\mult_22/SUMB[55][61] ) );
  FA_X1 \mult_22/S2_55_60  ( .A(\mult_22/ab[55][60] ), .B(
        \mult_22/CARRYB[54][60] ), .CI(\mult_22/SUMB[54][61] ), .CO(
        \mult_22/CARRYB[55][60] ), .S(\mult_22/SUMB[55][60] ) );
  FA_X1 \mult_22/S2_55_59  ( .A(\mult_22/ab[55][59] ), .B(
        \mult_22/CARRYB[54][59] ), .CI(\mult_22/SUMB[54][60] ), .CO(
        \mult_22/CARRYB[55][59] ), .S(\mult_22/SUMB[55][59] ) );
  FA_X1 \mult_22/S2_55_58  ( .A(\mult_22/ab[55][58] ), .B(
        \mult_22/CARRYB[54][58] ), .CI(\mult_22/SUMB[54][59] ), .CO(
        \mult_22/CARRYB[55][58] ), .S(\mult_22/SUMB[55][58] ) );
  FA_X1 \mult_22/S2_55_57  ( .A(\mult_22/ab[55][57] ), .B(
        \mult_22/CARRYB[54][57] ), .CI(\mult_22/SUMB[54][58] ), .CO(
        \mult_22/CARRYB[55][57] ), .S(\mult_22/SUMB[55][57] ) );
  FA_X1 \mult_22/S2_55_56  ( .A(\mult_22/ab[55][56] ), .B(
        \mult_22/CARRYB[54][56] ), .CI(\mult_22/SUMB[54][57] ), .CO(
        \mult_22/CARRYB[55][56] ), .S(\mult_22/SUMB[55][56] ) );
  FA_X1 \mult_22/S2_55_55  ( .A(\mult_22/ab[55][55] ), .B(
        \mult_22/CARRYB[54][55] ), .CI(\mult_22/SUMB[54][56] ), .CO(
        \mult_22/CARRYB[55][55] ), .S(\mult_22/SUMB[55][55] ) );
  FA_X1 \mult_22/S2_55_54  ( .A(\mult_22/ab[55][54] ), .B(
        \mult_22/CARRYB[54][54] ), .CI(\mult_22/SUMB[54][55] ), .CO(
        \mult_22/CARRYB[55][54] ), .S(\mult_22/SUMB[55][54] ) );
  FA_X1 \mult_22/S2_55_53  ( .A(\mult_22/ab[55][53] ), .B(
        \mult_22/CARRYB[54][53] ), .CI(\mult_22/SUMB[54][54] ), .CO(
        \mult_22/CARRYB[55][53] ), .S(\mult_22/SUMB[55][53] ) );
  FA_X1 \mult_22/S2_55_52  ( .A(\mult_22/ab[55][52] ), .B(
        \mult_22/CARRYB[54][52] ), .CI(\mult_22/SUMB[54][53] ), .CO(
        \mult_22/CARRYB[55][52] ), .S(\mult_22/SUMB[55][52] ) );
  FA_X1 \mult_22/S2_55_51  ( .A(\mult_22/ab[55][51] ), .B(
        \mult_22/CARRYB[54][51] ), .CI(\mult_22/SUMB[54][52] ), .CO(
        \mult_22/CARRYB[55][51] ), .S(\mult_22/SUMB[55][51] ) );
  FA_X1 \mult_22/S2_55_50  ( .A(\mult_22/ab[55][50] ), .B(
        \mult_22/CARRYB[54][50] ), .CI(\mult_22/SUMB[54][51] ), .CO(
        \mult_22/CARRYB[55][50] ), .S(\mult_22/SUMB[55][50] ) );
  FA_X1 \mult_22/S2_55_49  ( .A(\mult_22/ab[55][49] ), .B(
        \mult_22/CARRYB[54][49] ), .CI(\mult_22/SUMB[54][50] ), .CO(
        \mult_22/CARRYB[55][49] ), .S(\mult_22/SUMB[55][49] ) );
  FA_X1 \mult_22/S2_55_48  ( .A(\mult_22/ab[55][48] ), .B(
        \mult_22/CARRYB[54][48] ), .CI(\mult_22/SUMB[54][49] ), .CO(
        \mult_22/CARRYB[55][48] ), .S(\mult_22/SUMB[55][48] ) );
  FA_X1 \mult_22/S2_55_47  ( .A(\mult_22/ab[55][47] ), .B(
        \mult_22/CARRYB[54][47] ), .CI(\mult_22/SUMB[54][48] ), .CO(
        \mult_22/CARRYB[55][47] ), .S(\mult_22/SUMB[55][47] ) );
  FA_X1 \mult_22/S2_55_46  ( .A(\mult_22/ab[55][46] ), .B(
        \mult_22/CARRYB[54][46] ), .CI(\mult_22/SUMB[54][47] ), .CO(
        \mult_22/CARRYB[55][46] ), .S(\mult_22/SUMB[55][46] ) );
  FA_X1 \mult_22/S2_55_45  ( .A(\mult_22/ab[55][45] ), .B(
        \mult_22/CARRYB[54][45] ), .CI(\mult_22/SUMB[54][46] ), .CO(
        \mult_22/CARRYB[55][45] ), .S(\mult_22/SUMB[55][45] ) );
  FA_X1 \mult_22/S2_55_44  ( .A(\mult_22/ab[55][44] ), .B(
        \mult_22/CARRYB[54][44] ), .CI(\mult_22/SUMB[54][45] ), .CO(
        \mult_22/CARRYB[55][44] ), .S(\mult_22/SUMB[55][44] ) );
  FA_X1 \mult_22/S2_55_43  ( .A(\mult_22/ab[55][43] ), .B(
        \mult_22/CARRYB[54][43] ), .CI(\mult_22/SUMB[54][44] ), .CO(
        \mult_22/CARRYB[55][43] ), .S(\mult_22/SUMB[55][43] ) );
  FA_X1 \mult_22/S2_55_42  ( .A(\mult_22/ab[55][42] ), .B(
        \mult_22/CARRYB[54][42] ), .CI(\mult_22/SUMB[54][43] ), .CO(
        \mult_22/CARRYB[55][42] ), .S(\mult_22/SUMB[55][42] ) );
  FA_X1 \mult_22/S2_55_41  ( .A(\mult_22/ab[55][41] ), .B(
        \mult_22/CARRYB[54][41] ), .CI(\mult_22/SUMB[54][42] ), .CO(
        \mult_22/CARRYB[55][41] ), .S(\mult_22/SUMB[55][41] ) );
  FA_X1 \mult_22/S2_55_40  ( .A(\mult_22/ab[55][40] ), .B(
        \mult_22/CARRYB[54][40] ), .CI(\mult_22/SUMB[54][41] ), .CO(
        \mult_22/CARRYB[55][40] ), .S(\mult_22/SUMB[55][40] ) );
  FA_X1 \mult_22/S2_55_39  ( .A(\mult_22/ab[55][39] ), .B(
        \mult_22/CARRYB[54][39] ), .CI(\mult_22/SUMB[54][40] ), .CO(
        \mult_22/CARRYB[55][39] ), .S(\mult_22/SUMB[55][39] ) );
  FA_X1 \mult_22/S2_55_38  ( .A(\mult_22/ab[55][38] ), .B(
        \mult_22/CARRYB[54][38] ), .CI(\mult_22/SUMB[54][39] ), .CO(
        \mult_22/CARRYB[55][38] ), .S(\mult_22/SUMB[55][38] ) );
  FA_X1 \mult_22/S2_55_37  ( .A(\mult_22/ab[55][37] ), .B(
        \mult_22/CARRYB[54][37] ), .CI(\mult_22/SUMB[54][38] ), .CO(
        \mult_22/CARRYB[55][37] ), .S(\mult_22/SUMB[55][37] ) );
  FA_X1 \mult_22/S2_55_36  ( .A(\mult_22/ab[55][36] ), .B(
        \mult_22/CARRYB[54][36] ), .CI(\mult_22/SUMB[54][37] ), .CO(
        \mult_22/CARRYB[55][36] ), .S(\mult_22/SUMB[55][36] ) );
  FA_X1 \mult_22/S2_55_35  ( .A(\mult_22/ab[55][35] ), .B(
        \mult_22/CARRYB[54][35] ), .CI(\mult_22/SUMB[54][36] ), .CO(
        \mult_22/CARRYB[55][35] ), .S(\mult_22/SUMB[55][35] ) );
  FA_X1 \mult_22/S2_55_34  ( .A(\mult_22/ab[55][34] ), .B(
        \mult_22/CARRYB[54][34] ), .CI(\mult_22/SUMB[54][35] ), .CO(
        \mult_22/CARRYB[55][34] ), .S(\mult_22/SUMB[55][34] ) );
  FA_X1 \mult_22/S2_55_33  ( .A(\mult_22/ab[55][33] ), .B(
        \mult_22/CARRYB[54][33] ), .CI(\mult_22/SUMB[54][34] ), .CO(
        \mult_22/CARRYB[55][33] ), .S(\mult_22/SUMB[55][33] ) );
  FA_X1 \mult_22/S2_55_32  ( .A(\mult_22/ab[55][32] ), .B(
        \mult_22/CARRYB[54][32] ), .CI(\mult_22/SUMB[54][33] ), .CO(
        \mult_22/CARRYB[55][32] ), .S(\mult_22/SUMB[55][32] ) );
  FA_X1 \mult_22/S2_55_31  ( .A(\mult_22/ab[55][31] ), .B(
        \mult_22/CARRYB[54][31] ), .CI(\mult_22/SUMB[54][32] ), .CO(
        \mult_22/CARRYB[55][31] ), .S(\mult_22/SUMB[55][31] ) );
  FA_X1 \mult_22/S2_55_30  ( .A(\mult_22/ab[55][30] ), .B(
        \mult_22/CARRYB[54][30] ), .CI(\mult_22/SUMB[54][31] ), .CO(
        \mult_22/CARRYB[55][30] ), .S(\mult_22/SUMB[55][30] ) );
  FA_X1 \mult_22/S2_55_29  ( .A(\mult_22/ab[55][29] ), .B(
        \mult_22/CARRYB[54][29] ), .CI(\mult_22/SUMB[54][30] ), .CO(
        \mult_22/CARRYB[55][29] ), .S(\mult_22/SUMB[55][29] ) );
  FA_X1 \mult_22/S2_55_28  ( .A(\mult_22/ab[55][28] ), .B(
        \mult_22/CARRYB[54][28] ), .CI(\mult_22/SUMB[54][29] ), .CO(
        \mult_22/CARRYB[55][28] ), .S(\mult_22/SUMB[55][28] ) );
  FA_X1 \mult_22/S2_55_27  ( .A(\mult_22/ab[55][27] ), .B(
        \mult_22/CARRYB[54][27] ), .CI(\mult_22/SUMB[54][28] ), .CO(
        \mult_22/CARRYB[55][27] ), .S(\mult_22/SUMB[55][27] ) );
  FA_X1 \mult_22/S2_55_26  ( .A(\mult_22/ab[55][26] ), .B(
        \mult_22/CARRYB[54][26] ), .CI(\mult_22/SUMB[54][27] ), .CO(
        \mult_22/CARRYB[55][26] ), .S(\mult_22/SUMB[55][26] ) );
  FA_X1 \mult_22/S2_55_25  ( .A(\mult_22/ab[55][25] ), .B(
        \mult_22/CARRYB[54][25] ), .CI(\mult_22/SUMB[54][26] ), .CO(
        \mult_22/CARRYB[55][25] ), .S(\mult_22/SUMB[55][25] ) );
  FA_X1 \mult_22/S2_55_24  ( .A(\mult_22/ab[55][24] ), .B(
        \mult_22/CARRYB[54][24] ), .CI(\mult_22/SUMB[54][25] ), .CO(
        \mult_22/CARRYB[55][24] ), .S(\mult_22/SUMB[55][24] ) );
  FA_X1 \mult_22/S2_55_23  ( .A(\mult_22/ab[55][23] ), .B(
        \mult_22/CARRYB[54][23] ), .CI(\mult_22/SUMB[54][24] ), .CO(
        \mult_22/CARRYB[55][23] ), .S(\mult_22/SUMB[55][23] ) );
  FA_X1 \mult_22/S2_55_22  ( .A(\mult_22/ab[55][22] ), .B(
        \mult_22/CARRYB[54][22] ), .CI(\mult_22/SUMB[54][23] ), .CO(
        \mult_22/CARRYB[55][22] ), .S(\mult_22/SUMB[55][22] ) );
  FA_X1 \mult_22/S2_55_21  ( .A(\mult_22/ab[55][21] ), .B(
        \mult_22/CARRYB[54][21] ), .CI(\mult_22/SUMB[54][22] ), .CO(
        \mult_22/CARRYB[55][21] ), .S(\mult_22/SUMB[55][21] ) );
  FA_X1 \mult_22/S2_55_20  ( .A(\mult_22/ab[55][20] ), .B(
        \mult_22/CARRYB[54][20] ), .CI(\mult_22/SUMB[54][21] ), .CO(
        \mult_22/CARRYB[55][20] ), .S(\mult_22/SUMB[55][20] ) );
  FA_X1 \mult_22/S2_55_19  ( .A(\mult_22/ab[55][19] ), .B(
        \mult_22/CARRYB[54][19] ), .CI(\mult_22/SUMB[54][20] ), .CO(
        \mult_22/CARRYB[55][19] ), .S(\mult_22/SUMB[55][19] ) );
  FA_X1 \mult_22/S2_55_18  ( .A(\mult_22/ab[55][18] ), .B(
        \mult_22/CARRYB[54][18] ), .CI(\mult_22/SUMB[54][19] ), .CO(
        \mult_22/CARRYB[55][18] ), .S(\mult_22/SUMB[55][18] ) );
  FA_X1 \mult_22/S2_55_17  ( .A(\mult_22/ab[55][17] ), .B(
        \mult_22/CARRYB[54][17] ), .CI(\mult_22/SUMB[54][18] ), .CO(
        \mult_22/CARRYB[55][17] ), .S(\mult_22/SUMB[55][17] ) );
  FA_X1 \mult_22/S2_55_16  ( .A(\mult_22/ab[55][16] ), .B(
        \mult_22/CARRYB[54][16] ), .CI(\mult_22/SUMB[54][17] ), .CO(
        \mult_22/CARRYB[55][16] ), .S(\mult_22/SUMB[55][16] ) );
  FA_X1 \mult_22/S2_55_15  ( .A(\mult_22/ab[55][15] ), .B(
        \mult_22/CARRYB[54][15] ), .CI(\mult_22/SUMB[54][16] ), .CO(
        \mult_22/CARRYB[55][15] ), .S(\mult_22/SUMB[55][15] ) );
  FA_X1 \mult_22/S2_55_14  ( .A(\mult_22/ab[55][14] ), .B(
        \mult_22/CARRYB[54][14] ), .CI(\mult_22/SUMB[54][15] ), .CO(
        \mult_22/CARRYB[55][14] ), .S(\mult_22/SUMB[55][14] ) );
  FA_X1 \mult_22/S2_55_13  ( .A(\mult_22/ab[55][13] ), .B(
        \mult_22/CARRYB[54][13] ), .CI(\mult_22/SUMB[54][14] ), .CO(
        \mult_22/CARRYB[55][13] ), .S(\mult_22/SUMB[55][13] ) );
  FA_X1 \mult_22/S2_55_12  ( .A(\mult_22/CARRYB[54][12] ), .B(
        \mult_22/ab[55][12] ), .CI(\mult_22/SUMB[54][13] ), .CO(
        \mult_22/CARRYB[55][12] ), .S(\mult_22/SUMB[55][12] ) );
  FA_X1 \mult_22/S2_55_11  ( .A(\mult_22/CARRYB[54][11] ), .B(
        \mult_22/ab[55][11] ), .CI(\mult_22/SUMB[54][12] ), .CO(
        \mult_22/CARRYB[55][11] ), .S(\mult_22/SUMB[55][11] ) );
  FA_X1 \mult_22/S2_55_10  ( .A(\mult_22/ab[55][10] ), .B(
        \mult_22/CARRYB[54][10] ), .CI(\mult_22/SUMB[54][11] ), .CO(
        \mult_22/CARRYB[55][10] ), .S(\mult_22/SUMB[55][10] ) );
  FA_X1 \mult_22/S2_55_9  ( .A(\mult_22/ab[55][9] ), .B(
        \mult_22/CARRYB[54][9] ), .CI(\mult_22/SUMB[54][10] ), .CO(
        \mult_22/CARRYB[55][9] ), .S(\mult_22/SUMB[55][9] ) );
  FA_X1 \mult_22/S2_55_8  ( .A(\mult_22/ab[55][8] ), .B(
        \mult_22/CARRYB[54][8] ), .CI(\mult_22/SUMB[54][9] ), .CO(
        \mult_22/CARRYB[55][8] ), .S(\mult_22/SUMB[55][8] ) );
  FA_X1 \mult_22/S2_55_7  ( .A(\mult_22/ab[55][7] ), .B(
        \mult_22/CARRYB[54][7] ), .CI(\mult_22/SUMB[54][8] ), .CO(
        \mult_22/CARRYB[55][7] ), .S(\mult_22/SUMB[55][7] ) );
  FA_X1 \mult_22/S2_55_6  ( .A(\mult_22/ab[55][6] ), .B(
        \mult_22/CARRYB[54][6] ), .CI(\mult_22/SUMB[54][7] ), .CO(
        \mult_22/CARRYB[55][6] ), .S(\mult_22/SUMB[55][6] ) );
  FA_X1 \mult_22/S2_55_5  ( .A(\mult_22/ab[55][5] ), .B(
        \mult_22/CARRYB[54][5] ), .CI(\mult_22/SUMB[54][6] ), .CO(
        \mult_22/CARRYB[55][5] ), .S(\mult_22/SUMB[55][5] ) );
  FA_X1 \mult_22/S2_55_4  ( .A(\mult_22/ab[55][4] ), .B(
        \mult_22/CARRYB[54][4] ), .CI(\mult_22/SUMB[54][5] ), .CO(
        \mult_22/CARRYB[55][4] ), .S(\mult_22/SUMB[55][4] ) );
  FA_X1 \mult_22/S2_55_3  ( .A(\mult_22/ab[55][3] ), .B(
        \mult_22/CARRYB[54][3] ), .CI(\mult_22/SUMB[54][4] ), .CO(
        \mult_22/CARRYB[55][3] ), .S(\mult_22/SUMB[55][3] ) );
  FA_X1 \mult_22/S2_55_2  ( .A(\mult_22/ab[55][2] ), .B(
        \mult_22/CARRYB[54][2] ), .CI(\mult_22/SUMB[54][3] ), .CO(
        \mult_22/CARRYB[55][2] ), .S(\mult_22/SUMB[55][2] ) );
  FA_X1 \mult_22/S2_55_1  ( .A(\mult_22/ab[55][1] ), .B(
        \mult_22/CARRYB[54][1] ), .CI(\mult_22/SUMB[54][2] ), .CO(
        \mult_22/CARRYB[55][1] ), .S(\mult_22/SUMB[55][1] ) );
  FA_X1 \mult_22/S1_55_0  ( .A(\mult_22/ab[55][0] ), .B(
        \mult_22/CARRYB[54][0] ), .CI(\mult_22/SUMB[54][1] ), .CO(
        \mult_22/CARRYB[55][0] ), .S(N183) );
  FA_X1 \mult_22/S3_56_62  ( .A(\mult_22/ab[56][62] ), .B(
        \mult_22/CARRYB[55][62] ), .CI(\mult_22/ab[55][63] ), .CO(
        \mult_22/CARRYB[56][62] ), .S(\mult_22/SUMB[56][62] ) );
  FA_X1 \mult_22/S2_56_61  ( .A(\mult_22/ab[56][61] ), .B(
        \mult_22/CARRYB[55][61] ), .CI(\mult_22/SUMB[55][62] ), .CO(
        \mult_22/CARRYB[56][61] ), .S(\mult_22/SUMB[56][61] ) );
  FA_X1 \mult_22/S2_56_60  ( .A(\mult_22/ab[56][60] ), .B(
        \mult_22/CARRYB[55][60] ), .CI(\mult_22/SUMB[55][61] ), .CO(
        \mult_22/CARRYB[56][60] ), .S(\mult_22/SUMB[56][60] ) );
  FA_X1 \mult_22/S2_56_59  ( .A(\mult_22/ab[56][59] ), .B(
        \mult_22/CARRYB[55][59] ), .CI(\mult_22/SUMB[55][60] ), .CO(
        \mult_22/CARRYB[56][59] ), .S(\mult_22/SUMB[56][59] ) );
  FA_X1 \mult_22/S2_56_58  ( .A(\mult_22/ab[56][58] ), .B(
        \mult_22/CARRYB[55][58] ), .CI(\mult_22/SUMB[55][59] ), .CO(
        \mult_22/CARRYB[56][58] ), .S(\mult_22/SUMB[56][58] ) );
  FA_X1 \mult_22/S2_56_57  ( .A(\mult_22/ab[56][57] ), .B(
        \mult_22/CARRYB[55][57] ), .CI(\mult_22/SUMB[55][58] ), .CO(
        \mult_22/CARRYB[56][57] ), .S(\mult_22/SUMB[56][57] ) );
  FA_X1 \mult_22/S2_56_56  ( .A(\mult_22/ab[56][56] ), .B(
        \mult_22/CARRYB[55][56] ), .CI(\mult_22/SUMB[55][57] ), .CO(
        \mult_22/CARRYB[56][56] ), .S(\mult_22/SUMB[56][56] ) );
  FA_X1 \mult_22/S2_56_55  ( .A(\mult_22/ab[56][55] ), .B(
        \mult_22/CARRYB[55][55] ), .CI(\mult_22/SUMB[55][56] ), .CO(
        \mult_22/CARRYB[56][55] ), .S(\mult_22/SUMB[56][55] ) );
  FA_X1 \mult_22/S2_56_54  ( .A(\mult_22/ab[56][54] ), .B(
        \mult_22/CARRYB[55][54] ), .CI(\mult_22/SUMB[55][55] ), .CO(
        \mult_22/CARRYB[56][54] ), .S(\mult_22/SUMB[56][54] ) );
  FA_X1 \mult_22/S2_56_53  ( .A(\mult_22/ab[56][53] ), .B(
        \mult_22/CARRYB[55][53] ), .CI(\mult_22/SUMB[55][54] ), .CO(
        \mult_22/CARRYB[56][53] ), .S(\mult_22/SUMB[56][53] ) );
  FA_X1 \mult_22/S2_56_52  ( .A(\mult_22/ab[56][52] ), .B(
        \mult_22/CARRYB[55][52] ), .CI(\mult_22/SUMB[55][53] ), .CO(
        \mult_22/CARRYB[56][52] ), .S(\mult_22/SUMB[56][52] ) );
  FA_X1 \mult_22/S2_56_51  ( .A(\mult_22/ab[56][51] ), .B(
        \mult_22/CARRYB[55][51] ), .CI(\mult_22/SUMB[55][52] ), .CO(
        \mult_22/CARRYB[56][51] ), .S(\mult_22/SUMB[56][51] ) );
  FA_X1 \mult_22/S2_56_50  ( .A(\mult_22/ab[56][50] ), .B(
        \mult_22/CARRYB[55][50] ), .CI(\mult_22/SUMB[55][51] ), .CO(
        \mult_22/CARRYB[56][50] ), .S(\mult_22/SUMB[56][50] ) );
  FA_X1 \mult_22/S2_56_49  ( .A(\mult_22/ab[56][49] ), .B(
        \mult_22/CARRYB[55][49] ), .CI(\mult_22/SUMB[55][50] ), .CO(
        \mult_22/CARRYB[56][49] ), .S(\mult_22/SUMB[56][49] ) );
  FA_X1 \mult_22/S2_56_48  ( .A(\mult_22/ab[56][48] ), .B(
        \mult_22/CARRYB[55][48] ), .CI(\mult_22/SUMB[55][49] ), .CO(
        \mult_22/CARRYB[56][48] ), .S(\mult_22/SUMB[56][48] ) );
  FA_X1 \mult_22/S2_56_47  ( .A(\mult_22/ab[56][47] ), .B(
        \mult_22/CARRYB[55][47] ), .CI(\mult_22/SUMB[55][48] ), .CO(
        \mult_22/CARRYB[56][47] ), .S(\mult_22/SUMB[56][47] ) );
  FA_X1 \mult_22/S2_56_46  ( .A(\mult_22/ab[56][46] ), .B(
        \mult_22/CARRYB[55][46] ), .CI(\mult_22/SUMB[55][47] ), .CO(
        \mult_22/CARRYB[56][46] ), .S(\mult_22/SUMB[56][46] ) );
  FA_X1 \mult_22/S2_56_45  ( .A(\mult_22/ab[56][45] ), .B(
        \mult_22/CARRYB[55][45] ), .CI(\mult_22/SUMB[55][46] ), .CO(
        \mult_22/CARRYB[56][45] ), .S(\mult_22/SUMB[56][45] ) );
  FA_X1 \mult_22/S2_56_44  ( .A(\mult_22/ab[56][44] ), .B(
        \mult_22/CARRYB[55][44] ), .CI(\mult_22/SUMB[55][45] ), .CO(
        \mult_22/CARRYB[56][44] ), .S(\mult_22/SUMB[56][44] ) );
  FA_X1 \mult_22/S2_56_43  ( .A(\mult_22/ab[56][43] ), .B(
        \mult_22/CARRYB[55][43] ), .CI(\mult_22/SUMB[55][44] ), .CO(
        \mult_22/CARRYB[56][43] ), .S(\mult_22/SUMB[56][43] ) );
  FA_X1 \mult_22/S2_56_42  ( .A(\mult_22/ab[56][42] ), .B(
        \mult_22/CARRYB[55][42] ), .CI(\mult_22/SUMB[55][43] ), .CO(
        \mult_22/CARRYB[56][42] ), .S(\mult_22/SUMB[56][42] ) );
  FA_X1 \mult_22/S2_56_41  ( .A(\mult_22/ab[56][41] ), .B(
        \mult_22/CARRYB[55][41] ), .CI(\mult_22/SUMB[55][42] ), .CO(
        \mult_22/CARRYB[56][41] ), .S(\mult_22/SUMB[56][41] ) );
  FA_X1 \mult_22/S2_56_40  ( .A(\mult_22/ab[56][40] ), .B(
        \mult_22/CARRYB[55][40] ), .CI(\mult_22/SUMB[55][41] ), .CO(
        \mult_22/CARRYB[56][40] ), .S(\mult_22/SUMB[56][40] ) );
  FA_X1 \mult_22/S2_56_39  ( .A(\mult_22/ab[56][39] ), .B(
        \mult_22/CARRYB[55][39] ), .CI(\mult_22/SUMB[55][40] ), .CO(
        \mult_22/CARRYB[56][39] ), .S(\mult_22/SUMB[56][39] ) );
  FA_X1 \mult_22/S2_56_38  ( .A(\mult_22/ab[56][38] ), .B(
        \mult_22/CARRYB[55][38] ), .CI(\mult_22/SUMB[55][39] ), .CO(
        \mult_22/CARRYB[56][38] ), .S(\mult_22/SUMB[56][38] ) );
  FA_X1 \mult_22/S2_56_37  ( .A(\mult_22/ab[56][37] ), .B(
        \mult_22/CARRYB[55][37] ), .CI(\mult_22/SUMB[55][38] ), .CO(
        \mult_22/CARRYB[56][37] ), .S(\mult_22/SUMB[56][37] ) );
  FA_X1 \mult_22/S2_56_36  ( .A(\mult_22/ab[56][36] ), .B(
        \mult_22/CARRYB[55][36] ), .CI(\mult_22/SUMB[55][37] ), .CO(
        \mult_22/CARRYB[56][36] ), .S(\mult_22/SUMB[56][36] ) );
  FA_X1 \mult_22/S2_56_35  ( .A(\mult_22/ab[56][35] ), .B(
        \mult_22/CARRYB[55][35] ), .CI(\mult_22/SUMB[55][36] ), .CO(
        \mult_22/CARRYB[56][35] ), .S(\mult_22/SUMB[56][35] ) );
  FA_X1 \mult_22/S2_56_34  ( .A(\mult_22/ab[56][34] ), .B(
        \mult_22/CARRYB[55][34] ), .CI(\mult_22/SUMB[55][35] ), .CO(
        \mult_22/CARRYB[56][34] ), .S(\mult_22/SUMB[56][34] ) );
  FA_X1 \mult_22/S2_56_33  ( .A(\mult_22/ab[56][33] ), .B(
        \mult_22/CARRYB[55][33] ), .CI(\mult_22/SUMB[55][34] ), .CO(
        \mult_22/CARRYB[56][33] ), .S(\mult_22/SUMB[56][33] ) );
  FA_X1 \mult_22/S2_56_32  ( .A(\mult_22/ab[56][32] ), .B(
        \mult_22/CARRYB[55][32] ), .CI(\mult_22/SUMB[55][33] ), .CO(
        \mult_22/CARRYB[56][32] ), .S(\mult_22/SUMB[56][32] ) );
  FA_X1 \mult_22/S2_56_31  ( .A(\mult_22/ab[56][31] ), .B(
        \mult_22/CARRYB[55][31] ), .CI(\mult_22/SUMB[55][32] ), .CO(
        \mult_22/CARRYB[56][31] ), .S(\mult_22/SUMB[56][31] ) );
  FA_X1 \mult_22/S2_56_30  ( .A(\mult_22/ab[56][30] ), .B(
        \mult_22/CARRYB[55][30] ), .CI(\mult_22/SUMB[55][31] ), .CO(
        \mult_22/CARRYB[56][30] ), .S(\mult_22/SUMB[56][30] ) );
  FA_X1 \mult_22/S2_56_29  ( .A(\mult_22/ab[56][29] ), .B(
        \mult_22/CARRYB[55][29] ), .CI(\mult_22/SUMB[55][30] ), .CO(
        \mult_22/CARRYB[56][29] ), .S(\mult_22/SUMB[56][29] ) );
  FA_X1 \mult_22/S2_56_28  ( .A(\mult_22/ab[56][28] ), .B(
        \mult_22/CARRYB[55][28] ), .CI(\mult_22/SUMB[55][29] ), .CO(
        \mult_22/CARRYB[56][28] ), .S(\mult_22/SUMB[56][28] ) );
  FA_X1 \mult_22/S2_56_27  ( .A(\mult_22/ab[56][27] ), .B(
        \mult_22/CARRYB[55][27] ), .CI(\mult_22/SUMB[55][28] ), .CO(
        \mult_22/CARRYB[56][27] ), .S(\mult_22/SUMB[56][27] ) );
  FA_X1 \mult_22/S2_56_26  ( .A(\mult_22/ab[56][26] ), .B(
        \mult_22/CARRYB[55][26] ), .CI(\mult_22/SUMB[55][27] ), .CO(
        \mult_22/CARRYB[56][26] ), .S(\mult_22/SUMB[56][26] ) );
  FA_X1 \mult_22/S2_56_25  ( .A(\mult_22/ab[56][25] ), .B(
        \mult_22/CARRYB[55][25] ), .CI(\mult_22/SUMB[55][26] ), .CO(
        \mult_22/CARRYB[56][25] ), .S(\mult_22/SUMB[56][25] ) );
  FA_X1 \mult_22/S2_56_24  ( .A(\mult_22/ab[56][24] ), .B(
        \mult_22/CARRYB[55][24] ), .CI(\mult_22/SUMB[55][25] ), .CO(
        \mult_22/CARRYB[56][24] ), .S(\mult_22/SUMB[56][24] ) );
  FA_X1 \mult_22/S2_56_23  ( .A(\mult_22/ab[56][23] ), .B(
        \mult_22/CARRYB[55][23] ), .CI(\mult_22/SUMB[55][24] ), .CO(
        \mult_22/CARRYB[56][23] ), .S(\mult_22/SUMB[56][23] ) );
  FA_X1 \mult_22/S2_56_22  ( .A(\mult_22/ab[56][22] ), .B(
        \mult_22/CARRYB[55][22] ), .CI(\mult_22/SUMB[55][23] ), .CO(
        \mult_22/CARRYB[56][22] ), .S(\mult_22/SUMB[56][22] ) );
  FA_X1 \mult_22/S2_56_21  ( .A(\mult_22/ab[56][21] ), .B(
        \mult_22/CARRYB[55][21] ), .CI(\mult_22/SUMB[55][22] ), .CO(
        \mult_22/CARRYB[56][21] ), .S(\mult_22/SUMB[56][21] ) );
  FA_X1 \mult_22/S2_56_20  ( .A(\mult_22/ab[56][20] ), .B(
        \mult_22/CARRYB[55][20] ), .CI(\mult_22/SUMB[55][21] ), .CO(
        \mult_22/CARRYB[56][20] ), .S(\mult_22/SUMB[56][20] ) );
  FA_X1 \mult_22/S2_56_19  ( .A(\mult_22/ab[56][19] ), .B(
        \mult_22/CARRYB[55][19] ), .CI(\mult_22/SUMB[55][20] ), .CO(
        \mult_22/CARRYB[56][19] ), .S(\mult_22/SUMB[56][19] ) );
  FA_X1 \mult_22/S2_56_18  ( .A(\mult_22/ab[56][18] ), .B(
        \mult_22/CARRYB[55][18] ), .CI(\mult_22/SUMB[55][19] ), .CO(
        \mult_22/CARRYB[56][18] ), .S(\mult_22/SUMB[56][18] ) );
  FA_X1 \mult_22/S2_56_17  ( .A(\mult_22/ab[56][17] ), .B(
        \mult_22/CARRYB[55][17] ), .CI(\mult_22/SUMB[55][18] ), .CO(
        \mult_22/CARRYB[56][17] ), .S(\mult_22/SUMB[56][17] ) );
  FA_X1 \mult_22/S2_56_16  ( .A(\mult_22/ab[56][16] ), .B(
        \mult_22/CARRYB[55][16] ), .CI(\mult_22/SUMB[55][17] ), .CO(
        \mult_22/CARRYB[56][16] ), .S(\mult_22/SUMB[56][16] ) );
  FA_X1 \mult_22/S2_56_15  ( .A(\mult_22/ab[56][15] ), .B(
        \mult_22/CARRYB[55][15] ), .CI(\mult_22/SUMB[55][16] ), .CO(
        \mult_22/CARRYB[56][15] ), .S(\mult_22/SUMB[56][15] ) );
  FA_X1 \mult_22/S2_56_14  ( .A(\mult_22/ab[56][14] ), .B(
        \mult_22/CARRYB[55][14] ), .CI(\mult_22/SUMB[55][15] ), .CO(
        \mult_22/CARRYB[56][14] ), .S(\mult_22/SUMB[56][14] ) );
  FA_X1 \mult_22/S2_56_13  ( .A(\mult_22/ab[56][13] ), .B(
        \mult_22/CARRYB[55][13] ), .CI(\mult_22/SUMB[55][14] ), .CO(
        \mult_22/CARRYB[56][13] ), .S(\mult_22/SUMB[56][13] ) );
  FA_X1 \mult_22/S2_56_12  ( .A(\mult_22/ab[56][12] ), .B(
        \mult_22/CARRYB[55][12] ), .CI(\mult_22/SUMB[55][13] ), .CO(
        \mult_22/CARRYB[56][12] ), .S(\mult_22/SUMB[56][12] ) );
  FA_X1 \mult_22/S2_56_11  ( .A(\mult_22/ab[56][11] ), .B(
        \mult_22/CARRYB[55][11] ), .CI(\mult_22/SUMB[55][12] ), .CO(
        \mult_22/CARRYB[56][11] ), .S(\mult_22/SUMB[56][11] ) );
  FA_X1 \mult_22/S2_56_10  ( .A(\mult_22/CARRYB[55][10] ), .B(
        \mult_22/ab[56][10] ), .CI(\mult_22/SUMB[55][11] ), .CO(
        \mult_22/CARRYB[56][10] ), .S(\mult_22/SUMB[56][10] ) );
  FA_X1 \mult_22/S2_56_9  ( .A(\mult_22/CARRYB[55][9] ), .B(
        \mult_22/ab[56][9] ), .CI(\mult_22/SUMB[55][10] ), .CO(
        \mult_22/CARRYB[56][9] ), .S(\mult_22/SUMB[56][9] ) );
  FA_X1 \mult_22/S2_56_8  ( .A(\mult_22/ab[56][8] ), .B(
        \mult_22/CARRYB[55][8] ), .CI(\mult_22/SUMB[55][9] ), .CO(
        \mult_22/CARRYB[56][8] ), .S(\mult_22/SUMB[56][8] ) );
  FA_X1 \mult_22/S2_56_7  ( .A(\mult_22/ab[56][7] ), .B(
        \mult_22/CARRYB[55][7] ), .CI(\mult_22/SUMB[55][8] ), .CO(
        \mult_22/CARRYB[56][7] ), .S(\mult_22/SUMB[56][7] ) );
  FA_X1 \mult_22/S2_56_6  ( .A(\mult_22/ab[56][6] ), .B(
        \mult_22/CARRYB[55][6] ), .CI(\mult_22/SUMB[55][7] ), .CO(
        \mult_22/CARRYB[56][6] ), .S(\mult_22/SUMB[56][6] ) );
  FA_X1 \mult_22/S2_56_5  ( .A(\mult_22/ab[56][5] ), .B(
        \mult_22/CARRYB[55][5] ), .CI(\mult_22/SUMB[55][6] ), .CO(
        \mult_22/CARRYB[56][5] ), .S(\mult_22/SUMB[56][5] ) );
  FA_X1 \mult_22/S2_56_4  ( .A(\mult_22/ab[56][4] ), .B(
        \mult_22/CARRYB[55][4] ), .CI(\mult_22/SUMB[55][5] ), .CO(
        \mult_22/CARRYB[56][4] ), .S(\mult_22/SUMB[56][4] ) );
  FA_X1 \mult_22/S2_56_3  ( .A(\mult_22/ab[56][3] ), .B(
        \mult_22/CARRYB[55][3] ), .CI(\mult_22/SUMB[55][4] ), .CO(
        \mult_22/CARRYB[56][3] ), .S(\mult_22/SUMB[56][3] ) );
  FA_X1 \mult_22/S2_56_2  ( .A(\mult_22/ab[56][2] ), .B(
        \mult_22/CARRYB[55][2] ), .CI(\mult_22/SUMB[55][3] ), .CO(
        \mult_22/CARRYB[56][2] ), .S(\mult_22/SUMB[56][2] ) );
  FA_X1 \mult_22/S2_56_1  ( .A(\mult_22/ab[56][1] ), .B(
        \mult_22/CARRYB[55][1] ), .CI(\mult_22/SUMB[55][2] ), .CO(
        \mult_22/CARRYB[56][1] ), .S(\mult_22/SUMB[56][1] ) );
  FA_X1 \mult_22/S1_56_0  ( .A(\mult_22/ab[56][0] ), .B(
        \mult_22/CARRYB[55][0] ), .CI(\mult_22/SUMB[55][1] ), .CO(
        \mult_22/CARRYB[56][0] ), .S(N184) );
  FA_X1 \mult_22/S3_57_62  ( .A(\mult_22/ab[57][62] ), .B(
        \mult_22/CARRYB[56][62] ), .CI(\mult_22/ab[56][63] ), .CO(
        \mult_22/CARRYB[57][62] ), .S(\mult_22/SUMB[57][62] ) );
  FA_X1 \mult_22/S2_57_61  ( .A(\mult_22/ab[57][61] ), .B(
        \mult_22/CARRYB[56][61] ), .CI(\mult_22/SUMB[56][62] ), .CO(
        \mult_22/CARRYB[57][61] ), .S(\mult_22/SUMB[57][61] ) );
  FA_X1 \mult_22/S2_57_60  ( .A(\mult_22/ab[57][60] ), .B(
        \mult_22/CARRYB[56][60] ), .CI(\mult_22/SUMB[56][61] ), .CO(
        \mult_22/CARRYB[57][60] ), .S(\mult_22/SUMB[57][60] ) );
  FA_X1 \mult_22/S2_57_59  ( .A(\mult_22/ab[57][59] ), .B(
        \mult_22/CARRYB[56][59] ), .CI(\mult_22/SUMB[56][60] ), .CO(
        \mult_22/CARRYB[57][59] ), .S(\mult_22/SUMB[57][59] ) );
  FA_X1 \mult_22/S2_57_58  ( .A(\mult_22/ab[57][58] ), .B(
        \mult_22/CARRYB[56][58] ), .CI(\mult_22/SUMB[56][59] ), .CO(
        \mult_22/CARRYB[57][58] ), .S(\mult_22/SUMB[57][58] ) );
  FA_X1 \mult_22/S2_57_57  ( .A(\mult_22/ab[57][57] ), .B(
        \mult_22/CARRYB[56][57] ), .CI(\mult_22/SUMB[56][58] ), .CO(
        \mult_22/CARRYB[57][57] ), .S(\mult_22/SUMB[57][57] ) );
  FA_X1 \mult_22/S2_57_56  ( .A(\mult_22/ab[57][56] ), .B(
        \mult_22/CARRYB[56][56] ), .CI(\mult_22/SUMB[56][57] ), .CO(
        \mult_22/CARRYB[57][56] ), .S(\mult_22/SUMB[57][56] ) );
  FA_X1 \mult_22/S2_57_55  ( .A(\mult_22/ab[57][55] ), .B(
        \mult_22/CARRYB[56][55] ), .CI(\mult_22/SUMB[56][56] ), .CO(
        \mult_22/CARRYB[57][55] ), .S(\mult_22/SUMB[57][55] ) );
  FA_X1 \mult_22/S2_57_54  ( .A(\mult_22/ab[57][54] ), .B(
        \mult_22/CARRYB[56][54] ), .CI(\mult_22/SUMB[56][55] ), .CO(
        \mult_22/CARRYB[57][54] ), .S(\mult_22/SUMB[57][54] ) );
  FA_X1 \mult_22/S2_57_53  ( .A(\mult_22/ab[57][53] ), .B(
        \mult_22/CARRYB[56][53] ), .CI(\mult_22/SUMB[56][54] ), .CO(
        \mult_22/CARRYB[57][53] ), .S(\mult_22/SUMB[57][53] ) );
  FA_X1 \mult_22/S2_57_52  ( .A(\mult_22/ab[57][52] ), .B(
        \mult_22/CARRYB[56][52] ), .CI(\mult_22/SUMB[56][53] ), .CO(
        \mult_22/CARRYB[57][52] ), .S(\mult_22/SUMB[57][52] ) );
  FA_X1 \mult_22/S2_57_51  ( .A(\mult_22/ab[57][51] ), .B(
        \mult_22/CARRYB[56][51] ), .CI(\mult_22/SUMB[56][52] ), .CO(
        \mult_22/CARRYB[57][51] ), .S(\mult_22/SUMB[57][51] ) );
  FA_X1 \mult_22/S2_57_50  ( .A(\mult_22/ab[57][50] ), .B(
        \mult_22/CARRYB[56][50] ), .CI(\mult_22/SUMB[56][51] ), .CO(
        \mult_22/CARRYB[57][50] ), .S(\mult_22/SUMB[57][50] ) );
  FA_X1 \mult_22/S2_57_49  ( .A(\mult_22/ab[57][49] ), .B(
        \mult_22/CARRYB[56][49] ), .CI(\mult_22/SUMB[56][50] ), .CO(
        \mult_22/CARRYB[57][49] ), .S(\mult_22/SUMB[57][49] ) );
  FA_X1 \mult_22/S2_57_48  ( .A(\mult_22/ab[57][48] ), .B(
        \mult_22/CARRYB[56][48] ), .CI(\mult_22/SUMB[56][49] ), .CO(
        \mult_22/CARRYB[57][48] ), .S(\mult_22/SUMB[57][48] ) );
  FA_X1 \mult_22/S2_57_47  ( .A(\mult_22/ab[57][47] ), .B(
        \mult_22/CARRYB[56][47] ), .CI(\mult_22/SUMB[56][48] ), .CO(
        \mult_22/CARRYB[57][47] ), .S(\mult_22/SUMB[57][47] ) );
  FA_X1 \mult_22/S2_57_46  ( .A(\mult_22/ab[57][46] ), .B(
        \mult_22/CARRYB[56][46] ), .CI(\mult_22/SUMB[56][47] ), .CO(
        \mult_22/CARRYB[57][46] ), .S(\mult_22/SUMB[57][46] ) );
  FA_X1 \mult_22/S2_57_45  ( .A(\mult_22/ab[57][45] ), .B(
        \mult_22/CARRYB[56][45] ), .CI(\mult_22/SUMB[56][46] ), .CO(
        \mult_22/CARRYB[57][45] ), .S(\mult_22/SUMB[57][45] ) );
  FA_X1 \mult_22/S2_57_44  ( .A(\mult_22/ab[57][44] ), .B(
        \mult_22/CARRYB[56][44] ), .CI(\mult_22/SUMB[56][45] ), .CO(
        \mult_22/CARRYB[57][44] ), .S(\mult_22/SUMB[57][44] ) );
  FA_X1 \mult_22/S2_57_43  ( .A(\mult_22/ab[57][43] ), .B(
        \mult_22/CARRYB[56][43] ), .CI(\mult_22/SUMB[56][44] ), .CO(
        \mult_22/CARRYB[57][43] ), .S(\mult_22/SUMB[57][43] ) );
  FA_X1 \mult_22/S2_57_42  ( .A(\mult_22/ab[57][42] ), .B(
        \mult_22/CARRYB[56][42] ), .CI(\mult_22/SUMB[56][43] ), .CO(
        \mult_22/CARRYB[57][42] ), .S(\mult_22/SUMB[57][42] ) );
  FA_X1 \mult_22/S2_57_41  ( .A(\mult_22/ab[57][41] ), .B(
        \mult_22/CARRYB[56][41] ), .CI(\mult_22/SUMB[56][42] ), .CO(
        \mult_22/CARRYB[57][41] ), .S(\mult_22/SUMB[57][41] ) );
  FA_X1 \mult_22/S2_57_40  ( .A(\mult_22/ab[57][40] ), .B(
        \mult_22/CARRYB[56][40] ), .CI(\mult_22/SUMB[56][41] ), .CO(
        \mult_22/CARRYB[57][40] ), .S(\mult_22/SUMB[57][40] ) );
  FA_X1 \mult_22/S2_57_39  ( .A(\mult_22/ab[57][39] ), .B(
        \mult_22/CARRYB[56][39] ), .CI(\mult_22/SUMB[56][40] ), .CO(
        \mult_22/CARRYB[57][39] ), .S(\mult_22/SUMB[57][39] ) );
  FA_X1 \mult_22/S2_57_38  ( .A(\mult_22/ab[57][38] ), .B(
        \mult_22/CARRYB[56][38] ), .CI(\mult_22/SUMB[56][39] ), .CO(
        \mult_22/CARRYB[57][38] ), .S(\mult_22/SUMB[57][38] ) );
  FA_X1 \mult_22/S2_57_37  ( .A(\mult_22/ab[57][37] ), .B(
        \mult_22/CARRYB[56][37] ), .CI(\mult_22/SUMB[56][38] ), .CO(
        \mult_22/CARRYB[57][37] ), .S(\mult_22/SUMB[57][37] ) );
  FA_X1 \mult_22/S2_57_36  ( .A(\mult_22/ab[57][36] ), .B(
        \mult_22/CARRYB[56][36] ), .CI(\mult_22/SUMB[56][37] ), .CO(
        \mult_22/CARRYB[57][36] ), .S(\mult_22/SUMB[57][36] ) );
  FA_X1 \mult_22/S2_57_35  ( .A(\mult_22/ab[57][35] ), .B(
        \mult_22/CARRYB[56][35] ), .CI(\mult_22/SUMB[56][36] ), .CO(
        \mult_22/CARRYB[57][35] ), .S(\mult_22/SUMB[57][35] ) );
  FA_X1 \mult_22/S2_57_34  ( .A(\mult_22/ab[57][34] ), .B(
        \mult_22/CARRYB[56][34] ), .CI(\mult_22/SUMB[56][35] ), .CO(
        \mult_22/CARRYB[57][34] ), .S(\mult_22/SUMB[57][34] ) );
  FA_X1 \mult_22/S2_57_33  ( .A(\mult_22/ab[57][33] ), .B(
        \mult_22/CARRYB[56][33] ), .CI(\mult_22/SUMB[56][34] ), .CO(
        \mult_22/CARRYB[57][33] ), .S(\mult_22/SUMB[57][33] ) );
  FA_X1 \mult_22/S2_57_32  ( .A(\mult_22/ab[57][32] ), .B(
        \mult_22/CARRYB[56][32] ), .CI(\mult_22/SUMB[56][33] ), .CO(
        \mult_22/CARRYB[57][32] ), .S(\mult_22/SUMB[57][32] ) );
  FA_X1 \mult_22/S2_57_31  ( .A(\mult_22/ab[57][31] ), .B(
        \mult_22/CARRYB[56][31] ), .CI(\mult_22/SUMB[56][32] ), .CO(
        \mult_22/CARRYB[57][31] ), .S(\mult_22/SUMB[57][31] ) );
  FA_X1 \mult_22/S2_57_30  ( .A(\mult_22/ab[57][30] ), .B(
        \mult_22/CARRYB[56][30] ), .CI(\mult_22/SUMB[56][31] ), .CO(
        \mult_22/CARRYB[57][30] ), .S(\mult_22/SUMB[57][30] ) );
  FA_X1 \mult_22/S2_57_29  ( .A(\mult_22/ab[57][29] ), .B(
        \mult_22/CARRYB[56][29] ), .CI(\mult_22/SUMB[56][30] ), .CO(
        \mult_22/CARRYB[57][29] ), .S(\mult_22/SUMB[57][29] ) );
  FA_X1 \mult_22/S2_57_28  ( .A(\mult_22/ab[57][28] ), .B(
        \mult_22/CARRYB[56][28] ), .CI(\mult_22/SUMB[56][29] ), .CO(
        \mult_22/CARRYB[57][28] ), .S(\mult_22/SUMB[57][28] ) );
  FA_X1 \mult_22/S2_57_27  ( .A(\mult_22/ab[57][27] ), .B(
        \mult_22/CARRYB[56][27] ), .CI(\mult_22/SUMB[56][28] ), .CO(
        \mult_22/CARRYB[57][27] ), .S(\mult_22/SUMB[57][27] ) );
  FA_X1 \mult_22/S2_57_26  ( .A(\mult_22/ab[57][26] ), .B(
        \mult_22/CARRYB[56][26] ), .CI(\mult_22/SUMB[56][27] ), .CO(
        \mult_22/CARRYB[57][26] ), .S(\mult_22/SUMB[57][26] ) );
  FA_X1 \mult_22/S2_57_25  ( .A(\mult_22/ab[57][25] ), .B(
        \mult_22/CARRYB[56][25] ), .CI(\mult_22/SUMB[56][26] ), .CO(
        \mult_22/CARRYB[57][25] ), .S(\mult_22/SUMB[57][25] ) );
  FA_X1 \mult_22/S2_57_24  ( .A(\mult_22/ab[57][24] ), .B(
        \mult_22/CARRYB[56][24] ), .CI(\mult_22/SUMB[56][25] ), .CO(
        \mult_22/CARRYB[57][24] ), .S(\mult_22/SUMB[57][24] ) );
  FA_X1 \mult_22/S2_57_23  ( .A(\mult_22/ab[57][23] ), .B(
        \mult_22/CARRYB[56][23] ), .CI(\mult_22/SUMB[56][24] ), .CO(
        \mult_22/CARRYB[57][23] ), .S(\mult_22/SUMB[57][23] ) );
  FA_X1 \mult_22/S2_57_22  ( .A(\mult_22/ab[57][22] ), .B(
        \mult_22/CARRYB[56][22] ), .CI(\mult_22/SUMB[56][23] ), .CO(
        \mult_22/CARRYB[57][22] ), .S(\mult_22/SUMB[57][22] ) );
  FA_X1 \mult_22/S2_57_21  ( .A(\mult_22/ab[57][21] ), .B(
        \mult_22/CARRYB[56][21] ), .CI(\mult_22/SUMB[56][22] ), .CO(
        \mult_22/CARRYB[57][21] ), .S(\mult_22/SUMB[57][21] ) );
  FA_X1 \mult_22/S2_57_20  ( .A(\mult_22/ab[57][20] ), .B(
        \mult_22/CARRYB[56][20] ), .CI(\mult_22/SUMB[56][21] ), .CO(
        \mult_22/CARRYB[57][20] ), .S(\mult_22/SUMB[57][20] ) );
  FA_X1 \mult_22/S2_57_19  ( .A(\mult_22/ab[57][19] ), .B(
        \mult_22/CARRYB[56][19] ), .CI(\mult_22/SUMB[56][20] ), .CO(
        \mult_22/CARRYB[57][19] ), .S(\mult_22/SUMB[57][19] ) );
  FA_X1 \mult_22/S2_57_18  ( .A(\mult_22/ab[57][18] ), .B(
        \mult_22/CARRYB[56][18] ), .CI(\mult_22/SUMB[56][19] ), .CO(
        \mult_22/CARRYB[57][18] ), .S(\mult_22/SUMB[57][18] ) );
  FA_X1 \mult_22/S2_57_17  ( .A(\mult_22/ab[57][17] ), .B(
        \mult_22/CARRYB[56][17] ), .CI(\mult_22/SUMB[56][18] ), .CO(
        \mult_22/CARRYB[57][17] ), .S(\mult_22/SUMB[57][17] ) );
  FA_X1 \mult_22/S2_57_16  ( .A(\mult_22/ab[57][16] ), .B(
        \mult_22/CARRYB[56][16] ), .CI(\mult_22/SUMB[56][17] ), .CO(
        \mult_22/CARRYB[57][16] ), .S(\mult_22/SUMB[57][16] ) );
  FA_X1 \mult_22/S2_57_15  ( .A(\mult_22/ab[57][15] ), .B(
        \mult_22/CARRYB[56][15] ), .CI(\mult_22/SUMB[56][16] ), .CO(
        \mult_22/CARRYB[57][15] ), .S(\mult_22/SUMB[57][15] ) );
  FA_X1 \mult_22/S2_57_14  ( .A(\mult_22/ab[57][14] ), .B(
        \mult_22/CARRYB[56][14] ), .CI(\mult_22/SUMB[56][15] ), .CO(
        \mult_22/CARRYB[57][14] ), .S(\mult_22/SUMB[57][14] ) );
  FA_X1 \mult_22/S2_57_13  ( .A(\mult_22/ab[57][13] ), .B(
        \mult_22/CARRYB[56][13] ), .CI(\mult_22/SUMB[56][14] ), .CO(
        \mult_22/CARRYB[57][13] ), .S(\mult_22/SUMB[57][13] ) );
  FA_X1 \mult_22/S2_57_12  ( .A(\mult_22/ab[57][12] ), .B(
        \mult_22/CARRYB[56][12] ), .CI(\mult_22/SUMB[56][13] ), .CO(
        \mult_22/CARRYB[57][12] ), .S(\mult_22/SUMB[57][12] ) );
  FA_X1 \mult_22/S2_57_11  ( .A(\mult_22/ab[57][11] ), .B(
        \mult_22/CARRYB[56][11] ), .CI(\mult_22/SUMB[56][12] ), .CO(
        \mult_22/CARRYB[57][11] ), .S(\mult_22/SUMB[57][11] ) );
  FA_X1 \mult_22/S2_57_10  ( .A(\mult_22/CARRYB[56][10] ), .B(
        \mult_22/ab[57][10] ), .CI(\mult_22/SUMB[56][11] ), .CO(
        \mult_22/CARRYB[57][10] ), .S(\mult_22/SUMB[57][10] ) );
  FA_X1 \mult_22/S2_57_9  ( .A(\mult_22/CARRYB[56][9] ), .B(
        \mult_22/ab[57][9] ), .CI(\mult_22/SUMB[56][10] ), .CO(
        \mult_22/CARRYB[57][9] ), .S(\mult_22/SUMB[57][9] ) );
  FA_X1 \mult_22/S2_57_8  ( .A(\mult_22/ab[57][8] ), .B(
        \mult_22/CARRYB[56][8] ), .CI(\mult_22/SUMB[56][9] ), .CO(
        \mult_22/CARRYB[57][8] ), .S(\mult_22/SUMB[57][8] ) );
  FA_X1 \mult_22/S2_57_7  ( .A(\mult_22/CARRYB[56][7] ), .B(
        \mult_22/ab[57][7] ), .CI(\mult_22/SUMB[56][8] ), .CO(
        \mult_22/CARRYB[57][7] ), .S(\mult_22/SUMB[57][7] ) );
  FA_X1 \mult_22/S2_57_6  ( .A(\mult_22/ab[57][6] ), .B(
        \mult_22/CARRYB[56][6] ), .CI(\mult_22/SUMB[56][7] ), .CO(
        \mult_22/CARRYB[57][6] ), .S(\mult_22/SUMB[57][6] ) );
  FA_X1 \mult_22/S2_57_5  ( .A(\mult_22/ab[57][5] ), .B(
        \mult_22/CARRYB[56][5] ), .CI(\mult_22/SUMB[56][6] ), .CO(
        \mult_22/CARRYB[57][5] ), .S(\mult_22/SUMB[57][5] ) );
  FA_X1 \mult_22/S2_57_4  ( .A(\mult_22/ab[57][4] ), .B(
        \mult_22/CARRYB[56][4] ), .CI(\mult_22/SUMB[56][5] ), .CO(
        \mult_22/CARRYB[57][4] ), .S(\mult_22/SUMB[57][4] ) );
  FA_X1 \mult_22/S2_57_3  ( .A(\mult_22/ab[57][3] ), .B(
        \mult_22/CARRYB[56][3] ), .CI(\mult_22/SUMB[56][4] ), .CO(
        \mult_22/CARRYB[57][3] ), .S(\mult_22/SUMB[57][3] ) );
  FA_X1 \mult_22/S2_57_2  ( .A(\mult_22/ab[57][2] ), .B(
        \mult_22/CARRYB[56][2] ), .CI(\mult_22/SUMB[56][3] ), .CO(
        \mult_22/CARRYB[57][2] ), .S(\mult_22/SUMB[57][2] ) );
  FA_X1 \mult_22/S2_57_1  ( .A(\mult_22/ab[57][1] ), .B(
        \mult_22/CARRYB[56][1] ), .CI(\mult_22/SUMB[56][2] ), .CO(
        \mult_22/CARRYB[57][1] ), .S(\mult_22/SUMB[57][1] ) );
  FA_X1 \mult_22/S1_57_0  ( .A(\mult_22/ab[57][0] ), .B(
        \mult_22/CARRYB[56][0] ), .CI(\mult_22/SUMB[56][1] ), .CO(
        \mult_22/CARRYB[57][0] ), .S(N185) );
  FA_X1 \mult_22/S3_58_62  ( .A(\mult_22/ab[58][62] ), .B(
        \mult_22/CARRYB[57][62] ), .CI(\mult_22/ab[57][63] ), .CO(
        \mult_22/CARRYB[58][62] ), .S(\mult_22/SUMB[58][62] ) );
  FA_X1 \mult_22/S2_58_61  ( .A(\mult_22/ab[58][61] ), .B(
        \mult_22/CARRYB[57][61] ), .CI(\mult_22/SUMB[57][62] ), .CO(
        \mult_22/CARRYB[58][61] ), .S(\mult_22/SUMB[58][61] ) );
  FA_X1 \mult_22/S2_58_60  ( .A(\mult_22/ab[58][60] ), .B(
        \mult_22/CARRYB[57][60] ), .CI(\mult_22/SUMB[57][61] ), .CO(
        \mult_22/CARRYB[58][60] ), .S(\mult_22/SUMB[58][60] ) );
  FA_X1 \mult_22/S2_58_59  ( .A(\mult_22/ab[58][59] ), .B(
        \mult_22/CARRYB[57][59] ), .CI(\mult_22/SUMB[57][60] ), .CO(
        \mult_22/CARRYB[58][59] ), .S(\mult_22/SUMB[58][59] ) );
  FA_X1 \mult_22/S2_58_58  ( .A(\mult_22/ab[58][58] ), .B(
        \mult_22/CARRYB[57][58] ), .CI(\mult_22/SUMB[57][59] ), .CO(
        \mult_22/CARRYB[58][58] ), .S(\mult_22/SUMB[58][58] ) );
  FA_X1 \mult_22/S2_58_57  ( .A(\mult_22/ab[58][57] ), .B(
        \mult_22/CARRYB[57][57] ), .CI(\mult_22/SUMB[57][58] ), .CO(
        \mult_22/CARRYB[58][57] ), .S(\mult_22/SUMB[58][57] ) );
  FA_X1 \mult_22/S2_58_56  ( .A(\mult_22/ab[58][56] ), .B(
        \mult_22/CARRYB[57][56] ), .CI(\mult_22/SUMB[57][57] ), .CO(
        \mult_22/CARRYB[58][56] ), .S(\mult_22/SUMB[58][56] ) );
  FA_X1 \mult_22/S2_58_55  ( .A(\mult_22/ab[58][55] ), .B(
        \mult_22/CARRYB[57][55] ), .CI(\mult_22/SUMB[57][56] ), .CO(
        \mult_22/CARRYB[58][55] ), .S(\mult_22/SUMB[58][55] ) );
  FA_X1 \mult_22/S2_58_54  ( .A(\mult_22/ab[58][54] ), .B(
        \mult_22/CARRYB[57][54] ), .CI(\mult_22/SUMB[57][55] ), .CO(
        \mult_22/CARRYB[58][54] ), .S(\mult_22/SUMB[58][54] ) );
  FA_X1 \mult_22/S2_58_53  ( .A(\mult_22/ab[58][53] ), .B(
        \mult_22/CARRYB[57][53] ), .CI(\mult_22/SUMB[57][54] ), .CO(
        \mult_22/CARRYB[58][53] ), .S(\mult_22/SUMB[58][53] ) );
  FA_X1 \mult_22/S2_58_52  ( .A(\mult_22/ab[58][52] ), .B(
        \mult_22/CARRYB[57][52] ), .CI(\mult_22/SUMB[57][53] ), .CO(
        \mult_22/CARRYB[58][52] ), .S(\mult_22/SUMB[58][52] ) );
  FA_X1 \mult_22/S2_58_51  ( .A(\mult_22/ab[58][51] ), .B(
        \mult_22/CARRYB[57][51] ), .CI(\mult_22/SUMB[57][52] ), .CO(
        \mult_22/CARRYB[58][51] ), .S(\mult_22/SUMB[58][51] ) );
  FA_X1 \mult_22/S2_58_50  ( .A(\mult_22/ab[58][50] ), .B(
        \mult_22/CARRYB[57][50] ), .CI(\mult_22/SUMB[57][51] ), .CO(
        \mult_22/CARRYB[58][50] ), .S(\mult_22/SUMB[58][50] ) );
  FA_X1 \mult_22/S2_58_49  ( .A(\mult_22/ab[58][49] ), .B(
        \mult_22/CARRYB[57][49] ), .CI(\mult_22/SUMB[57][50] ), .CO(
        \mult_22/CARRYB[58][49] ), .S(\mult_22/SUMB[58][49] ) );
  FA_X1 \mult_22/S2_58_48  ( .A(\mult_22/ab[58][48] ), .B(
        \mult_22/CARRYB[57][48] ), .CI(\mult_22/SUMB[57][49] ), .CO(
        \mult_22/CARRYB[58][48] ), .S(\mult_22/SUMB[58][48] ) );
  FA_X1 \mult_22/S2_58_47  ( .A(\mult_22/ab[58][47] ), .B(
        \mult_22/CARRYB[57][47] ), .CI(\mult_22/SUMB[57][48] ), .CO(
        \mult_22/CARRYB[58][47] ), .S(\mult_22/SUMB[58][47] ) );
  FA_X1 \mult_22/S2_58_46  ( .A(\mult_22/ab[58][46] ), .B(
        \mult_22/CARRYB[57][46] ), .CI(\mult_22/SUMB[57][47] ), .CO(
        \mult_22/CARRYB[58][46] ), .S(\mult_22/SUMB[58][46] ) );
  FA_X1 \mult_22/S2_58_45  ( .A(\mult_22/ab[58][45] ), .B(
        \mult_22/CARRYB[57][45] ), .CI(\mult_22/SUMB[57][46] ), .CO(
        \mult_22/CARRYB[58][45] ), .S(\mult_22/SUMB[58][45] ) );
  FA_X1 \mult_22/S2_58_44  ( .A(\mult_22/ab[58][44] ), .B(
        \mult_22/CARRYB[57][44] ), .CI(\mult_22/SUMB[57][45] ), .CO(
        \mult_22/CARRYB[58][44] ), .S(\mult_22/SUMB[58][44] ) );
  FA_X1 \mult_22/S2_58_43  ( .A(\mult_22/ab[58][43] ), .B(
        \mult_22/CARRYB[57][43] ), .CI(\mult_22/SUMB[57][44] ), .CO(
        \mult_22/CARRYB[58][43] ), .S(\mult_22/SUMB[58][43] ) );
  FA_X1 \mult_22/S2_58_42  ( .A(\mult_22/ab[58][42] ), .B(
        \mult_22/CARRYB[57][42] ), .CI(\mult_22/SUMB[57][43] ), .CO(
        \mult_22/CARRYB[58][42] ), .S(\mult_22/SUMB[58][42] ) );
  FA_X1 \mult_22/S2_58_41  ( .A(\mult_22/ab[58][41] ), .B(
        \mult_22/CARRYB[57][41] ), .CI(\mult_22/SUMB[57][42] ), .CO(
        \mult_22/CARRYB[58][41] ), .S(\mult_22/SUMB[58][41] ) );
  FA_X1 \mult_22/S2_58_40  ( .A(\mult_22/ab[58][40] ), .B(
        \mult_22/CARRYB[57][40] ), .CI(\mult_22/SUMB[57][41] ), .CO(
        \mult_22/CARRYB[58][40] ), .S(\mult_22/SUMB[58][40] ) );
  FA_X1 \mult_22/S2_58_39  ( .A(\mult_22/ab[58][39] ), .B(
        \mult_22/CARRYB[57][39] ), .CI(\mult_22/SUMB[57][40] ), .CO(
        \mult_22/CARRYB[58][39] ), .S(\mult_22/SUMB[58][39] ) );
  FA_X1 \mult_22/S2_58_38  ( .A(\mult_22/ab[58][38] ), .B(
        \mult_22/CARRYB[57][38] ), .CI(\mult_22/SUMB[57][39] ), .CO(
        \mult_22/CARRYB[58][38] ), .S(\mult_22/SUMB[58][38] ) );
  FA_X1 \mult_22/S2_58_37  ( .A(\mult_22/ab[58][37] ), .B(
        \mult_22/CARRYB[57][37] ), .CI(\mult_22/SUMB[57][38] ), .CO(
        \mult_22/CARRYB[58][37] ), .S(\mult_22/SUMB[58][37] ) );
  FA_X1 \mult_22/S2_58_36  ( .A(\mult_22/ab[58][36] ), .B(
        \mult_22/CARRYB[57][36] ), .CI(\mult_22/SUMB[57][37] ), .CO(
        \mult_22/CARRYB[58][36] ), .S(\mult_22/SUMB[58][36] ) );
  FA_X1 \mult_22/S2_58_35  ( .A(\mult_22/ab[58][35] ), .B(
        \mult_22/CARRYB[57][35] ), .CI(\mult_22/SUMB[57][36] ), .CO(
        \mult_22/CARRYB[58][35] ), .S(\mult_22/SUMB[58][35] ) );
  FA_X1 \mult_22/S2_58_34  ( .A(\mult_22/ab[58][34] ), .B(
        \mult_22/CARRYB[57][34] ), .CI(\mult_22/SUMB[57][35] ), .CO(
        \mult_22/CARRYB[58][34] ), .S(\mult_22/SUMB[58][34] ) );
  FA_X1 \mult_22/S2_58_33  ( .A(\mult_22/ab[58][33] ), .B(
        \mult_22/CARRYB[57][33] ), .CI(\mult_22/SUMB[57][34] ), .CO(
        \mult_22/CARRYB[58][33] ), .S(\mult_22/SUMB[58][33] ) );
  FA_X1 \mult_22/S2_58_32  ( .A(\mult_22/ab[58][32] ), .B(
        \mult_22/CARRYB[57][32] ), .CI(\mult_22/SUMB[57][33] ), .CO(
        \mult_22/CARRYB[58][32] ), .S(\mult_22/SUMB[58][32] ) );
  FA_X1 \mult_22/S2_58_31  ( .A(\mult_22/ab[58][31] ), .B(
        \mult_22/CARRYB[57][31] ), .CI(\mult_22/SUMB[57][32] ), .CO(
        \mult_22/CARRYB[58][31] ), .S(\mult_22/SUMB[58][31] ) );
  FA_X1 \mult_22/S2_58_30  ( .A(\mult_22/ab[58][30] ), .B(
        \mult_22/CARRYB[57][30] ), .CI(\mult_22/SUMB[57][31] ), .CO(
        \mult_22/CARRYB[58][30] ), .S(\mult_22/SUMB[58][30] ) );
  FA_X1 \mult_22/S2_58_29  ( .A(\mult_22/ab[58][29] ), .B(
        \mult_22/CARRYB[57][29] ), .CI(\mult_22/SUMB[57][30] ), .CO(
        \mult_22/CARRYB[58][29] ), .S(\mult_22/SUMB[58][29] ) );
  FA_X1 \mult_22/S2_58_28  ( .A(\mult_22/ab[58][28] ), .B(
        \mult_22/CARRYB[57][28] ), .CI(\mult_22/SUMB[57][29] ), .CO(
        \mult_22/CARRYB[58][28] ), .S(\mult_22/SUMB[58][28] ) );
  FA_X1 \mult_22/S2_58_27  ( .A(\mult_22/ab[58][27] ), .B(
        \mult_22/CARRYB[57][27] ), .CI(\mult_22/SUMB[57][28] ), .CO(
        \mult_22/CARRYB[58][27] ), .S(\mult_22/SUMB[58][27] ) );
  FA_X1 \mult_22/S2_58_26  ( .A(\mult_22/ab[58][26] ), .B(
        \mult_22/CARRYB[57][26] ), .CI(\mult_22/SUMB[57][27] ), .CO(
        \mult_22/CARRYB[58][26] ), .S(\mult_22/SUMB[58][26] ) );
  FA_X1 \mult_22/S2_58_25  ( .A(\mult_22/ab[58][25] ), .B(
        \mult_22/CARRYB[57][25] ), .CI(\mult_22/SUMB[57][26] ), .CO(
        \mult_22/CARRYB[58][25] ), .S(\mult_22/SUMB[58][25] ) );
  FA_X1 \mult_22/S2_58_24  ( .A(\mult_22/ab[58][24] ), .B(
        \mult_22/CARRYB[57][24] ), .CI(\mult_22/SUMB[57][25] ), .CO(
        \mult_22/CARRYB[58][24] ), .S(\mult_22/SUMB[58][24] ) );
  FA_X1 \mult_22/S2_58_23  ( .A(\mult_22/ab[58][23] ), .B(
        \mult_22/CARRYB[57][23] ), .CI(\mult_22/SUMB[57][24] ), .CO(
        \mult_22/CARRYB[58][23] ), .S(\mult_22/SUMB[58][23] ) );
  FA_X1 \mult_22/S2_58_22  ( .A(\mult_22/ab[58][22] ), .B(
        \mult_22/CARRYB[57][22] ), .CI(\mult_22/SUMB[57][23] ), .CO(
        \mult_22/CARRYB[58][22] ), .S(\mult_22/SUMB[58][22] ) );
  FA_X1 \mult_22/S2_58_21  ( .A(\mult_22/ab[58][21] ), .B(
        \mult_22/CARRYB[57][21] ), .CI(\mult_22/SUMB[57][22] ), .CO(
        \mult_22/CARRYB[58][21] ), .S(\mult_22/SUMB[58][21] ) );
  FA_X1 \mult_22/S2_58_20  ( .A(\mult_22/ab[58][20] ), .B(
        \mult_22/CARRYB[57][20] ), .CI(\mult_22/SUMB[57][21] ), .CO(
        \mult_22/CARRYB[58][20] ), .S(\mult_22/SUMB[58][20] ) );
  FA_X1 \mult_22/S2_58_19  ( .A(\mult_22/ab[58][19] ), .B(
        \mult_22/CARRYB[57][19] ), .CI(\mult_22/SUMB[57][20] ), .CO(
        \mult_22/CARRYB[58][19] ), .S(\mult_22/SUMB[58][19] ) );
  FA_X1 \mult_22/S2_58_18  ( .A(\mult_22/ab[58][18] ), .B(
        \mult_22/CARRYB[57][18] ), .CI(\mult_22/SUMB[57][19] ), .CO(
        \mult_22/CARRYB[58][18] ), .S(\mult_22/SUMB[58][18] ) );
  FA_X1 \mult_22/S2_58_17  ( .A(\mult_22/ab[58][17] ), .B(
        \mult_22/CARRYB[57][17] ), .CI(\mult_22/SUMB[57][18] ), .CO(
        \mult_22/CARRYB[58][17] ), .S(\mult_22/SUMB[58][17] ) );
  FA_X1 \mult_22/S2_58_16  ( .A(\mult_22/ab[58][16] ), .B(
        \mult_22/CARRYB[57][16] ), .CI(\mult_22/SUMB[57][17] ), .CO(
        \mult_22/CARRYB[58][16] ), .S(\mult_22/SUMB[58][16] ) );
  FA_X1 \mult_22/S2_58_15  ( .A(\mult_22/ab[58][15] ), .B(
        \mult_22/CARRYB[57][15] ), .CI(\mult_22/SUMB[57][16] ), .CO(
        \mult_22/CARRYB[58][15] ), .S(\mult_22/SUMB[58][15] ) );
  FA_X1 \mult_22/S2_58_14  ( .A(\mult_22/ab[58][14] ), .B(
        \mult_22/CARRYB[57][14] ), .CI(\mult_22/SUMB[57][15] ), .CO(
        \mult_22/CARRYB[58][14] ), .S(\mult_22/SUMB[58][14] ) );
  FA_X1 \mult_22/S2_58_13  ( .A(\mult_22/ab[58][13] ), .B(
        \mult_22/CARRYB[57][13] ), .CI(\mult_22/SUMB[57][14] ), .CO(
        \mult_22/CARRYB[58][13] ), .S(\mult_22/SUMB[58][13] ) );
  FA_X1 \mult_22/S2_58_12  ( .A(\mult_22/ab[58][12] ), .B(
        \mult_22/CARRYB[57][12] ), .CI(\mult_22/SUMB[57][13] ), .CO(
        \mult_22/CARRYB[58][12] ), .S(\mult_22/SUMB[58][12] ) );
  FA_X1 \mult_22/S2_58_11  ( .A(\mult_22/ab[58][11] ), .B(
        \mult_22/CARRYB[57][11] ), .CI(\mult_22/SUMB[57][12] ), .CO(
        \mult_22/CARRYB[58][11] ), .S(\mult_22/SUMB[58][11] ) );
  FA_X1 \mult_22/S2_58_10  ( .A(\mult_22/ab[58][10] ), .B(
        \mult_22/CARRYB[57][10] ), .CI(\mult_22/SUMB[57][11] ), .CO(
        \mult_22/CARRYB[58][10] ), .S(\mult_22/SUMB[58][10] ) );
  FA_X1 \mult_22/S2_58_9  ( .A(\mult_22/ab[58][9] ), .B(
        \mult_22/CARRYB[57][9] ), .CI(\mult_22/SUMB[57][10] ), .CO(
        \mult_22/CARRYB[58][9] ), .S(\mult_22/SUMB[58][9] ) );
  FA_X1 \mult_22/S2_58_8  ( .A(\mult_22/CARRYB[57][8] ), .B(
        \mult_22/ab[58][8] ), .CI(\mult_22/SUMB[57][9] ), .CO(
        \mult_22/CARRYB[58][8] ), .S(\mult_22/SUMB[58][8] ) );
  FA_X1 \mult_22/S2_58_7  ( .A(\mult_22/CARRYB[57][7] ), .B(
        \mult_22/ab[58][7] ), .CI(\mult_22/SUMB[57][8] ), .CO(
        \mult_22/CARRYB[58][7] ), .S(\mult_22/SUMB[58][7] ) );
  FA_X1 \mult_22/S2_58_6  ( .A(\mult_22/ab[58][6] ), .B(
        \mult_22/CARRYB[57][6] ), .CI(\mult_22/SUMB[57][7] ), .CO(
        \mult_22/CARRYB[58][6] ), .S(\mult_22/SUMB[58][6] ) );
  FA_X1 \mult_22/S2_58_5  ( .A(\mult_22/ab[58][5] ), .B(
        \mult_22/CARRYB[57][5] ), .CI(\mult_22/SUMB[57][6] ), .CO(
        \mult_22/CARRYB[58][5] ), .S(\mult_22/SUMB[58][5] ) );
  FA_X1 \mult_22/S2_58_4  ( .A(\mult_22/ab[58][4] ), .B(
        \mult_22/CARRYB[57][4] ), .CI(\mult_22/SUMB[57][5] ), .CO(
        \mult_22/CARRYB[58][4] ), .S(\mult_22/SUMB[58][4] ) );
  FA_X1 \mult_22/S2_58_3  ( .A(\mult_22/ab[58][3] ), .B(
        \mult_22/CARRYB[57][3] ), .CI(\mult_22/SUMB[57][4] ), .CO(
        \mult_22/CARRYB[58][3] ), .S(\mult_22/SUMB[58][3] ) );
  FA_X1 \mult_22/S2_58_2  ( .A(\mult_22/ab[58][2] ), .B(
        \mult_22/CARRYB[57][2] ), .CI(\mult_22/SUMB[57][3] ), .CO(
        \mult_22/CARRYB[58][2] ), .S(\mult_22/SUMB[58][2] ) );
  FA_X1 \mult_22/S2_58_1  ( .A(\mult_22/ab[58][1] ), .B(
        \mult_22/CARRYB[57][1] ), .CI(\mult_22/SUMB[57][2] ), .CO(
        \mult_22/CARRYB[58][1] ), .S(\mult_22/SUMB[58][1] ) );
  FA_X1 \mult_22/S1_58_0  ( .A(\mult_22/ab[58][0] ), .B(
        \mult_22/CARRYB[57][0] ), .CI(\mult_22/SUMB[57][1] ), .CO(
        \mult_22/CARRYB[58][0] ), .S(N186) );
  FA_X1 \mult_22/S3_59_62  ( .A(\mult_22/ab[59][62] ), .B(
        \mult_22/CARRYB[58][62] ), .CI(\mult_22/ab[58][63] ), .CO(
        \mult_22/CARRYB[59][62] ), .S(\mult_22/SUMB[59][62] ) );
  FA_X1 \mult_22/S2_59_61  ( .A(\mult_22/ab[59][61] ), .B(
        \mult_22/CARRYB[58][61] ), .CI(\mult_22/SUMB[58][62] ), .CO(
        \mult_22/CARRYB[59][61] ), .S(\mult_22/SUMB[59][61] ) );
  FA_X1 \mult_22/S2_59_60  ( .A(\mult_22/ab[59][60] ), .B(
        \mult_22/CARRYB[58][60] ), .CI(\mult_22/SUMB[58][61] ), .CO(
        \mult_22/CARRYB[59][60] ), .S(\mult_22/SUMB[59][60] ) );
  FA_X1 \mult_22/S2_59_59  ( .A(\mult_22/ab[59][59] ), .B(
        \mult_22/CARRYB[58][59] ), .CI(\mult_22/SUMB[58][60] ), .CO(
        \mult_22/CARRYB[59][59] ), .S(\mult_22/SUMB[59][59] ) );
  FA_X1 \mult_22/S2_59_58  ( .A(\mult_22/ab[59][58] ), .B(
        \mult_22/CARRYB[58][58] ), .CI(\mult_22/SUMB[58][59] ), .CO(
        \mult_22/CARRYB[59][58] ), .S(\mult_22/SUMB[59][58] ) );
  FA_X1 \mult_22/S2_59_57  ( .A(\mult_22/ab[59][57] ), .B(
        \mult_22/CARRYB[58][57] ), .CI(\mult_22/SUMB[58][58] ), .CO(
        \mult_22/CARRYB[59][57] ), .S(\mult_22/SUMB[59][57] ) );
  FA_X1 \mult_22/S2_59_56  ( .A(\mult_22/ab[59][56] ), .B(
        \mult_22/CARRYB[58][56] ), .CI(\mult_22/SUMB[58][57] ), .CO(
        \mult_22/CARRYB[59][56] ), .S(\mult_22/SUMB[59][56] ) );
  FA_X1 \mult_22/S2_59_55  ( .A(\mult_22/ab[59][55] ), .B(
        \mult_22/CARRYB[58][55] ), .CI(\mult_22/SUMB[58][56] ), .CO(
        \mult_22/CARRYB[59][55] ), .S(\mult_22/SUMB[59][55] ) );
  FA_X1 \mult_22/S2_59_54  ( .A(\mult_22/ab[59][54] ), .B(
        \mult_22/CARRYB[58][54] ), .CI(\mult_22/SUMB[58][55] ), .CO(
        \mult_22/CARRYB[59][54] ), .S(\mult_22/SUMB[59][54] ) );
  FA_X1 \mult_22/S2_59_53  ( .A(\mult_22/ab[59][53] ), .B(
        \mult_22/CARRYB[58][53] ), .CI(\mult_22/SUMB[58][54] ), .CO(
        \mult_22/CARRYB[59][53] ), .S(\mult_22/SUMB[59][53] ) );
  FA_X1 \mult_22/S2_59_52  ( .A(\mult_22/ab[59][52] ), .B(
        \mult_22/CARRYB[58][52] ), .CI(\mult_22/SUMB[58][53] ), .CO(
        \mult_22/CARRYB[59][52] ), .S(\mult_22/SUMB[59][52] ) );
  FA_X1 \mult_22/S2_59_51  ( .A(\mult_22/ab[59][51] ), .B(
        \mult_22/CARRYB[58][51] ), .CI(\mult_22/SUMB[58][52] ), .CO(
        \mult_22/CARRYB[59][51] ), .S(\mult_22/SUMB[59][51] ) );
  FA_X1 \mult_22/S2_59_50  ( .A(\mult_22/ab[59][50] ), .B(
        \mult_22/CARRYB[58][50] ), .CI(\mult_22/SUMB[58][51] ), .CO(
        \mult_22/CARRYB[59][50] ), .S(\mult_22/SUMB[59][50] ) );
  FA_X1 \mult_22/S2_59_49  ( .A(\mult_22/ab[59][49] ), .B(
        \mult_22/CARRYB[58][49] ), .CI(\mult_22/SUMB[58][50] ), .CO(
        \mult_22/CARRYB[59][49] ), .S(\mult_22/SUMB[59][49] ) );
  FA_X1 \mult_22/S2_59_48  ( .A(\mult_22/ab[59][48] ), .B(
        \mult_22/CARRYB[58][48] ), .CI(\mult_22/SUMB[58][49] ), .CO(
        \mult_22/CARRYB[59][48] ), .S(\mult_22/SUMB[59][48] ) );
  FA_X1 \mult_22/S2_59_47  ( .A(\mult_22/ab[59][47] ), .B(
        \mult_22/CARRYB[58][47] ), .CI(\mult_22/SUMB[58][48] ), .CO(
        \mult_22/CARRYB[59][47] ), .S(\mult_22/SUMB[59][47] ) );
  FA_X1 \mult_22/S2_59_46  ( .A(\mult_22/ab[59][46] ), .B(
        \mult_22/CARRYB[58][46] ), .CI(\mult_22/SUMB[58][47] ), .CO(
        \mult_22/CARRYB[59][46] ), .S(\mult_22/SUMB[59][46] ) );
  FA_X1 \mult_22/S2_59_45  ( .A(\mult_22/ab[59][45] ), .B(
        \mult_22/CARRYB[58][45] ), .CI(\mult_22/SUMB[58][46] ), .CO(
        \mult_22/CARRYB[59][45] ), .S(\mult_22/SUMB[59][45] ) );
  FA_X1 \mult_22/S2_59_44  ( .A(\mult_22/ab[59][44] ), .B(
        \mult_22/CARRYB[58][44] ), .CI(\mult_22/SUMB[58][45] ), .CO(
        \mult_22/CARRYB[59][44] ), .S(\mult_22/SUMB[59][44] ) );
  FA_X1 \mult_22/S2_59_43  ( .A(\mult_22/ab[59][43] ), .B(
        \mult_22/CARRYB[58][43] ), .CI(\mult_22/SUMB[58][44] ), .CO(
        \mult_22/CARRYB[59][43] ), .S(\mult_22/SUMB[59][43] ) );
  FA_X1 \mult_22/S2_59_42  ( .A(\mult_22/ab[59][42] ), .B(
        \mult_22/CARRYB[58][42] ), .CI(\mult_22/SUMB[58][43] ), .CO(
        \mult_22/CARRYB[59][42] ), .S(\mult_22/SUMB[59][42] ) );
  FA_X1 \mult_22/S2_59_41  ( .A(\mult_22/ab[59][41] ), .B(
        \mult_22/CARRYB[58][41] ), .CI(\mult_22/SUMB[58][42] ), .CO(
        \mult_22/CARRYB[59][41] ), .S(\mult_22/SUMB[59][41] ) );
  FA_X1 \mult_22/S2_59_40  ( .A(\mult_22/ab[59][40] ), .B(
        \mult_22/CARRYB[58][40] ), .CI(\mult_22/SUMB[58][41] ), .CO(
        \mult_22/CARRYB[59][40] ), .S(\mult_22/SUMB[59][40] ) );
  FA_X1 \mult_22/S2_59_39  ( .A(\mult_22/ab[59][39] ), .B(
        \mult_22/CARRYB[58][39] ), .CI(\mult_22/SUMB[58][40] ), .CO(
        \mult_22/CARRYB[59][39] ), .S(\mult_22/SUMB[59][39] ) );
  FA_X1 \mult_22/S2_59_38  ( .A(\mult_22/ab[59][38] ), .B(
        \mult_22/CARRYB[58][38] ), .CI(\mult_22/SUMB[58][39] ), .CO(
        \mult_22/CARRYB[59][38] ), .S(\mult_22/SUMB[59][38] ) );
  FA_X1 \mult_22/S2_59_37  ( .A(\mult_22/ab[59][37] ), .B(
        \mult_22/CARRYB[58][37] ), .CI(\mult_22/SUMB[58][38] ), .CO(
        \mult_22/CARRYB[59][37] ), .S(\mult_22/SUMB[59][37] ) );
  FA_X1 \mult_22/S2_59_36  ( .A(\mult_22/ab[59][36] ), .B(
        \mult_22/CARRYB[58][36] ), .CI(\mult_22/SUMB[58][37] ), .CO(
        \mult_22/CARRYB[59][36] ), .S(\mult_22/SUMB[59][36] ) );
  FA_X1 \mult_22/S2_59_35  ( .A(\mult_22/ab[59][35] ), .B(
        \mult_22/CARRYB[58][35] ), .CI(\mult_22/SUMB[58][36] ), .CO(
        \mult_22/CARRYB[59][35] ), .S(\mult_22/SUMB[59][35] ) );
  FA_X1 \mult_22/S2_59_34  ( .A(\mult_22/ab[59][34] ), .B(
        \mult_22/CARRYB[58][34] ), .CI(\mult_22/SUMB[58][35] ), .CO(
        \mult_22/CARRYB[59][34] ), .S(\mult_22/SUMB[59][34] ) );
  FA_X1 \mult_22/S2_59_33  ( .A(\mult_22/ab[59][33] ), .B(
        \mult_22/CARRYB[58][33] ), .CI(\mult_22/SUMB[58][34] ), .CO(
        \mult_22/CARRYB[59][33] ), .S(\mult_22/SUMB[59][33] ) );
  FA_X1 \mult_22/S2_59_32  ( .A(\mult_22/ab[59][32] ), .B(
        \mult_22/CARRYB[58][32] ), .CI(\mult_22/SUMB[58][33] ), .CO(
        \mult_22/CARRYB[59][32] ), .S(\mult_22/SUMB[59][32] ) );
  FA_X1 \mult_22/S2_59_31  ( .A(\mult_22/ab[59][31] ), .B(
        \mult_22/CARRYB[58][31] ), .CI(\mult_22/SUMB[58][32] ), .CO(
        \mult_22/CARRYB[59][31] ), .S(\mult_22/SUMB[59][31] ) );
  FA_X1 \mult_22/S2_59_30  ( .A(\mult_22/ab[59][30] ), .B(
        \mult_22/CARRYB[58][30] ), .CI(\mult_22/SUMB[58][31] ), .CO(
        \mult_22/CARRYB[59][30] ), .S(\mult_22/SUMB[59][30] ) );
  FA_X1 \mult_22/S2_59_29  ( .A(\mult_22/ab[59][29] ), .B(
        \mult_22/CARRYB[58][29] ), .CI(\mult_22/SUMB[58][30] ), .CO(
        \mult_22/CARRYB[59][29] ), .S(\mult_22/SUMB[59][29] ) );
  FA_X1 \mult_22/S2_59_28  ( .A(\mult_22/ab[59][28] ), .B(
        \mult_22/CARRYB[58][28] ), .CI(\mult_22/SUMB[58][29] ), .CO(
        \mult_22/CARRYB[59][28] ), .S(\mult_22/SUMB[59][28] ) );
  FA_X1 \mult_22/S2_59_27  ( .A(\mult_22/ab[59][27] ), .B(
        \mult_22/CARRYB[58][27] ), .CI(\mult_22/SUMB[58][28] ), .CO(
        \mult_22/CARRYB[59][27] ), .S(\mult_22/SUMB[59][27] ) );
  FA_X1 \mult_22/S2_59_26  ( .A(\mult_22/ab[59][26] ), .B(
        \mult_22/CARRYB[58][26] ), .CI(\mult_22/SUMB[58][27] ), .CO(
        \mult_22/CARRYB[59][26] ), .S(\mult_22/SUMB[59][26] ) );
  FA_X1 \mult_22/S2_59_25  ( .A(\mult_22/ab[59][25] ), .B(
        \mult_22/CARRYB[58][25] ), .CI(\mult_22/SUMB[58][26] ), .CO(
        \mult_22/CARRYB[59][25] ), .S(\mult_22/SUMB[59][25] ) );
  FA_X1 \mult_22/S2_59_24  ( .A(\mult_22/ab[59][24] ), .B(
        \mult_22/CARRYB[58][24] ), .CI(\mult_22/SUMB[58][25] ), .CO(
        \mult_22/CARRYB[59][24] ), .S(\mult_22/SUMB[59][24] ) );
  FA_X1 \mult_22/S2_59_23  ( .A(\mult_22/ab[59][23] ), .B(
        \mult_22/CARRYB[58][23] ), .CI(\mult_22/SUMB[58][24] ), .CO(
        \mult_22/CARRYB[59][23] ), .S(\mult_22/SUMB[59][23] ) );
  FA_X1 \mult_22/S2_59_22  ( .A(\mult_22/ab[59][22] ), .B(
        \mult_22/CARRYB[58][22] ), .CI(\mult_22/SUMB[58][23] ), .CO(
        \mult_22/CARRYB[59][22] ), .S(\mult_22/SUMB[59][22] ) );
  FA_X1 \mult_22/S2_59_21  ( .A(\mult_22/ab[59][21] ), .B(
        \mult_22/CARRYB[58][21] ), .CI(\mult_22/SUMB[58][22] ), .CO(
        \mult_22/CARRYB[59][21] ), .S(\mult_22/SUMB[59][21] ) );
  FA_X1 \mult_22/S2_59_20  ( .A(\mult_22/ab[59][20] ), .B(
        \mult_22/CARRYB[58][20] ), .CI(\mult_22/SUMB[58][21] ), .CO(
        \mult_22/CARRYB[59][20] ), .S(\mult_22/SUMB[59][20] ) );
  FA_X1 \mult_22/S2_59_19  ( .A(\mult_22/ab[59][19] ), .B(
        \mult_22/CARRYB[58][19] ), .CI(\mult_22/SUMB[58][20] ), .CO(
        \mult_22/CARRYB[59][19] ), .S(\mult_22/SUMB[59][19] ) );
  FA_X1 \mult_22/S2_59_18  ( .A(\mult_22/ab[59][18] ), .B(
        \mult_22/CARRYB[58][18] ), .CI(\mult_22/SUMB[58][19] ), .CO(
        \mult_22/CARRYB[59][18] ), .S(\mult_22/SUMB[59][18] ) );
  FA_X1 \mult_22/S2_59_17  ( .A(\mult_22/ab[59][17] ), .B(
        \mult_22/CARRYB[58][17] ), .CI(\mult_22/SUMB[58][18] ), .CO(
        \mult_22/CARRYB[59][17] ), .S(\mult_22/SUMB[59][17] ) );
  FA_X1 \mult_22/S2_59_16  ( .A(\mult_22/ab[59][16] ), .B(
        \mult_22/CARRYB[58][16] ), .CI(\mult_22/SUMB[58][17] ), .CO(
        \mult_22/CARRYB[59][16] ), .S(\mult_22/SUMB[59][16] ) );
  FA_X1 \mult_22/S2_59_15  ( .A(\mult_22/ab[59][15] ), .B(
        \mult_22/CARRYB[58][15] ), .CI(\mult_22/SUMB[58][16] ), .CO(
        \mult_22/CARRYB[59][15] ), .S(\mult_22/SUMB[59][15] ) );
  FA_X1 \mult_22/S2_59_14  ( .A(\mult_22/ab[59][14] ), .B(
        \mult_22/CARRYB[58][14] ), .CI(\mult_22/SUMB[58][15] ), .CO(
        \mult_22/CARRYB[59][14] ), .S(\mult_22/SUMB[59][14] ) );
  FA_X1 \mult_22/S2_59_13  ( .A(\mult_22/ab[59][13] ), .B(
        \mult_22/CARRYB[58][13] ), .CI(\mult_22/SUMB[58][14] ), .CO(
        \mult_22/CARRYB[59][13] ), .S(\mult_22/SUMB[59][13] ) );
  FA_X1 \mult_22/S2_59_12  ( .A(\mult_22/ab[59][12] ), .B(
        \mult_22/CARRYB[58][12] ), .CI(\mult_22/SUMB[58][13] ), .CO(
        \mult_22/CARRYB[59][12] ), .S(\mult_22/SUMB[59][12] ) );
  FA_X1 \mult_22/S2_59_11  ( .A(\mult_22/ab[59][11] ), .B(
        \mult_22/CARRYB[58][11] ), .CI(\mult_22/SUMB[58][12] ), .CO(
        \mult_22/CARRYB[59][11] ), .S(\mult_22/SUMB[59][11] ) );
  FA_X1 \mult_22/S2_59_10  ( .A(\mult_22/ab[59][10] ), .B(
        \mult_22/CARRYB[58][10] ), .CI(\mult_22/SUMB[58][11] ), .CO(
        \mult_22/CARRYB[59][10] ), .S(\mult_22/SUMB[59][10] ) );
  FA_X1 \mult_22/S2_59_9  ( .A(\mult_22/ab[59][9] ), .B(
        \mult_22/CARRYB[58][9] ), .CI(\mult_22/SUMB[58][10] ), .CO(
        \mult_22/CARRYB[59][9] ), .S(\mult_22/SUMB[59][9] ) );
  FA_X1 \mult_22/S2_59_8  ( .A(\mult_22/CARRYB[58][8] ), .B(
        \mult_22/ab[59][8] ), .CI(\mult_22/SUMB[58][9] ), .CO(
        \mult_22/CARRYB[59][8] ), .S(\mult_22/SUMB[59][8] ) );
  FA_X1 \mult_22/S2_59_7  ( .A(\mult_22/CARRYB[58][7] ), .B(
        \mult_22/ab[59][7] ), .CI(\mult_22/SUMB[58][8] ), .CO(
        \mult_22/CARRYB[59][7] ), .S(\mult_22/SUMB[59][7] ) );
  FA_X1 \mult_22/S2_59_6  ( .A(\mult_22/ab[59][6] ), .B(
        \mult_22/CARRYB[58][6] ), .CI(\mult_22/SUMB[58][7] ), .CO(
        \mult_22/CARRYB[59][6] ), .S(\mult_22/SUMB[59][6] ) );
  FA_X1 \mult_22/S2_59_5  ( .A(\mult_22/ab[59][5] ), .B(
        \mult_22/CARRYB[58][5] ), .CI(\mult_22/SUMB[58][6] ), .CO(
        \mult_22/CARRYB[59][5] ), .S(\mult_22/SUMB[59][5] ) );
  FA_X1 \mult_22/S2_59_4  ( .A(\mult_22/ab[59][4] ), .B(
        \mult_22/CARRYB[58][4] ), .CI(\mult_22/SUMB[58][5] ), .CO(
        \mult_22/CARRYB[59][4] ), .S(\mult_22/SUMB[59][4] ) );
  FA_X1 \mult_22/S2_59_3  ( .A(\mult_22/ab[59][3] ), .B(
        \mult_22/CARRYB[58][3] ), .CI(\mult_22/SUMB[58][4] ), .CO(
        \mult_22/CARRYB[59][3] ), .S(\mult_22/SUMB[59][3] ) );
  FA_X1 \mult_22/S2_59_2  ( .A(\mult_22/ab[59][2] ), .B(
        \mult_22/CARRYB[58][2] ), .CI(\mult_22/SUMB[58][3] ), .CO(
        \mult_22/CARRYB[59][2] ), .S(\mult_22/SUMB[59][2] ) );
  FA_X1 \mult_22/S2_59_1  ( .A(\mult_22/ab[59][1] ), .B(
        \mult_22/CARRYB[58][1] ), .CI(\mult_22/SUMB[58][2] ), .CO(
        \mult_22/CARRYB[59][1] ), .S(\mult_22/SUMB[59][1] ) );
  FA_X1 \mult_22/S1_59_0  ( .A(\mult_22/ab[59][0] ), .B(
        \mult_22/CARRYB[58][0] ), .CI(\mult_22/SUMB[58][1] ), .CO(
        \mult_22/CARRYB[59][0] ), .S(N187) );
  FA_X1 \mult_22/S3_60_62  ( .A(\mult_22/ab[60][62] ), .B(
        \mult_22/CARRYB[59][62] ), .CI(\mult_22/ab[59][63] ), .CO(
        \mult_22/CARRYB[60][62] ), .S(\mult_22/SUMB[60][62] ) );
  FA_X1 \mult_22/S2_60_61  ( .A(\mult_22/ab[60][61] ), .B(
        \mult_22/CARRYB[59][61] ), .CI(\mult_22/SUMB[59][62] ), .CO(
        \mult_22/CARRYB[60][61] ), .S(\mult_22/SUMB[60][61] ) );
  FA_X1 \mult_22/S2_60_60  ( .A(\mult_22/ab[60][60] ), .B(
        \mult_22/CARRYB[59][60] ), .CI(\mult_22/SUMB[59][61] ), .CO(
        \mult_22/CARRYB[60][60] ), .S(\mult_22/SUMB[60][60] ) );
  FA_X1 \mult_22/S2_60_59  ( .A(\mult_22/ab[60][59] ), .B(
        \mult_22/CARRYB[59][59] ), .CI(\mult_22/SUMB[59][60] ), .CO(
        \mult_22/CARRYB[60][59] ), .S(\mult_22/SUMB[60][59] ) );
  FA_X1 \mult_22/S2_60_58  ( .A(\mult_22/ab[60][58] ), .B(
        \mult_22/CARRYB[59][58] ), .CI(\mult_22/SUMB[59][59] ), .CO(
        \mult_22/CARRYB[60][58] ), .S(\mult_22/SUMB[60][58] ) );
  FA_X1 \mult_22/S2_60_57  ( .A(\mult_22/ab[60][57] ), .B(
        \mult_22/CARRYB[59][57] ), .CI(\mult_22/SUMB[59][58] ), .CO(
        \mult_22/CARRYB[60][57] ), .S(\mult_22/SUMB[60][57] ) );
  FA_X1 \mult_22/S2_60_56  ( .A(\mult_22/ab[60][56] ), .B(
        \mult_22/CARRYB[59][56] ), .CI(\mult_22/SUMB[59][57] ), .CO(
        \mult_22/CARRYB[60][56] ), .S(\mult_22/SUMB[60][56] ) );
  FA_X1 \mult_22/S2_60_55  ( .A(\mult_22/ab[60][55] ), .B(
        \mult_22/CARRYB[59][55] ), .CI(\mult_22/SUMB[59][56] ), .CO(
        \mult_22/CARRYB[60][55] ), .S(\mult_22/SUMB[60][55] ) );
  FA_X1 \mult_22/S2_60_54  ( .A(\mult_22/ab[60][54] ), .B(
        \mult_22/CARRYB[59][54] ), .CI(\mult_22/SUMB[59][55] ), .CO(
        \mult_22/CARRYB[60][54] ), .S(\mult_22/SUMB[60][54] ) );
  FA_X1 \mult_22/S2_60_53  ( .A(\mult_22/ab[60][53] ), .B(
        \mult_22/CARRYB[59][53] ), .CI(\mult_22/SUMB[59][54] ), .CO(
        \mult_22/CARRYB[60][53] ), .S(\mult_22/SUMB[60][53] ) );
  FA_X1 \mult_22/S2_60_52  ( .A(\mult_22/ab[60][52] ), .B(
        \mult_22/CARRYB[59][52] ), .CI(\mult_22/SUMB[59][53] ), .CO(
        \mult_22/CARRYB[60][52] ), .S(\mult_22/SUMB[60][52] ) );
  FA_X1 \mult_22/S2_60_51  ( .A(\mult_22/ab[60][51] ), .B(
        \mult_22/CARRYB[59][51] ), .CI(\mult_22/SUMB[59][52] ), .CO(
        \mult_22/CARRYB[60][51] ), .S(\mult_22/SUMB[60][51] ) );
  FA_X1 \mult_22/S2_60_50  ( .A(\mult_22/ab[60][50] ), .B(
        \mult_22/CARRYB[59][50] ), .CI(\mult_22/SUMB[59][51] ), .CO(
        \mult_22/CARRYB[60][50] ), .S(\mult_22/SUMB[60][50] ) );
  FA_X1 \mult_22/S2_60_49  ( .A(\mult_22/ab[60][49] ), .B(
        \mult_22/CARRYB[59][49] ), .CI(\mult_22/SUMB[59][50] ), .CO(
        \mult_22/CARRYB[60][49] ), .S(\mult_22/SUMB[60][49] ) );
  FA_X1 \mult_22/S2_60_48  ( .A(\mult_22/ab[60][48] ), .B(
        \mult_22/CARRYB[59][48] ), .CI(\mult_22/SUMB[59][49] ), .CO(
        \mult_22/CARRYB[60][48] ), .S(\mult_22/SUMB[60][48] ) );
  FA_X1 \mult_22/S2_60_47  ( .A(\mult_22/ab[60][47] ), .B(
        \mult_22/CARRYB[59][47] ), .CI(\mult_22/SUMB[59][48] ), .CO(
        \mult_22/CARRYB[60][47] ), .S(\mult_22/SUMB[60][47] ) );
  FA_X1 \mult_22/S2_60_46  ( .A(\mult_22/ab[60][46] ), .B(
        \mult_22/CARRYB[59][46] ), .CI(\mult_22/SUMB[59][47] ), .CO(
        \mult_22/CARRYB[60][46] ), .S(\mult_22/SUMB[60][46] ) );
  FA_X1 \mult_22/S2_60_45  ( .A(\mult_22/ab[60][45] ), .B(
        \mult_22/CARRYB[59][45] ), .CI(\mult_22/SUMB[59][46] ), .CO(
        \mult_22/CARRYB[60][45] ), .S(\mult_22/SUMB[60][45] ) );
  FA_X1 \mult_22/S2_60_44  ( .A(\mult_22/ab[60][44] ), .B(
        \mult_22/CARRYB[59][44] ), .CI(\mult_22/SUMB[59][45] ), .CO(
        \mult_22/CARRYB[60][44] ), .S(\mult_22/SUMB[60][44] ) );
  FA_X1 \mult_22/S2_60_43  ( .A(\mult_22/ab[60][43] ), .B(
        \mult_22/CARRYB[59][43] ), .CI(\mult_22/SUMB[59][44] ), .CO(
        \mult_22/CARRYB[60][43] ), .S(\mult_22/SUMB[60][43] ) );
  FA_X1 \mult_22/S2_60_42  ( .A(\mult_22/ab[60][42] ), .B(
        \mult_22/CARRYB[59][42] ), .CI(\mult_22/SUMB[59][43] ), .CO(
        \mult_22/CARRYB[60][42] ), .S(\mult_22/SUMB[60][42] ) );
  FA_X1 \mult_22/S2_60_41  ( .A(\mult_22/ab[60][41] ), .B(
        \mult_22/CARRYB[59][41] ), .CI(\mult_22/SUMB[59][42] ), .CO(
        \mult_22/CARRYB[60][41] ), .S(\mult_22/SUMB[60][41] ) );
  FA_X1 \mult_22/S2_60_40  ( .A(\mult_22/ab[60][40] ), .B(
        \mult_22/CARRYB[59][40] ), .CI(\mult_22/SUMB[59][41] ), .CO(
        \mult_22/CARRYB[60][40] ), .S(\mult_22/SUMB[60][40] ) );
  FA_X1 \mult_22/S2_60_39  ( .A(\mult_22/ab[60][39] ), .B(
        \mult_22/CARRYB[59][39] ), .CI(\mult_22/SUMB[59][40] ), .CO(
        \mult_22/CARRYB[60][39] ), .S(\mult_22/SUMB[60][39] ) );
  FA_X1 \mult_22/S2_60_38  ( .A(\mult_22/ab[60][38] ), .B(
        \mult_22/CARRYB[59][38] ), .CI(\mult_22/SUMB[59][39] ), .CO(
        \mult_22/CARRYB[60][38] ), .S(\mult_22/SUMB[60][38] ) );
  FA_X1 \mult_22/S2_60_37  ( .A(\mult_22/ab[60][37] ), .B(
        \mult_22/CARRYB[59][37] ), .CI(\mult_22/SUMB[59][38] ), .CO(
        \mult_22/CARRYB[60][37] ), .S(\mult_22/SUMB[60][37] ) );
  FA_X1 \mult_22/S2_60_36  ( .A(\mult_22/ab[60][36] ), .B(
        \mult_22/CARRYB[59][36] ), .CI(\mult_22/SUMB[59][37] ), .CO(
        \mult_22/CARRYB[60][36] ), .S(\mult_22/SUMB[60][36] ) );
  FA_X1 \mult_22/S2_60_35  ( .A(\mult_22/ab[60][35] ), .B(
        \mult_22/CARRYB[59][35] ), .CI(\mult_22/SUMB[59][36] ), .CO(
        \mult_22/CARRYB[60][35] ), .S(\mult_22/SUMB[60][35] ) );
  FA_X1 \mult_22/S2_60_34  ( .A(\mult_22/ab[60][34] ), .B(
        \mult_22/CARRYB[59][34] ), .CI(\mult_22/SUMB[59][35] ), .CO(
        \mult_22/CARRYB[60][34] ), .S(\mult_22/SUMB[60][34] ) );
  FA_X1 \mult_22/S2_60_33  ( .A(\mult_22/ab[60][33] ), .B(
        \mult_22/CARRYB[59][33] ), .CI(\mult_22/SUMB[59][34] ), .CO(
        \mult_22/CARRYB[60][33] ), .S(\mult_22/SUMB[60][33] ) );
  FA_X1 \mult_22/S2_60_32  ( .A(\mult_22/ab[60][32] ), .B(
        \mult_22/CARRYB[59][32] ), .CI(\mult_22/SUMB[59][33] ), .CO(
        \mult_22/CARRYB[60][32] ), .S(\mult_22/SUMB[60][32] ) );
  FA_X1 \mult_22/S2_60_31  ( .A(\mult_22/ab[60][31] ), .B(
        \mult_22/CARRYB[59][31] ), .CI(\mult_22/SUMB[59][32] ), .CO(
        \mult_22/CARRYB[60][31] ), .S(\mult_22/SUMB[60][31] ) );
  FA_X1 \mult_22/S2_60_30  ( .A(\mult_22/ab[60][30] ), .B(
        \mult_22/CARRYB[59][30] ), .CI(\mult_22/SUMB[59][31] ), .CO(
        \mult_22/CARRYB[60][30] ), .S(\mult_22/SUMB[60][30] ) );
  FA_X1 \mult_22/S2_60_29  ( .A(\mult_22/ab[60][29] ), .B(
        \mult_22/CARRYB[59][29] ), .CI(\mult_22/SUMB[59][30] ), .CO(
        \mult_22/CARRYB[60][29] ), .S(\mult_22/SUMB[60][29] ) );
  FA_X1 \mult_22/S2_60_28  ( .A(\mult_22/ab[60][28] ), .B(
        \mult_22/CARRYB[59][28] ), .CI(\mult_22/SUMB[59][29] ), .CO(
        \mult_22/CARRYB[60][28] ), .S(\mult_22/SUMB[60][28] ) );
  FA_X1 \mult_22/S2_60_27  ( .A(\mult_22/ab[60][27] ), .B(
        \mult_22/CARRYB[59][27] ), .CI(\mult_22/SUMB[59][28] ), .CO(
        \mult_22/CARRYB[60][27] ), .S(\mult_22/SUMB[60][27] ) );
  FA_X1 \mult_22/S2_60_26  ( .A(\mult_22/ab[60][26] ), .B(
        \mult_22/CARRYB[59][26] ), .CI(\mult_22/SUMB[59][27] ), .CO(
        \mult_22/CARRYB[60][26] ), .S(\mult_22/SUMB[60][26] ) );
  FA_X1 \mult_22/S2_60_25  ( .A(\mult_22/ab[60][25] ), .B(
        \mult_22/CARRYB[59][25] ), .CI(\mult_22/SUMB[59][26] ), .CO(
        \mult_22/CARRYB[60][25] ), .S(\mult_22/SUMB[60][25] ) );
  FA_X1 \mult_22/S2_60_24  ( .A(\mult_22/ab[60][24] ), .B(
        \mult_22/CARRYB[59][24] ), .CI(\mult_22/SUMB[59][25] ), .CO(
        \mult_22/CARRYB[60][24] ), .S(\mult_22/SUMB[60][24] ) );
  FA_X1 \mult_22/S2_60_23  ( .A(\mult_22/ab[60][23] ), .B(
        \mult_22/CARRYB[59][23] ), .CI(\mult_22/SUMB[59][24] ), .CO(
        \mult_22/CARRYB[60][23] ), .S(\mult_22/SUMB[60][23] ) );
  FA_X1 \mult_22/S2_60_22  ( .A(\mult_22/ab[60][22] ), .B(
        \mult_22/CARRYB[59][22] ), .CI(\mult_22/SUMB[59][23] ), .CO(
        \mult_22/CARRYB[60][22] ), .S(\mult_22/SUMB[60][22] ) );
  FA_X1 \mult_22/S2_60_21  ( .A(\mult_22/ab[60][21] ), .B(
        \mult_22/CARRYB[59][21] ), .CI(\mult_22/SUMB[59][22] ), .CO(
        \mult_22/CARRYB[60][21] ), .S(\mult_22/SUMB[60][21] ) );
  FA_X1 \mult_22/S2_60_20  ( .A(\mult_22/ab[60][20] ), .B(
        \mult_22/CARRYB[59][20] ), .CI(\mult_22/SUMB[59][21] ), .CO(
        \mult_22/CARRYB[60][20] ), .S(\mult_22/SUMB[60][20] ) );
  FA_X1 \mult_22/S2_60_19  ( .A(\mult_22/ab[60][19] ), .B(
        \mult_22/CARRYB[59][19] ), .CI(\mult_22/SUMB[59][20] ), .CO(
        \mult_22/CARRYB[60][19] ), .S(\mult_22/SUMB[60][19] ) );
  FA_X1 \mult_22/S2_60_18  ( .A(\mult_22/ab[60][18] ), .B(
        \mult_22/CARRYB[59][18] ), .CI(\mult_22/SUMB[59][19] ), .CO(
        \mult_22/CARRYB[60][18] ), .S(\mult_22/SUMB[60][18] ) );
  FA_X1 \mult_22/S2_60_17  ( .A(\mult_22/ab[60][17] ), .B(
        \mult_22/CARRYB[59][17] ), .CI(\mult_22/SUMB[59][18] ), .CO(
        \mult_22/CARRYB[60][17] ), .S(\mult_22/SUMB[60][17] ) );
  FA_X1 \mult_22/S2_60_16  ( .A(\mult_22/ab[60][16] ), .B(
        \mult_22/CARRYB[59][16] ), .CI(\mult_22/SUMB[59][17] ), .CO(
        \mult_22/CARRYB[60][16] ), .S(\mult_22/SUMB[60][16] ) );
  FA_X1 \mult_22/S2_60_15  ( .A(\mult_22/ab[60][15] ), .B(
        \mult_22/CARRYB[59][15] ), .CI(\mult_22/SUMB[59][16] ), .CO(
        \mult_22/CARRYB[60][15] ), .S(\mult_22/SUMB[60][15] ) );
  FA_X1 \mult_22/S2_60_14  ( .A(\mult_22/ab[60][14] ), .B(
        \mult_22/CARRYB[59][14] ), .CI(\mult_22/SUMB[59][15] ), .CO(
        \mult_22/CARRYB[60][14] ), .S(\mult_22/SUMB[60][14] ) );
  FA_X1 \mult_22/S2_60_13  ( .A(\mult_22/ab[60][13] ), .B(
        \mult_22/CARRYB[59][13] ), .CI(\mult_22/SUMB[59][14] ), .CO(
        \mult_22/CARRYB[60][13] ), .S(\mult_22/SUMB[60][13] ) );
  FA_X1 \mult_22/S2_60_12  ( .A(\mult_22/ab[60][12] ), .B(
        \mult_22/CARRYB[59][12] ), .CI(\mult_22/SUMB[59][13] ), .CO(
        \mult_22/CARRYB[60][12] ), .S(\mult_22/SUMB[60][12] ) );
  FA_X1 \mult_22/S2_60_11  ( .A(\mult_22/ab[60][11] ), .B(
        \mult_22/CARRYB[59][11] ), .CI(\mult_22/SUMB[59][12] ), .CO(
        \mult_22/CARRYB[60][11] ), .S(\mult_22/SUMB[60][11] ) );
  FA_X1 \mult_22/S2_60_10  ( .A(\mult_22/ab[60][10] ), .B(
        \mult_22/CARRYB[59][10] ), .CI(\mult_22/SUMB[59][11] ), .CO(
        \mult_22/CARRYB[60][10] ), .S(\mult_22/SUMB[60][10] ) );
  FA_X1 \mult_22/S2_60_9  ( .A(\mult_22/ab[60][9] ), .B(
        \mult_22/CARRYB[59][9] ), .CI(\mult_22/SUMB[59][10] ), .CO(
        \mult_22/CARRYB[60][9] ), .S(\mult_22/SUMB[60][9] ) );
  FA_X1 \mult_22/S2_60_8  ( .A(\mult_22/ab[60][8] ), .B(
        \mult_22/CARRYB[59][8] ), .CI(\mult_22/SUMB[59][9] ), .CO(
        \mult_22/CARRYB[60][8] ), .S(\mult_22/SUMB[60][8] ) );
  FA_X1 \mult_22/S2_60_7  ( .A(\mult_22/ab[60][7] ), .B(
        \mult_22/CARRYB[59][7] ), .CI(\mult_22/SUMB[59][8] ), .CO(
        \mult_22/CARRYB[60][7] ), .S(\mult_22/SUMB[60][7] ) );
  FA_X1 \mult_22/S2_60_6  ( .A(\mult_22/CARRYB[59][6] ), .B(
        \mult_22/ab[60][6] ), .CI(\mult_22/SUMB[59][7] ), .CO(
        \mult_22/CARRYB[60][6] ), .S(\mult_22/SUMB[60][6] ) );
  FA_X1 \mult_22/S2_60_5  ( .A(\mult_22/CARRYB[59][5] ), .B(
        \mult_22/ab[60][5] ), .CI(\mult_22/SUMB[59][6] ), .CO(
        \mult_22/CARRYB[60][5] ), .S(\mult_22/SUMB[60][5] ) );
  FA_X1 \mult_22/S2_60_4  ( .A(\mult_22/ab[60][4] ), .B(
        \mult_22/CARRYB[59][4] ), .CI(\mult_22/SUMB[59][5] ), .CO(
        \mult_22/CARRYB[60][4] ), .S(\mult_22/SUMB[60][4] ) );
  FA_X1 \mult_22/S2_60_3  ( .A(\mult_22/ab[60][3] ), .B(
        \mult_22/CARRYB[59][3] ), .CI(\mult_22/SUMB[59][4] ), .CO(
        \mult_22/CARRYB[60][3] ), .S(\mult_22/SUMB[60][3] ) );
  FA_X1 \mult_22/S2_60_2  ( .A(\mult_22/ab[60][2] ), .B(
        \mult_22/CARRYB[59][2] ), .CI(\mult_22/SUMB[59][3] ), .CO(
        \mult_22/CARRYB[60][2] ), .S(\mult_22/SUMB[60][2] ) );
  FA_X1 \mult_22/S2_60_1  ( .A(\mult_22/ab[60][1] ), .B(
        \mult_22/CARRYB[59][1] ), .CI(\mult_22/SUMB[59][2] ), .CO(
        \mult_22/CARRYB[60][1] ), .S(\mult_22/SUMB[60][1] ) );
  FA_X1 \mult_22/S1_60_0  ( .A(\mult_22/ab[60][0] ), .B(
        \mult_22/CARRYB[59][0] ), .CI(\mult_22/SUMB[59][1] ), .CO(
        \mult_22/CARRYB[60][0] ), .S(N188) );
  FA_X1 \mult_22/S3_61_62  ( .A(\mult_22/ab[61][62] ), .B(
        \mult_22/CARRYB[60][62] ), .CI(\mult_22/ab[60][63] ), .CO(
        \mult_22/CARRYB[61][62] ), .S(\mult_22/SUMB[61][62] ) );
  FA_X1 \mult_22/S2_61_61  ( .A(\mult_22/ab[61][61] ), .B(
        \mult_22/CARRYB[60][61] ), .CI(\mult_22/SUMB[60][62] ), .CO(
        \mult_22/CARRYB[61][61] ), .S(\mult_22/SUMB[61][61] ) );
  FA_X1 \mult_22/S2_61_60  ( .A(\mult_22/ab[61][60] ), .B(
        \mult_22/CARRYB[60][60] ), .CI(\mult_22/SUMB[60][61] ), .CO(
        \mult_22/CARRYB[61][60] ), .S(\mult_22/SUMB[61][60] ) );
  FA_X1 \mult_22/S2_61_59  ( .A(\mult_22/ab[61][59] ), .B(
        \mult_22/CARRYB[60][59] ), .CI(\mult_22/SUMB[60][60] ), .CO(
        \mult_22/CARRYB[61][59] ), .S(\mult_22/SUMB[61][59] ) );
  FA_X1 \mult_22/S2_61_58  ( .A(\mult_22/ab[61][58] ), .B(
        \mult_22/CARRYB[60][58] ), .CI(\mult_22/SUMB[60][59] ), .CO(
        \mult_22/CARRYB[61][58] ), .S(\mult_22/SUMB[61][58] ) );
  FA_X1 \mult_22/S2_61_57  ( .A(\mult_22/ab[61][57] ), .B(
        \mult_22/CARRYB[60][57] ), .CI(\mult_22/SUMB[60][58] ), .CO(
        \mult_22/CARRYB[61][57] ), .S(\mult_22/SUMB[61][57] ) );
  FA_X1 \mult_22/S2_61_56  ( .A(\mult_22/ab[61][56] ), .B(
        \mult_22/CARRYB[60][56] ), .CI(\mult_22/SUMB[60][57] ), .CO(
        \mult_22/CARRYB[61][56] ), .S(\mult_22/SUMB[61][56] ) );
  FA_X1 \mult_22/S2_61_55  ( .A(\mult_22/ab[61][55] ), .B(
        \mult_22/CARRYB[60][55] ), .CI(\mult_22/SUMB[60][56] ), .CO(
        \mult_22/CARRYB[61][55] ), .S(\mult_22/SUMB[61][55] ) );
  FA_X1 \mult_22/S2_61_54  ( .A(\mult_22/ab[61][54] ), .B(
        \mult_22/CARRYB[60][54] ), .CI(\mult_22/SUMB[60][55] ), .CO(
        \mult_22/CARRYB[61][54] ), .S(\mult_22/SUMB[61][54] ) );
  FA_X1 \mult_22/S2_61_53  ( .A(\mult_22/ab[61][53] ), .B(
        \mult_22/CARRYB[60][53] ), .CI(\mult_22/SUMB[60][54] ), .CO(
        \mult_22/CARRYB[61][53] ), .S(\mult_22/SUMB[61][53] ) );
  FA_X1 \mult_22/S2_61_52  ( .A(\mult_22/ab[61][52] ), .B(
        \mult_22/CARRYB[60][52] ), .CI(\mult_22/SUMB[60][53] ), .CO(
        \mult_22/CARRYB[61][52] ), .S(\mult_22/SUMB[61][52] ) );
  FA_X1 \mult_22/S2_61_51  ( .A(\mult_22/ab[61][51] ), .B(
        \mult_22/CARRYB[60][51] ), .CI(\mult_22/SUMB[60][52] ), .CO(
        \mult_22/CARRYB[61][51] ), .S(\mult_22/SUMB[61][51] ) );
  FA_X1 \mult_22/S2_61_50  ( .A(\mult_22/ab[61][50] ), .B(
        \mult_22/CARRYB[60][50] ), .CI(\mult_22/SUMB[60][51] ), .CO(
        \mult_22/CARRYB[61][50] ), .S(\mult_22/SUMB[61][50] ) );
  FA_X1 \mult_22/S2_61_49  ( .A(\mult_22/ab[61][49] ), .B(
        \mult_22/CARRYB[60][49] ), .CI(\mult_22/SUMB[60][50] ), .CO(
        \mult_22/CARRYB[61][49] ), .S(\mult_22/SUMB[61][49] ) );
  FA_X1 \mult_22/S2_61_48  ( .A(\mult_22/ab[61][48] ), .B(
        \mult_22/CARRYB[60][48] ), .CI(\mult_22/SUMB[60][49] ), .CO(
        \mult_22/CARRYB[61][48] ), .S(\mult_22/SUMB[61][48] ) );
  FA_X1 \mult_22/S2_61_47  ( .A(\mult_22/ab[61][47] ), .B(
        \mult_22/CARRYB[60][47] ), .CI(\mult_22/SUMB[60][48] ), .CO(
        \mult_22/CARRYB[61][47] ), .S(\mult_22/SUMB[61][47] ) );
  FA_X1 \mult_22/S2_61_46  ( .A(\mult_22/ab[61][46] ), .B(
        \mult_22/CARRYB[60][46] ), .CI(\mult_22/SUMB[60][47] ), .CO(
        \mult_22/CARRYB[61][46] ), .S(\mult_22/SUMB[61][46] ) );
  FA_X1 \mult_22/S2_61_45  ( .A(\mult_22/ab[61][45] ), .B(
        \mult_22/CARRYB[60][45] ), .CI(\mult_22/SUMB[60][46] ), .CO(
        \mult_22/CARRYB[61][45] ), .S(\mult_22/SUMB[61][45] ) );
  FA_X1 \mult_22/S2_61_44  ( .A(\mult_22/ab[61][44] ), .B(
        \mult_22/CARRYB[60][44] ), .CI(\mult_22/SUMB[60][45] ), .CO(
        \mult_22/CARRYB[61][44] ), .S(\mult_22/SUMB[61][44] ) );
  FA_X1 \mult_22/S2_61_43  ( .A(\mult_22/ab[61][43] ), .B(
        \mult_22/CARRYB[60][43] ), .CI(\mult_22/SUMB[60][44] ), .CO(
        \mult_22/CARRYB[61][43] ), .S(\mult_22/SUMB[61][43] ) );
  FA_X1 \mult_22/S2_61_42  ( .A(\mult_22/ab[61][42] ), .B(
        \mult_22/CARRYB[60][42] ), .CI(\mult_22/SUMB[60][43] ), .CO(
        \mult_22/CARRYB[61][42] ), .S(\mult_22/SUMB[61][42] ) );
  FA_X1 \mult_22/S2_61_41  ( .A(\mult_22/ab[61][41] ), .B(
        \mult_22/CARRYB[60][41] ), .CI(\mult_22/SUMB[60][42] ), .CO(
        \mult_22/CARRYB[61][41] ), .S(\mult_22/SUMB[61][41] ) );
  FA_X1 \mult_22/S2_61_40  ( .A(\mult_22/ab[61][40] ), .B(
        \mult_22/CARRYB[60][40] ), .CI(\mult_22/SUMB[60][41] ), .CO(
        \mult_22/CARRYB[61][40] ), .S(\mult_22/SUMB[61][40] ) );
  FA_X1 \mult_22/S2_61_39  ( .A(\mult_22/ab[61][39] ), .B(
        \mult_22/CARRYB[60][39] ), .CI(\mult_22/SUMB[60][40] ), .CO(
        \mult_22/CARRYB[61][39] ), .S(\mult_22/SUMB[61][39] ) );
  FA_X1 \mult_22/S2_61_38  ( .A(\mult_22/ab[61][38] ), .B(
        \mult_22/CARRYB[60][38] ), .CI(\mult_22/SUMB[60][39] ), .CO(
        \mult_22/CARRYB[61][38] ), .S(\mult_22/SUMB[61][38] ) );
  FA_X1 \mult_22/S2_61_37  ( .A(\mult_22/ab[61][37] ), .B(
        \mult_22/CARRYB[60][37] ), .CI(\mult_22/SUMB[60][38] ), .CO(
        \mult_22/CARRYB[61][37] ), .S(\mult_22/SUMB[61][37] ) );
  FA_X1 \mult_22/S2_61_36  ( .A(\mult_22/ab[61][36] ), .B(
        \mult_22/CARRYB[60][36] ), .CI(\mult_22/SUMB[60][37] ), .CO(
        \mult_22/CARRYB[61][36] ), .S(\mult_22/SUMB[61][36] ) );
  FA_X1 \mult_22/S2_61_35  ( .A(\mult_22/ab[61][35] ), .B(
        \mult_22/CARRYB[60][35] ), .CI(\mult_22/SUMB[60][36] ), .CO(
        \mult_22/CARRYB[61][35] ), .S(\mult_22/SUMB[61][35] ) );
  FA_X1 \mult_22/S2_61_34  ( .A(\mult_22/ab[61][34] ), .B(
        \mult_22/CARRYB[60][34] ), .CI(\mult_22/SUMB[60][35] ), .CO(
        \mult_22/CARRYB[61][34] ), .S(\mult_22/SUMB[61][34] ) );
  FA_X1 \mult_22/S2_61_33  ( .A(\mult_22/ab[61][33] ), .B(
        \mult_22/CARRYB[60][33] ), .CI(\mult_22/SUMB[60][34] ), .CO(
        \mult_22/CARRYB[61][33] ), .S(\mult_22/SUMB[61][33] ) );
  FA_X1 \mult_22/S2_61_32  ( .A(\mult_22/ab[61][32] ), .B(
        \mult_22/CARRYB[60][32] ), .CI(\mult_22/SUMB[60][33] ), .CO(
        \mult_22/CARRYB[61][32] ), .S(\mult_22/SUMB[61][32] ) );
  FA_X1 \mult_22/S2_61_31  ( .A(\mult_22/ab[61][31] ), .B(
        \mult_22/CARRYB[60][31] ), .CI(\mult_22/SUMB[60][32] ), .CO(
        \mult_22/CARRYB[61][31] ), .S(\mult_22/SUMB[61][31] ) );
  FA_X1 \mult_22/S2_61_30  ( .A(\mult_22/ab[61][30] ), .B(
        \mult_22/CARRYB[60][30] ), .CI(\mult_22/SUMB[60][31] ), .CO(
        \mult_22/CARRYB[61][30] ), .S(\mult_22/SUMB[61][30] ) );
  FA_X1 \mult_22/S2_61_29  ( .A(\mult_22/ab[61][29] ), .B(
        \mult_22/CARRYB[60][29] ), .CI(\mult_22/SUMB[60][30] ), .CO(
        \mult_22/CARRYB[61][29] ), .S(\mult_22/SUMB[61][29] ) );
  FA_X1 \mult_22/S2_61_28  ( .A(\mult_22/ab[61][28] ), .B(
        \mult_22/CARRYB[60][28] ), .CI(\mult_22/SUMB[60][29] ), .CO(
        \mult_22/CARRYB[61][28] ), .S(\mult_22/SUMB[61][28] ) );
  FA_X1 \mult_22/S2_61_27  ( .A(\mult_22/ab[61][27] ), .B(
        \mult_22/CARRYB[60][27] ), .CI(\mult_22/SUMB[60][28] ), .CO(
        \mult_22/CARRYB[61][27] ), .S(\mult_22/SUMB[61][27] ) );
  FA_X1 \mult_22/S2_61_26  ( .A(\mult_22/ab[61][26] ), .B(
        \mult_22/CARRYB[60][26] ), .CI(\mult_22/SUMB[60][27] ), .CO(
        \mult_22/CARRYB[61][26] ), .S(\mult_22/SUMB[61][26] ) );
  FA_X1 \mult_22/S2_61_25  ( .A(\mult_22/ab[61][25] ), .B(
        \mult_22/CARRYB[60][25] ), .CI(\mult_22/SUMB[60][26] ), .CO(
        \mult_22/CARRYB[61][25] ), .S(\mult_22/SUMB[61][25] ) );
  FA_X1 \mult_22/S2_61_24  ( .A(\mult_22/ab[61][24] ), .B(
        \mult_22/CARRYB[60][24] ), .CI(\mult_22/SUMB[60][25] ), .CO(
        \mult_22/CARRYB[61][24] ), .S(\mult_22/SUMB[61][24] ) );
  FA_X1 \mult_22/S2_61_23  ( .A(\mult_22/ab[61][23] ), .B(
        \mult_22/CARRYB[60][23] ), .CI(\mult_22/SUMB[60][24] ), .CO(
        \mult_22/CARRYB[61][23] ), .S(\mult_22/SUMB[61][23] ) );
  FA_X1 \mult_22/S2_61_22  ( .A(\mult_22/ab[61][22] ), .B(
        \mult_22/CARRYB[60][22] ), .CI(\mult_22/SUMB[60][23] ), .CO(
        \mult_22/CARRYB[61][22] ), .S(\mult_22/SUMB[61][22] ) );
  FA_X1 \mult_22/S2_61_21  ( .A(\mult_22/ab[61][21] ), .B(
        \mult_22/CARRYB[60][21] ), .CI(\mult_22/SUMB[60][22] ), .CO(
        \mult_22/CARRYB[61][21] ), .S(\mult_22/SUMB[61][21] ) );
  FA_X1 \mult_22/S2_61_20  ( .A(\mult_22/ab[61][20] ), .B(
        \mult_22/CARRYB[60][20] ), .CI(\mult_22/SUMB[60][21] ), .CO(
        \mult_22/CARRYB[61][20] ), .S(\mult_22/SUMB[61][20] ) );
  FA_X1 \mult_22/S2_61_19  ( .A(\mult_22/ab[61][19] ), .B(
        \mult_22/CARRYB[60][19] ), .CI(\mult_22/SUMB[60][20] ), .CO(
        \mult_22/CARRYB[61][19] ), .S(\mult_22/SUMB[61][19] ) );
  FA_X1 \mult_22/S2_61_18  ( .A(\mult_22/ab[61][18] ), .B(
        \mult_22/CARRYB[60][18] ), .CI(\mult_22/SUMB[60][19] ), .CO(
        \mult_22/CARRYB[61][18] ), .S(\mult_22/SUMB[61][18] ) );
  FA_X1 \mult_22/S2_61_17  ( .A(\mult_22/ab[61][17] ), .B(
        \mult_22/CARRYB[60][17] ), .CI(\mult_22/SUMB[60][18] ), .CO(
        \mult_22/CARRYB[61][17] ), .S(\mult_22/SUMB[61][17] ) );
  FA_X1 \mult_22/S2_61_16  ( .A(\mult_22/ab[61][16] ), .B(
        \mult_22/CARRYB[60][16] ), .CI(\mult_22/SUMB[60][17] ), .CO(
        \mult_22/CARRYB[61][16] ), .S(\mult_22/SUMB[61][16] ) );
  FA_X1 \mult_22/S2_61_15  ( .A(\mult_22/ab[61][15] ), .B(
        \mult_22/CARRYB[60][15] ), .CI(\mult_22/SUMB[60][16] ), .CO(
        \mult_22/CARRYB[61][15] ), .S(\mult_22/SUMB[61][15] ) );
  FA_X1 \mult_22/S2_61_14  ( .A(\mult_22/ab[61][14] ), .B(
        \mult_22/CARRYB[60][14] ), .CI(\mult_22/SUMB[60][15] ), .CO(
        \mult_22/CARRYB[61][14] ), .S(\mult_22/SUMB[61][14] ) );
  FA_X1 \mult_22/S2_61_13  ( .A(\mult_22/ab[61][13] ), .B(
        \mult_22/CARRYB[60][13] ), .CI(\mult_22/SUMB[60][14] ), .CO(
        \mult_22/CARRYB[61][13] ), .S(\mult_22/SUMB[61][13] ) );
  FA_X1 \mult_22/S2_61_12  ( .A(\mult_22/ab[61][12] ), .B(
        \mult_22/CARRYB[60][12] ), .CI(\mult_22/SUMB[60][13] ), .CO(
        \mult_22/CARRYB[61][12] ), .S(\mult_22/SUMB[61][12] ) );
  FA_X1 \mult_22/S2_61_11  ( .A(\mult_22/ab[61][11] ), .B(
        \mult_22/CARRYB[60][11] ), .CI(\mult_22/SUMB[60][12] ), .CO(
        \mult_22/CARRYB[61][11] ), .S(\mult_22/SUMB[61][11] ) );
  FA_X1 \mult_22/S2_61_10  ( .A(\mult_22/ab[61][10] ), .B(
        \mult_22/CARRYB[60][10] ), .CI(\mult_22/SUMB[60][11] ), .CO(
        \mult_22/CARRYB[61][10] ), .S(\mult_22/SUMB[61][10] ) );
  FA_X1 \mult_22/S2_61_9  ( .A(\mult_22/ab[61][9] ), .B(
        \mult_22/CARRYB[60][9] ), .CI(\mult_22/SUMB[60][10] ), .CO(
        \mult_22/CARRYB[61][9] ), .S(\mult_22/SUMB[61][9] ) );
  FA_X1 \mult_22/S2_61_8  ( .A(\mult_22/ab[61][8] ), .B(
        \mult_22/CARRYB[60][8] ), .CI(\mult_22/SUMB[60][9] ), .CO(
        \mult_22/CARRYB[61][8] ), .S(\mult_22/SUMB[61][8] ) );
  FA_X1 \mult_22/S2_61_7  ( .A(\mult_22/ab[61][7] ), .B(
        \mult_22/CARRYB[60][7] ), .CI(\mult_22/SUMB[60][8] ), .CO(
        \mult_22/CARRYB[61][7] ), .S(\mult_22/SUMB[61][7] ) );
  FA_X1 \mult_22/S2_61_6  ( .A(\mult_22/CARRYB[60][6] ), .B(
        \mult_22/ab[61][6] ), .CI(\mult_22/SUMB[60][7] ), .CO(
        \mult_22/CARRYB[61][6] ), .S(\mult_22/SUMB[61][6] ) );
  FA_X1 \mult_22/S2_61_5  ( .A(\mult_22/CARRYB[60][5] ), .B(
        \mult_22/ab[61][5] ), .CI(\mult_22/SUMB[60][6] ), .CO(
        \mult_22/CARRYB[61][5] ), .S(\mult_22/SUMB[61][5] ) );
  FA_X1 \mult_22/S2_61_4  ( .A(\mult_22/ab[61][4] ), .B(
        \mult_22/CARRYB[60][4] ), .CI(\mult_22/SUMB[60][5] ), .CO(
        \mult_22/CARRYB[61][4] ), .S(\mult_22/SUMB[61][4] ) );
  FA_X1 \mult_22/S2_61_3  ( .A(\mult_22/ab[61][3] ), .B(
        \mult_22/CARRYB[60][3] ), .CI(\mult_22/SUMB[60][4] ), .CO(
        \mult_22/CARRYB[61][3] ), .S(\mult_22/SUMB[61][3] ) );
  FA_X1 \mult_22/S2_61_2  ( .A(\mult_22/ab[61][2] ), .B(
        \mult_22/CARRYB[60][2] ), .CI(\mult_22/SUMB[60][3] ), .CO(
        \mult_22/CARRYB[61][2] ), .S(\mult_22/SUMB[61][2] ) );
  FA_X1 \mult_22/S2_61_1  ( .A(\mult_22/ab[61][1] ), .B(
        \mult_22/CARRYB[60][1] ), .CI(\mult_22/SUMB[60][2] ), .CO(
        \mult_22/CARRYB[61][1] ), .S(\mult_22/SUMB[61][1] ) );
  FA_X1 \mult_22/S1_61_0  ( .A(\mult_22/ab[61][0] ), .B(
        \mult_22/CARRYB[60][0] ), .CI(\mult_22/SUMB[60][1] ), .CO(
        \mult_22/CARRYB[61][0] ), .S(N189) );
  FA_X1 \mult_22/S3_62_62  ( .A(\mult_22/ab[62][62] ), .B(
        \mult_22/CARRYB[61][62] ), .CI(\mult_22/ab[61][63] ), .CO(
        \mult_22/CARRYB[62][62] ), .S(\mult_22/SUMB[62][62] ) );
  FA_X1 \mult_22/S2_62_61  ( .A(\mult_22/ab[62][61] ), .B(
        \mult_22/CARRYB[61][61] ), .CI(\mult_22/SUMB[61][62] ), .CO(
        \mult_22/CARRYB[62][61] ), .S(\mult_22/SUMB[62][61] ) );
  FA_X1 \mult_22/S2_62_60  ( .A(\mult_22/ab[62][60] ), .B(
        \mult_22/CARRYB[61][60] ), .CI(\mult_22/SUMB[61][61] ), .CO(
        \mult_22/CARRYB[62][60] ), .S(\mult_22/SUMB[62][60] ) );
  FA_X1 \mult_22/S2_62_59  ( .A(\mult_22/ab[62][59] ), .B(
        \mult_22/CARRYB[61][59] ), .CI(\mult_22/SUMB[61][60] ), .CO(
        \mult_22/CARRYB[62][59] ), .S(\mult_22/SUMB[62][59] ) );
  FA_X1 \mult_22/S2_62_58  ( .A(\mult_22/ab[62][58] ), .B(
        \mult_22/CARRYB[61][58] ), .CI(\mult_22/SUMB[61][59] ), .CO(
        \mult_22/CARRYB[62][58] ), .S(\mult_22/SUMB[62][58] ) );
  FA_X1 \mult_22/S2_62_57  ( .A(\mult_22/ab[62][57] ), .B(
        \mult_22/CARRYB[61][57] ), .CI(\mult_22/SUMB[61][58] ), .CO(
        \mult_22/CARRYB[62][57] ), .S(\mult_22/SUMB[62][57] ) );
  FA_X1 \mult_22/S2_62_56  ( .A(\mult_22/ab[62][56] ), .B(
        \mult_22/CARRYB[61][56] ), .CI(\mult_22/SUMB[61][57] ), .CO(
        \mult_22/CARRYB[62][56] ), .S(\mult_22/SUMB[62][56] ) );
  FA_X1 \mult_22/S2_62_55  ( .A(\mult_22/ab[62][55] ), .B(
        \mult_22/CARRYB[61][55] ), .CI(\mult_22/SUMB[61][56] ), .CO(
        \mult_22/CARRYB[62][55] ), .S(\mult_22/SUMB[62][55] ) );
  FA_X1 \mult_22/S2_62_54  ( .A(\mult_22/ab[62][54] ), .B(
        \mult_22/CARRYB[61][54] ), .CI(\mult_22/SUMB[61][55] ), .CO(
        \mult_22/CARRYB[62][54] ), .S(\mult_22/SUMB[62][54] ) );
  FA_X1 \mult_22/S2_62_53  ( .A(\mult_22/ab[62][53] ), .B(
        \mult_22/CARRYB[61][53] ), .CI(\mult_22/SUMB[61][54] ), .CO(
        \mult_22/CARRYB[62][53] ), .S(\mult_22/SUMB[62][53] ) );
  FA_X1 \mult_22/S2_62_52  ( .A(\mult_22/ab[62][52] ), .B(
        \mult_22/CARRYB[61][52] ), .CI(\mult_22/SUMB[61][53] ), .CO(
        \mult_22/CARRYB[62][52] ), .S(\mult_22/SUMB[62][52] ) );
  FA_X1 \mult_22/S2_62_51  ( .A(\mult_22/ab[62][51] ), .B(
        \mult_22/CARRYB[61][51] ), .CI(\mult_22/SUMB[61][52] ), .CO(
        \mult_22/CARRYB[62][51] ), .S(\mult_22/SUMB[62][51] ) );
  FA_X1 \mult_22/S2_62_50  ( .A(\mult_22/ab[62][50] ), .B(
        \mult_22/CARRYB[61][50] ), .CI(\mult_22/SUMB[61][51] ), .CO(
        \mult_22/CARRYB[62][50] ), .S(\mult_22/SUMB[62][50] ) );
  FA_X1 \mult_22/S2_62_49  ( .A(\mult_22/ab[62][49] ), .B(
        \mult_22/CARRYB[61][49] ), .CI(\mult_22/SUMB[61][50] ), .CO(
        \mult_22/CARRYB[62][49] ), .S(\mult_22/SUMB[62][49] ) );
  FA_X1 \mult_22/S2_62_48  ( .A(\mult_22/ab[62][48] ), .B(
        \mult_22/CARRYB[61][48] ), .CI(\mult_22/SUMB[61][49] ), .CO(
        \mult_22/CARRYB[62][48] ), .S(\mult_22/SUMB[62][48] ) );
  FA_X1 \mult_22/S2_62_47  ( .A(\mult_22/ab[62][47] ), .B(
        \mult_22/CARRYB[61][47] ), .CI(\mult_22/SUMB[61][48] ), .CO(
        \mult_22/CARRYB[62][47] ), .S(\mult_22/SUMB[62][47] ) );
  FA_X1 \mult_22/S2_62_46  ( .A(\mult_22/ab[62][46] ), .B(
        \mult_22/CARRYB[61][46] ), .CI(\mult_22/SUMB[61][47] ), .CO(
        \mult_22/CARRYB[62][46] ), .S(\mult_22/SUMB[62][46] ) );
  FA_X1 \mult_22/S2_62_45  ( .A(\mult_22/ab[62][45] ), .B(
        \mult_22/CARRYB[61][45] ), .CI(\mult_22/SUMB[61][46] ), .CO(
        \mult_22/CARRYB[62][45] ), .S(\mult_22/SUMB[62][45] ) );
  FA_X1 \mult_22/S2_62_44  ( .A(\mult_22/ab[62][44] ), .B(
        \mult_22/CARRYB[61][44] ), .CI(\mult_22/SUMB[61][45] ), .CO(
        \mult_22/CARRYB[62][44] ), .S(\mult_22/SUMB[62][44] ) );
  FA_X1 \mult_22/S2_62_43  ( .A(\mult_22/ab[62][43] ), .B(
        \mult_22/CARRYB[61][43] ), .CI(\mult_22/SUMB[61][44] ), .CO(
        \mult_22/CARRYB[62][43] ), .S(\mult_22/SUMB[62][43] ) );
  FA_X1 \mult_22/S2_62_42  ( .A(\mult_22/ab[62][42] ), .B(
        \mult_22/CARRYB[61][42] ), .CI(\mult_22/SUMB[61][43] ), .CO(
        \mult_22/CARRYB[62][42] ), .S(\mult_22/SUMB[62][42] ) );
  FA_X1 \mult_22/S2_62_41  ( .A(\mult_22/ab[62][41] ), .B(
        \mult_22/CARRYB[61][41] ), .CI(\mult_22/SUMB[61][42] ), .CO(
        \mult_22/CARRYB[62][41] ), .S(\mult_22/SUMB[62][41] ) );
  FA_X1 \mult_22/S2_62_40  ( .A(\mult_22/ab[62][40] ), .B(
        \mult_22/CARRYB[61][40] ), .CI(\mult_22/SUMB[61][41] ), .CO(
        \mult_22/CARRYB[62][40] ), .S(\mult_22/SUMB[62][40] ) );
  FA_X1 \mult_22/S2_62_39  ( .A(\mult_22/ab[62][39] ), .B(
        \mult_22/CARRYB[61][39] ), .CI(\mult_22/SUMB[61][40] ), .CO(
        \mult_22/CARRYB[62][39] ), .S(\mult_22/SUMB[62][39] ) );
  FA_X1 \mult_22/S2_62_38  ( .A(\mult_22/ab[62][38] ), .B(
        \mult_22/CARRYB[61][38] ), .CI(\mult_22/SUMB[61][39] ), .CO(
        \mult_22/CARRYB[62][38] ), .S(\mult_22/SUMB[62][38] ) );
  FA_X1 \mult_22/S2_62_37  ( .A(\mult_22/ab[62][37] ), .B(
        \mult_22/CARRYB[61][37] ), .CI(\mult_22/SUMB[61][38] ), .CO(
        \mult_22/CARRYB[62][37] ), .S(\mult_22/SUMB[62][37] ) );
  FA_X1 \mult_22/S2_62_36  ( .A(\mult_22/ab[62][36] ), .B(
        \mult_22/CARRYB[61][36] ), .CI(\mult_22/SUMB[61][37] ), .CO(
        \mult_22/CARRYB[62][36] ), .S(\mult_22/SUMB[62][36] ) );
  FA_X1 \mult_22/S2_62_35  ( .A(\mult_22/ab[62][35] ), .B(
        \mult_22/CARRYB[61][35] ), .CI(\mult_22/SUMB[61][36] ), .CO(
        \mult_22/CARRYB[62][35] ), .S(\mult_22/SUMB[62][35] ) );
  FA_X1 \mult_22/S2_62_34  ( .A(\mult_22/ab[62][34] ), .B(
        \mult_22/CARRYB[61][34] ), .CI(\mult_22/SUMB[61][35] ), .CO(
        \mult_22/CARRYB[62][34] ), .S(\mult_22/SUMB[62][34] ) );
  FA_X1 \mult_22/S2_62_33  ( .A(\mult_22/ab[62][33] ), .B(
        \mult_22/CARRYB[61][33] ), .CI(\mult_22/SUMB[61][34] ), .CO(
        \mult_22/CARRYB[62][33] ), .S(\mult_22/SUMB[62][33] ) );
  FA_X1 \mult_22/S2_62_32  ( .A(\mult_22/ab[62][32] ), .B(
        \mult_22/CARRYB[61][32] ), .CI(\mult_22/SUMB[61][33] ), .CO(
        \mult_22/CARRYB[62][32] ), .S(\mult_22/SUMB[62][32] ) );
  FA_X1 \mult_22/S2_62_31  ( .A(\mult_22/ab[62][31] ), .B(
        \mult_22/CARRYB[61][31] ), .CI(\mult_22/SUMB[61][32] ), .CO(
        \mult_22/CARRYB[62][31] ), .S(\mult_22/SUMB[62][31] ) );
  FA_X1 \mult_22/S2_62_30  ( .A(\mult_22/ab[62][30] ), .B(
        \mult_22/CARRYB[61][30] ), .CI(\mult_22/SUMB[61][31] ), .CO(
        \mult_22/CARRYB[62][30] ), .S(\mult_22/SUMB[62][30] ) );
  FA_X1 \mult_22/S2_62_29  ( .A(\mult_22/ab[62][29] ), .B(
        \mult_22/CARRYB[61][29] ), .CI(\mult_22/SUMB[61][30] ), .CO(
        \mult_22/CARRYB[62][29] ), .S(\mult_22/SUMB[62][29] ) );
  FA_X1 \mult_22/S2_62_28  ( .A(\mult_22/ab[62][28] ), .B(
        \mult_22/CARRYB[61][28] ), .CI(\mult_22/SUMB[61][29] ), .CO(
        \mult_22/CARRYB[62][28] ), .S(\mult_22/SUMB[62][28] ) );
  FA_X1 \mult_22/S2_62_27  ( .A(\mult_22/ab[62][27] ), .B(
        \mult_22/CARRYB[61][27] ), .CI(\mult_22/SUMB[61][28] ), .CO(
        \mult_22/CARRYB[62][27] ), .S(\mult_22/SUMB[62][27] ) );
  FA_X1 \mult_22/S2_62_26  ( .A(\mult_22/ab[62][26] ), .B(
        \mult_22/CARRYB[61][26] ), .CI(\mult_22/SUMB[61][27] ), .CO(
        \mult_22/CARRYB[62][26] ), .S(\mult_22/SUMB[62][26] ) );
  FA_X1 \mult_22/S2_62_25  ( .A(\mult_22/ab[62][25] ), .B(
        \mult_22/CARRYB[61][25] ), .CI(\mult_22/SUMB[61][26] ), .CO(
        \mult_22/CARRYB[62][25] ), .S(\mult_22/SUMB[62][25] ) );
  FA_X1 \mult_22/S2_62_24  ( .A(\mult_22/ab[62][24] ), .B(
        \mult_22/CARRYB[61][24] ), .CI(\mult_22/SUMB[61][25] ), .CO(
        \mult_22/CARRYB[62][24] ), .S(\mult_22/SUMB[62][24] ) );
  FA_X1 \mult_22/S2_62_23  ( .A(\mult_22/ab[62][23] ), .B(
        \mult_22/CARRYB[61][23] ), .CI(\mult_22/SUMB[61][24] ), .CO(
        \mult_22/CARRYB[62][23] ), .S(\mult_22/SUMB[62][23] ) );
  FA_X1 \mult_22/S2_62_22  ( .A(\mult_22/ab[62][22] ), .B(
        \mult_22/CARRYB[61][22] ), .CI(\mult_22/SUMB[61][23] ), .CO(
        \mult_22/CARRYB[62][22] ), .S(\mult_22/SUMB[62][22] ) );
  FA_X1 \mult_22/S2_62_21  ( .A(\mult_22/ab[62][21] ), .B(
        \mult_22/CARRYB[61][21] ), .CI(\mult_22/SUMB[61][22] ), .CO(
        \mult_22/CARRYB[62][21] ), .S(\mult_22/SUMB[62][21] ) );
  FA_X1 \mult_22/S2_62_20  ( .A(\mult_22/ab[62][20] ), .B(
        \mult_22/CARRYB[61][20] ), .CI(\mult_22/SUMB[61][21] ), .CO(
        \mult_22/CARRYB[62][20] ), .S(\mult_22/SUMB[62][20] ) );
  FA_X1 \mult_22/S2_62_19  ( .A(\mult_22/ab[62][19] ), .B(
        \mult_22/CARRYB[61][19] ), .CI(\mult_22/SUMB[61][20] ), .CO(
        \mult_22/CARRYB[62][19] ), .S(\mult_22/SUMB[62][19] ) );
  FA_X1 \mult_22/S2_62_18  ( .A(\mult_22/ab[62][18] ), .B(
        \mult_22/CARRYB[61][18] ), .CI(\mult_22/SUMB[61][19] ), .CO(
        \mult_22/CARRYB[62][18] ), .S(\mult_22/SUMB[62][18] ) );
  FA_X1 \mult_22/S2_62_17  ( .A(\mult_22/ab[62][17] ), .B(
        \mult_22/CARRYB[61][17] ), .CI(\mult_22/SUMB[61][18] ), .CO(
        \mult_22/CARRYB[62][17] ), .S(\mult_22/SUMB[62][17] ) );
  FA_X1 \mult_22/S2_62_16  ( .A(\mult_22/ab[62][16] ), .B(
        \mult_22/CARRYB[61][16] ), .CI(\mult_22/SUMB[61][17] ), .CO(
        \mult_22/CARRYB[62][16] ), .S(\mult_22/SUMB[62][16] ) );
  FA_X1 \mult_22/S2_62_15  ( .A(\mult_22/ab[62][15] ), .B(
        \mult_22/CARRYB[61][15] ), .CI(\mult_22/SUMB[61][16] ), .CO(
        \mult_22/CARRYB[62][15] ), .S(\mult_22/SUMB[62][15] ) );
  FA_X1 \mult_22/S2_62_14  ( .A(\mult_22/ab[62][14] ), .B(
        \mult_22/CARRYB[61][14] ), .CI(\mult_22/SUMB[61][15] ), .CO(
        \mult_22/CARRYB[62][14] ), .S(\mult_22/SUMB[62][14] ) );
  FA_X1 \mult_22/S2_62_13  ( .A(\mult_22/ab[62][13] ), .B(
        \mult_22/CARRYB[61][13] ), .CI(\mult_22/SUMB[61][14] ), .CO(
        \mult_22/CARRYB[62][13] ), .S(\mult_22/SUMB[62][13] ) );
  FA_X1 \mult_22/S2_62_12  ( .A(\mult_22/ab[62][12] ), .B(
        \mult_22/CARRYB[61][12] ), .CI(\mult_22/SUMB[61][13] ), .CO(
        \mult_22/CARRYB[62][12] ), .S(\mult_22/SUMB[62][12] ) );
  FA_X1 \mult_22/S2_62_11  ( .A(\mult_22/ab[62][11] ), .B(
        \mult_22/CARRYB[61][11] ), .CI(\mult_22/SUMB[61][12] ), .CO(
        \mult_22/CARRYB[62][11] ), .S(\mult_22/SUMB[62][11] ) );
  FA_X1 \mult_22/S2_62_10  ( .A(\mult_22/ab[62][10] ), .B(
        \mult_22/CARRYB[61][10] ), .CI(\mult_22/SUMB[61][11] ), .CO(
        \mult_22/CARRYB[62][10] ), .S(\mult_22/SUMB[62][10] ) );
  FA_X1 \mult_22/S2_62_9  ( .A(\mult_22/ab[62][9] ), .B(
        \mult_22/CARRYB[61][9] ), .CI(\mult_22/SUMB[61][10] ), .CO(
        \mult_22/CARRYB[62][9] ), .S(\mult_22/SUMB[62][9] ) );
  FA_X1 \mult_22/S2_62_8  ( .A(\mult_22/ab[62][8] ), .B(
        \mult_22/CARRYB[61][8] ), .CI(\mult_22/SUMB[61][9] ), .CO(
        \mult_22/CARRYB[62][8] ), .S(\mult_22/SUMB[62][8] ) );
  FA_X1 \mult_22/S2_62_7  ( .A(\mult_22/ab[62][7] ), .B(
        \mult_22/CARRYB[61][7] ), .CI(\mult_22/SUMB[61][8] ), .CO(
        \mult_22/CARRYB[62][7] ), .S(\mult_22/SUMB[62][7] ) );
  FA_X1 \mult_22/S2_62_6  ( .A(\mult_22/ab[62][6] ), .B(
        \mult_22/CARRYB[61][6] ), .CI(\mult_22/SUMB[61][7] ), .CO(
        \mult_22/CARRYB[62][6] ), .S(\mult_22/SUMB[62][6] ) );
  FA_X1 \mult_22/S2_62_5  ( .A(\mult_22/ab[62][5] ), .B(
        \mult_22/CARRYB[61][5] ), .CI(\mult_22/SUMB[61][6] ), .CO(
        \mult_22/CARRYB[62][5] ), .S(\mult_22/SUMB[62][5] ) );
  FA_X1 \mult_22/S2_62_4  ( .A(\mult_22/CARRYB[61][4] ), .B(
        \mult_22/ab[62][4] ), .CI(\mult_22/SUMB[61][5] ), .CO(
        \mult_22/CARRYB[62][4] ), .S(\mult_22/SUMB[62][4] ) );
  FA_X1 \mult_22/S2_62_3  ( .A(\mult_22/ab[62][3] ), .B(
        \mult_22/CARRYB[61][3] ), .CI(\mult_22/SUMB[61][4] ), .CO(
        \mult_22/CARRYB[62][3] ), .S(\mult_22/SUMB[62][3] ) );
  FA_X1 \mult_22/S2_62_2  ( .A(\mult_22/ab[62][2] ), .B(
        \mult_22/CARRYB[61][2] ), .CI(\mult_22/SUMB[61][3] ), .CO(
        \mult_22/CARRYB[62][2] ), .S(\mult_22/SUMB[62][2] ) );
  FA_X1 \mult_22/S2_62_1  ( .A(\mult_22/ab[62][1] ), .B(
        \mult_22/CARRYB[61][1] ), .CI(\mult_22/SUMB[61][2] ), .CO(
        \mult_22/CARRYB[62][1] ), .S(\mult_22/SUMB[62][1] ) );
  FA_X1 \mult_22/S1_62_0  ( .A(\mult_22/ab[62][0] ), .B(
        \mult_22/CARRYB[61][0] ), .CI(\mult_22/SUMB[61][1] ), .CO(
        \mult_22/CARRYB[62][0] ), .S(N190) );
  FA_X1 \mult_22/S5_62  ( .A(\mult_22/ab[63][62] ), .B(
        \mult_22/CARRYB[62][62] ), .CI(\mult_22/ab[62][63] ), .CO(
        \mult_22/CARRYB[63][62] ), .S(\mult_22/SUMB[63][62] ) );
  FA_X1 \mult_22/S4_61  ( .A(\mult_22/ab[63][61] ), .B(
        \mult_22/CARRYB[62][61] ), .CI(\mult_22/SUMB[62][62] ), .CO(
        \mult_22/CARRYB[63][61] ), .S(\mult_22/SUMB[63][61] ) );
  FA_X1 \mult_22/S4_60  ( .A(\mult_22/ab[63][60] ), .B(
        \mult_22/CARRYB[62][60] ), .CI(\mult_22/SUMB[62][61] ), .CO(
        \mult_22/CARRYB[63][60] ), .S(\mult_22/SUMB[63][60] ) );
  FA_X1 \mult_22/S4_59  ( .A(\mult_22/ab[63][59] ), .B(
        \mult_22/CARRYB[62][59] ), .CI(\mult_22/SUMB[62][60] ), .CO(
        \mult_22/CARRYB[63][59] ), .S(\mult_22/SUMB[63][59] ) );
  FA_X1 \mult_22/S4_58  ( .A(\mult_22/ab[63][58] ), .B(
        \mult_22/CARRYB[62][58] ), .CI(\mult_22/SUMB[62][59] ), .CO(
        \mult_22/CARRYB[63][58] ), .S(\mult_22/SUMB[63][58] ) );
  FA_X1 \mult_22/S4_57  ( .A(\mult_22/ab[63][57] ), .B(
        \mult_22/CARRYB[62][57] ), .CI(\mult_22/SUMB[62][58] ), .CO(
        \mult_22/CARRYB[63][57] ), .S(\mult_22/SUMB[63][57] ) );
  FA_X1 \mult_22/S4_56  ( .A(\mult_22/ab[63][56] ), .B(
        \mult_22/CARRYB[62][56] ), .CI(\mult_22/SUMB[62][57] ), .CO(
        \mult_22/CARRYB[63][56] ), .S(\mult_22/SUMB[63][56] ) );
  FA_X1 \mult_22/S4_55  ( .A(\mult_22/ab[63][55] ), .B(
        \mult_22/CARRYB[62][55] ), .CI(\mult_22/SUMB[62][56] ), .CO(
        \mult_22/CARRYB[63][55] ), .S(\mult_22/SUMB[63][55] ) );
  FA_X1 \mult_22/S4_54  ( .A(\mult_22/ab[63][54] ), .B(
        \mult_22/CARRYB[62][54] ), .CI(\mult_22/SUMB[62][55] ), .CO(
        \mult_22/CARRYB[63][54] ), .S(\mult_22/SUMB[63][54] ) );
  FA_X1 \mult_22/S4_53  ( .A(\mult_22/ab[63][53] ), .B(
        \mult_22/CARRYB[62][53] ), .CI(\mult_22/SUMB[62][54] ), .CO(
        \mult_22/CARRYB[63][53] ), .S(\mult_22/SUMB[63][53] ) );
  FA_X1 \mult_22/S4_52  ( .A(\mult_22/ab[63][52] ), .B(
        \mult_22/CARRYB[62][52] ), .CI(\mult_22/SUMB[62][53] ), .CO(
        \mult_22/CARRYB[63][52] ), .S(\mult_22/SUMB[63][52] ) );
  FA_X1 \mult_22/S4_51  ( .A(\mult_22/ab[63][51] ), .B(
        \mult_22/CARRYB[62][51] ), .CI(\mult_22/SUMB[62][52] ), .CO(
        \mult_22/CARRYB[63][51] ), .S(\mult_22/SUMB[63][51] ) );
  FA_X1 \mult_22/S4_50  ( .A(\mult_22/ab[63][50] ), .B(
        \mult_22/CARRYB[62][50] ), .CI(\mult_22/SUMB[62][51] ), .CO(
        \mult_22/CARRYB[63][50] ), .S(\mult_22/SUMB[63][50] ) );
  FA_X1 \mult_22/S4_49  ( .A(\mult_22/ab[63][49] ), .B(
        \mult_22/CARRYB[62][49] ), .CI(\mult_22/SUMB[62][50] ), .CO(
        \mult_22/CARRYB[63][49] ), .S(\mult_22/SUMB[63][49] ) );
  FA_X1 \mult_22/S4_48  ( .A(\mult_22/ab[63][48] ), .B(
        \mult_22/CARRYB[62][48] ), .CI(\mult_22/SUMB[62][49] ), .CO(
        \mult_22/CARRYB[63][48] ), .S(\mult_22/SUMB[63][48] ) );
  FA_X1 \mult_22/S4_47  ( .A(\mult_22/ab[63][47] ), .B(
        \mult_22/CARRYB[62][47] ), .CI(\mult_22/SUMB[62][48] ), .CO(
        \mult_22/CARRYB[63][47] ), .S(\mult_22/SUMB[63][47] ) );
  FA_X1 \mult_22/S4_46  ( .A(\mult_22/ab[63][46] ), .B(
        \mult_22/CARRYB[62][46] ), .CI(\mult_22/SUMB[62][47] ), .CO(
        \mult_22/CARRYB[63][46] ), .S(\mult_22/SUMB[63][46] ) );
  FA_X1 \mult_22/S4_45  ( .A(\mult_22/ab[63][45] ), .B(
        \mult_22/CARRYB[62][45] ), .CI(\mult_22/SUMB[62][46] ), .CO(
        \mult_22/CARRYB[63][45] ), .S(\mult_22/SUMB[63][45] ) );
  FA_X1 \mult_22/S4_44  ( .A(\mult_22/ab[63][44] ), .B(
        \mult_22/CARRYB[62][44] ), .CI(\mult_22/SUMB[62][45] ), .CO(
        \mult_22/CARRYB[63][44] ), .S(\mult_22/SUMB[63][44] ) );
  FA_X1 \mult_22/S4_43  ( .A(\mult_22/ab[63][43] ), .B(
        \mult_22/CARRYB[62][43] ), .CI(\mult_22/SUMB[62][44] ), .CO(
        \mult_22/CARRYB[63][43] ), .S(\mult_22/SUMB[63][43] ) );
  FA_X1 \mult_22/S4_42  ( .A(\mult_22/ab[63][42] ), .B(
        \mult_22/CARRYB[62][42] ), .CI(\mult_22/SUMB[62][43] ), .CO(
        \mult_22/CARRYB[63][42] ), .S(\mult_22/SUMB[63][42] ) );
  FA_X1 \mult_22/S4_41  ( .A(\mult_22/ab[63][41] ), .B(
        \mult_22/CARRYB[62][41] ), .CI(\mult_22/SUMB[62][42] ), .CO(
        \mult_22/CARRYB[63][41] ), .S(\mult_22/SUMB[63][41] ) );
  FA_X1 \mult_22/S4_40  ( .A(\mult_22/ab[63][40] ), .B(
        \mult_22/CARRYB[62][40] ), .CI(\mult_22/SUMB[62][41] ), .CO(
        \mult_22/CARRYB[63][40] ), .S(\mult_22/SUMB[63][40] ) );
  FA_X1 \mult_22/S4_39  ( .A(\mult_22/ab[63][39] ), .B(
        \mult_22/CARRYB[62][39] ), .CI(\mult_22/SUMB[62][40] ), .CO(
        \mult_22/CARRYB[63][39] ), .S(\mult_22/SUMB[63][39] ) );
  FA_X1 \mult_22/S4_38  ( .A(\mult_22/ab[63][38] ), .B(
        \mult_22/CARRYB[62][38] ), .CI(\mult_22/SUMB[62][39] ), .CO(
        \mult_22/CARRYB[63][38] ), .S(\mult_22/SUMB[63][38] ) );
  FA_X1 \mult_22/S4_37  ( .A(\mult_22/ab[63][37] ), .B(
        \mult_22/CARRYB[62][37] ), .CI(\mult_22/SUMB[62][38] ), .CO(
        \mult_22/CARRYB[63][37] ), .S(\mult_22/SUMB[63][37] ) );
  FA_X1 \mult_22/S4_36  ( .A(\mult_22/ab[63][36] ), .B(
        \mult_22/CARRYB[62][36] ), .CI(\mult_22/SUMB[62][37] ), .CO(
        \mult_22/CARRYB[63][36] ), .S(\mult_22/SUMB[63][36] ) );
  FA_X1 \mult_22/S4_35  ( .A(\mult_22/ab[63][35] ), .B(
        \mult_22/CARRYB[62][35] ), .CI(\mult_22/SUMB[62][36] ), .CO(
        \mult_22/CARRYB[63][35] ), .S(\mult_22/SUMB[63][35] ) );
  FA_X1 \mult_22/S4_34  ( .A(\mult_22/ab[63][34] ), .B(
        \mult_22/CARRYB[62][34] ), .CI(\mult_22/SUMB[62][35] ), .CO(
        \mult_22/CARRYB[63][34] ), .S(\mult_22/SUMB[63][34] ) );
  FA_X1 \mult_22/S4_33  ( .A(\mult_22/ab[63][33] ), .B(
        \mult_22/CARRYB[62][33] ), .CI(\mult_22/SUMB[62][34] ), .CO(
        \mult_22/CARRYB[63][33] ), .S(\mult_22/SUMB[63][33] ) );
  FA_X1 \mult_22/S4_32  ( .A(\mult_22/ab[63][32] ), .B(
        \mult_22/CARRYB[62][32] ), .CI(\mult_22/SUMB[62][33] ), .CO(
        \mult_22/CARRYB[63][32] ), .S(\mult_22/SUMB[63][32] ) );
  FA_X1 \mult_22/S4_31  ( .A(\mult_22/ab[63][31] ), .B(
        \mult_22/CARRYB[62][31] ), .CI(\mult_22/SUMB[62][32] ), .CO(
        \mult_22/CARRYB[63][31] ), .S(\mult_22/SUMB[63][31] ) );
  FA_X1 \mult_22/S4_30  ( .A(\mult_22/ab[63][30] ), .B(
        \mult_22/CARRYB[62][30] ), .CI(\mult_22/SUMB[62][31] ), .CO(
        \mult_22/CARRYB[63][30] ), .S(\mult_22/SUMB[63][30] ) );
  FA_X1 \mult_22/S4_29  ( .A(\mult_22/ab[63][29] ), .B(
        \mult_22/CARRYB[62][29] ), .CI(\mult_22/SUMB[62][30] ), .CO(
        \mult_22/CARRYB[63][29] ), .S(\mult_22/SUMB[63][29] ) );
  FA_X1 \mult_22/S4_28  ( .A(\mult_22/ab[63][28] ), .B(
        \mult_22/CARRYB[62][28] ), .CI(\mult_22/SUMB[62][29] ), .CO(
        \mult_22/CARRYB[63][28] ), .S(\mult_22/SUMB[63][28] ) );
  FA_X1 \mult_22/S4_27  ( .A(\mult_22/ab[63][27] ), .B(
        \mult_22/CARRYB[62][27] ), .CI(\mult_22/SUMB[62][28] ), .CO(
        \mult_22/CARRYB[63][27] ), .S(\mult_22/SUMB[63][27] ) );
  FA_X1 \mult_22/S4_26  ( .A(\mult_22/ab[63][26] ), .B(
        \mult_22/CARRYB[62][26] ), .CI(\mult_22/SUMB[62][27] ), .CO(
        \mult_22/CARRYB[63][26] ), .S(\mult_22/SUMB[63][26] ) );
  FA_X1 \mult_22/S4_25  ( .A(\mult_22/ab[63][25] ), .B(
        \mult_22/CARRYB[62][25] ), .CI(\mult_22/SUMB[62][26] ), .CO(
        \mult_22/CARRYB[63][25] ), .S(\mult_22/SUMB[63][25] ) );
  FA_X1 \mult_22/S4_24  ( .A(\mult_22/ab[63][24] ), .B(
        \mult_22/CARRYB[62][24] ), .CI(\mult_22/SUMB[62][25] ), .CO(
        \mult_22/CARRYB[63][24] ), .S(\mult_22/SUMB[63][24] ) );
  FA_X1 \mult_22/S4_23  ( .A(\mult_22/ab[63][23] ), .B(
        \mult_22/CARRYB[62][23] ), .CI(\mult_22/SUMB[62][24] ), .CO(
        \mult_22/CARRYB[63][23] ), .S(\mult_22/SUMB[63][23] ) );
  FA_X1 \mult_22/S4_22  ( .A(\mult_22/ab[63][22] ), .B(
        \mult_22/CARRYB[62][22] ), .CI(\mult_22/SUMB[62][23] ), .CO(
        \mult_22/CARRYB[63][22] ), .S(\mult_22/SUMB[63][22] ) );
  FA_X1 \mult_22/S4_21  ( .A(\mult_22/ab[63][21] ), .B(
        \mult_22/CARRYB[62][21] ), .CI(\mult_22/SUMB[62][22] ), .CO(
        \mult_22/CARRYB[63][21] ), .S(\mult_22/SUMB[63][21] ) );
  FA_X1 \mult_22/S4_20  ( .A(\mult_22/ab[63][20] ), .B(
        \mult_22/CARRYB[62][20] ), .CI(\mult_22/SUMB[62][21] ), .CO(
        \mult_22/CARRYB[63][20] ), .S(\mult_22/SUMB[63][20] ) );
  FA_X1 \mult_22/S4_19  ( .A(\mult_22/ab[63][19] ), .B(
        \mult_22/CARRYB[62][19] ), .CI(\mult_22/SUMB[62][20] ), .CO(
        \mult_22/CARRYB[63][19] ), .S(\mult_22/SUMB[63][19] ) );
  FA_X1 \mult_22/S4_18  ( .A(\mult_22/ab[63][18] ), .B(
        \mult_22/CARRYB[62][18] ), .CI(\mult_22/SUMB[62][19] ), .CO(
        \mult_22/CARRYB[63][18] ), .S(\mult_22/SUMB[63][18] ) );
  FA_X1 \mult_22/S4_17  ( .A(\mult_22/ab[63][17] ), .B(
        \mult_22/CARRYB[62][17] ), .CI(\mult_22/SUMB[62][18] ), .CO(
        \mult_22/CARRYB[63][17] ), .S(\mult_22/SUMB[63][17] ) );
  FA_X1 \mult_22/S4_16  ( .A(\mult_22/ab[63][16] ), .B(
        \mult_22/CARRYB[62][16] ), .CI(\mult_22/SUMB[62][17] ), .CO(
        \mult_22/CARRYB[63][16] ), .S(\mult_22/SUMB[63][16] ) );
  FA_X1 \mult_22/S4_15  ( .A(\mult_22/ab[63][15] ), .B(
        \mult_22/CARRYB[62][15] ), .CI(\mult_22/SUMB[62][16] ), .CO(
        \mult_22/CARRYB[63][15] ), .S(\mult_22/SUMB[63][15] ) );
  FA_X1 \mult_22/S4_14  ( .A(\mult_22/ab[63][14] ), .B(
        \mult_22/CARRYB[62][14] ), .CI(\mult_22/SUMB[62][15] ), .CO(
        \mult_22/CARRYB[63][14] ), .S(\mult_22/SUMB[63][14] ) );
  FA_X1 \mult_22/S4_13  ( .A(\mult_22/ab[63][13] ), .B(
        \mult_22/CARRYB[62][13] ), .CI(\mult_22/SUMB[62][14] ), .CO(
        \mult_22/CARRYB[63][13] ), .S(\mult_22/SUMB[63][13] ) );
  FA_X1 \mult_22/S4_12  ( .A(\mult_22/ab[63][12] ), .B(
        \mult_22/CARRYB[62][12] ), .CI(\mult_22/SUMB[62][13] ), .CO(
        \mult_22/CARRYB[63][12] ), .S(\mult_22/SUMB[63][12] ) );
  FA_X1 \mult_22/S4_11  ( .A(\mult_22/ab[63][11] ), .B(
        \mult_22/CARRYB[62][11] ), .CI(\mult_22/SUMB[62][12] ), .CO(
        \mult_22/CARRYB[63][11] ), .S(\mult_22/SUMB[63][11] ) );
  FA_X1 \mult_22/S4_10  ( .A(\mult_22/ab[63][10] ), .B(
        \mult_22/CARRYB[62][10] ), .CI(\mult_22/SUMB[62][11] ), .CO(
        \mult_22/CARRYB[63][10] ), .S(\mult_22/SUMB[63][10] ) );
  FA_X1 \mult_22/S4_9  ( .A(\mult_22/ab[63][9] ), .B(\mult_22/CARRYB[62][9] ), 
        .CI(\mult_22/SUMB[62][10] ), .CO(\mult_22/CARRYB[63][9] ), .S(
        \mult_22/SUMB[63][9] ) );
  FA_X1 \mult_22/S4_8  ( .A(\mult_22/ab[63][8] ), .B(\mult_22/CARRYB[62][8] ), 
        .CI(\mult_22/SUMB[62][9] ), .CO(\mult_22/CARRYB[63][8] ), .S(
        \mult_22/SUMB[63][8] ) );
  FA_X1 \mult_22/S4_7  ( .A(\mult_22/ab[63][7] ), .B(\mult_22/CARRYB[62][7] ), 
        .CI(\mult_22/SUMB[62][8] ), .CO(\mult_22/CARRYB[63][7] ), .S(
        \mult_22/SUMB[63][7] ) );
  FA_X1 \mult_22/S4_6  ( .A(\mult_22/ab[63][6] ), .B(\mult_22/CARRYB[62][6] ), 
        .CI(\mult_22/SUMB[62][7] ), .CO(\mult_22/CARRYB[63][6] ), .S(
        \mult_22/SUMB[63][6] ) );
  FA_X1 \mult_22/S4_5  ( .A(\mult_22/ab[63][5] ), .B(\mult_22/CARRYB[62][5] ), 
        .CI(\mult_22/SUMB[62][6] ), .CO(\mult_22/CARRYB[63][5] ), .S(
        \mult_22/SUMB[63][5] ) );
  FA_X1 \mult_22/S4_4  ( .A(\mult_22/CARRYB[62][4] ), .B(\mult_22/ab[63][4] ), 
        .CI(\mult_22/SUMB[62][5] ), .CO(\mult_22/CARRYB[63][4] ), .S(
        \mult_22/SUMB[63][4] ) );
  FA_X1 \mult_22/S4_3  ( .A(\mult_22/CARRYB[62][3] ), .B(\mult_22/ab[63][3] ), 
        .CI(\mult_22/SUMB[62][4] ), .CO(\mult_22/CARRYB[63][3] ), .S(
        \mult_22/SUMB[63][3] ) );
  FA_X1 \mult_22/S4_2  ( .A(\mult_22/ab[63][2] ), .B(\mult_22/CARRYB[62][2] ), 
        .CI(\mult_22/SUMB[62][3] ), .CO(\mult_22/CARRYB[63][2] ), .S(
        \mult_22/SUMB[63][2] ) );
  FA_X1 \mult_22/S4_1  ( .A(\mult_22/ab[63][1] ), .B(\mult_22/CARRYB[62][1] ), 
        .CI(\mult_22/SUMB[62][2] ), .CO(\mult_22/CARRYB[63][1] ), .S(
        \mult_22/SUMB[63][1] ) );
  FA_X1 \mult_22/S4_0  ( .A(\mult_22/ab[63][0] ), .B(\mult_22/CARRYB[62][0] ), 
        .CI(\mult_22/SUMB[62][1] ), .CO(\mult_22/CARRYB[63][0] ), .S(N191) );
  AOI21_X2 U6544 ( .B1(\mult_22/CARRYB[63][38] ), .B2(\mult_22/SUMB[63][39] ), 
        .A(n1415), .ZN(n1400) );
  AND2_X2 U6590 ( .A1(n1479), .A2(n1478), .ZN(n1466) );
  NOR2_X2 U6595 ( .A1(n1483), .A2(n1484), .ZN(n1467) );
  NOR2_X2 U6629 ( .A1(n1530), .A2(n1531), .ZN(n1519) );
  NOR2_X2 U6669 ( .A1(n1579), .A2(n1580), .ZN(n1563) );
  AOI21_X2 U6688 ( .B1(\mult_22/CARRYB[63][6] ), .B2(\mult_22/SUMB[63][7] ), 
        .A(n1603), .ZN(n1590) );
  XOR2_X1 U7280 ( .A(n810), .B(n811), .Z(\mult_22/n99 ) );
  XOR2_X1 U7281 ( .A(n812), .B(n813), .Z(\mult_22/n98 ) );
  XOR2_X1 U7282 ( .A(n814), .B(n815), .Z(\mult_22/n97 ) );
  XOR2_X1 U7283 ( .A(n816), .B(n817), .Z(\mult_22/n96 ) );
  XOR2_X1 U7284 ( .A(n818), .B(n819), .Z(\mult_22/n95 ) );
  XOR2_X1 U7285 ( .A(n820), .B(n821), .Z(\mult_22/n94 ) );
  XOR2_X1 U7286 ( .A(n822), .B(n823), .Z(\mult_22/n93 ) );
  XOR2_X1 U7287 ( .A(n824), .B(n825), .Z(\mult_22/n92 ) );
  XOR2_X1 U7288 ( .A(n826), .B(n827), .Z(\mult_22/n91 ) );
  XOR2_X1 U7289 ( .A(n828), .B(n829), .Z(\mult_22/n90 ) );
  XOR2_X1 U7290 ( .A(n831), .B(n832), .Z(\mult_22/n89 ) );
  XOR2_X1 U7291 ( .A(n833), .B(n834), .Z(\mult_22/n88 ) );
  XOR2_X1 U7292 ( .A(n835), .B(n836), .Z(\mult_22/n87 ) );
  XOR2_X1 U7293 ( .A(n837), .B(n838), .Z(\mult_22/n86 ) );
  XOR2_X1 U7294 ( .A(n839), .B(n840), .Z(\mult_22/n85 ) );
  XOR2_X1 U7295 ( .A(n841), .B(n842), .Z(\mult_22/n84 ) );
  XOR2_X1 U7296 ( .A(n843), .B(n844), .Z(\mult_22/n83 ) );
  XOR2_X1 U7297 ( .A(n845), .B(n846), .Z(\mult_22/n82 ) );
  XOR2_X1 U7298 ( .A(n847), .B(n848), .Z(\mult_22/n81 ) );
  XOR2_X1 U7299 ( .A(n849), .B(n850), .Z(\mult_22/n80 ) );
  XOR2_X1 U7300 ( .A(n852), .B(n853), .Z(\mult_22/n79 ) );
  XOR2_X1 U7301 ( .A(n854), .B(n855), .Z(\mult_22/n78 ) );
  XOR2_X1 U7302 ( .A(n856), .B(n857), .Z(\mult_22/n77 ) );
  XOR2_X1 U7303 ( .A(n858), .B(n859), .Z(\mult_22/n76 ) );
  XOR2_X1 U7304 ( .A(n860), .B(n861), .Z(\mult_22/n75 ) );
  XOR2_X1 U7305 ( .A(n862), .B(n863), .Z(\mult_22/n74 ) );
  XOR2_X1 U7306 ( .A(n864), .B(n865), .Z(\mult_22/n73 ) );
  XOR2_X1 U7307 ( .A(n866), .B(n867), .Z(\mult_22/n72 ) );
  XOR2_X1 U7308 ( .A(n868), .B(n869), .Z(\mult_22/n71 ) );
  XOR2_X1 U7309 ( .A(n870), .B(n871), .Z(\mult_22/n70 ) );
  XOR2_X1 U7310 ( .A(n873), .B(n874), .Z(\mult_22/n69 ) );
  XOR2_X1 U7311 ( .A(n876), .B(n877), .Z(\mult_22/n66 ) );
  XOR2_X1 U7312 ( .A(n878), .B(n879), .Z(\mult_22/n65 ) );
  XOR2_X1 U7313 ( .A(n880), .B(n881), .Z(\mult_22/n64 ) );
  XOR2_X1 U7314 ( .A(n851), .B(n882), .Z(\mult_22/n63 ) );
  XOR2_X1 U7315 ( .A(n872), .B(n883), .Z(\mult_22/n62 ) );
  XOR2_X1 U7316 ( .A(n884), .B(n885), .Z(\mult_22/n61 ) );
  XOR2_X1 U7320 ( .A(n909), .B(n910), .Z(\mult_22/n195 ) );
  XOR2_X1 U7321 ( .A(n911), .B(n912), .Z(\mult_22/n194 ) );
  XOR2_X1 U7322 ( .A(n886), .B(n913), .Z(\mult_22/n159 ) );
  XOR2_X1 U7323 ( .A(n830), .B(n914), .Z(\mult_22/n13 ) );
  XOR2_X1 U7324 ( .A(n892), .B(n915), .Z(\mult_22/n12 ) );
  XOR2_X1 U7325 ( .A(n888), .B(n916), .Z(\mult_22/n114 ) );
  XOR2_X1 U7326 ( .A(n875), .B(n917), .Z(\mult_22/n113 ) );
  XOR2_X1 U7327 ( .A(n889), .B(n918), .Z(\mult_22/n112 ) );
  XOR2_X1 U7328 ( .A(n890), .B(n919), .Z(\mult_22/n111 ) );
  XOR2_X1 U7329 ( .A(n891), .B(n920), .Z(\mult_22/n110 ) );
  XOR2_X1 U7330 ( .A(n893), .B(n921), .Z(\mult_22/n109 ) );
  XOR2_X1 U7331 ( .A(n894), .B(n922), .Z(\mult_22/n108 ) );
  XOR2_X1 U7332 ( .A(n895), .B(n923), .Z(\mult_22/n107 ) );
  XOR2_X1 U7333 ( .A(n896), .B(n924), .Z(\mult_22/n106 ) );
  XOR2_X1 U7334 ( .A(n897), .B(n925), .Z(\mult_22/n105 ) );
  XOR2_X1 U7335 ( .A(n898), .B(n926), .Z(\mult_22/n104 ) );
  XOR2_X1 U7336 ( .A(n899), .B(n927), .Z(\mult_22/n103 ) );
  XOR2_X1 U7337 ( .A(n900), .B(n928), .Z(\mult_22/n102 ) );
  XOR2_X1 U7338 ( .A(n905), .B(n929), .Z(\mult_22/n101 ) );
  XOR2_X1 U7339 ( .A(n906), .B(n930), .Z(\mult_22/n100 ) );
  XOR2_X1 U7350 ( .A(n942), .B(n941), .Z(\mult_22/SUMB[26][34] ) );
  NAND3_X1 U7363 ( .A1(reg_mid_0[21]), .A2(reg_mid_1[36]), .A3(
        \mult_22/CARRYB[20][36] ), .ZN(n953) );
  XOR2_X1 U7364 ( .A(n981), .B(n982), .Z(\mult_20/n63 ) );
  XOR2_X1 U7365 ( .A(n983), .B(n984), .Z(\mult_20/n62 ) );
  XOR2_X1 U7366 ( .A(n985), .B(n986), .Z(\mult_20/n61 ) );
  XOR2_X1 U7367 ( .A(n987), .B(n988), .Z(\mult_20/n60 ) );
  XOR2_X1 U7368 ( .A(n990), .B(n991), .Z(\mult_20/n59 ) );
  XOR2_X1 U7369 ( .A(n992), .B(n993), .Z(\mult_20/n58 ) );
  XOR2_X1 U7370 ( .A(n994), .B(n995), .Z(\mult_20/n57 ) );
  XOR2_X1 U7371 ( .A(n996), .B(n997), .Z(\mult_20/n56 ) );
  XOR2_X1 U7372 ( .A(n998), .B(n999), .Z(\mult_20/n55 ) );
  XOR2_X1 U7373 ( .A(n1000), .B(n1001), .Z(\mult_20/n54 ) );
  XOR2_X1 U7374 ( .A(n1002), .B(n1003), .Z(\mult_20/n53 ) );
  XOR2_X1 U7375 ( .A(n1004), .B(n1005), .Z(\mult_20/n52 ) );
  XOR2_X1 U7376 ( .A(n1006), .B(n1007), .Z(\mult_20/n51 ) );
  XOR2_X1 U7377 ( .A(n1008), .B(n1009), .Z(\mult_20/n50 ) );
  XOR2_X1 U7378 ( .A(n1011), .B(n1012), .Z(\mult_20/n49 ) );
  XOR2_X1 U7379 ( .A(n1013), .B(n1014), .Z(\mult_20/n48 ) );
  XOR2_X1 U7380 ( .A(n1015), .B(n1016), .Z(\mult_20/n47 ) );
  XOR2_X1 U7381 ( .A(n1017), .B(n1018), .Z(\mult_20/n46 ) );
  XOR2_X1 U7382 ( .A(n1019), .B(n1020), .Z(\mult_20/n45 ) );
  XOR2_X1 U7383 ( .A(n1021), .B(n1022), .Z(\mult_20/n44 ) );
  XOR2_X1 U7384 ( .A(n1023), .B(n1024), .Z(\mult_20/n43 ) );
  XOR2_X1 U7385 ( .A(n1025), .B(n1026), .Z(\mult_20/n42 ) );
  XOR2_X1 U7386 ( .A(n978), .B(n1027), .Z(\mult_20/n41 ) );
  XOR2_X1 U7387 ( .A(n979), .B(n1028), .Z(\mult_20/n40 ) );
  XOR2_X1 U7388 ( .A(n980), .B(n1030), .Z(\mult_20/n39 ) );
  XOR2_X1 U7389 ( .A(n989), .B(n1031), .Z(\mult_20/n38 ) );
  XOR2_X1 U7390 ( .A(n1010), .B(n1032), .Z(\mult_20/n37 ) );
  XOR2_X1 U7391 ( .A(n1029), .B(n1033), .Z(\mult_20/n36 ) );
  XOR2_X1 U7392 ( .A(n1034), .B(n1035), .Z(\mult_20/n35 ) );
  XOR2_X1 U7393 ( .A(n1036), .B(n1037), .Z(\mult_20/n34 ) );
  XOR2_X1 U7394 ( .A(n1042), .B(n1043), .Z(\mult_19/n63 ) );
  XOR2_X1 U7395 ( .A(n1044), .B(n1045), .Z(\mult_19/n62 ) );
  XOR2_X1 U7396 ( .A(n1046), .B(n1047), .Z(\mult_19/n61 ) );
  XOR2_X1 U7397 ( .A(n1048), .B(n1049), .Z(\mult_19/n60 ) );
  XOR2_X1 U7398 ( .A(n1051), .B(n1052), .Z(\mult_19/n59 ) );
  XOR2_X1 U7399 ( .A(n1053), .B(n1054), .Z(\mult_19/n58 ) );
  XOR2_X1 U7400 ( .A(n1055), .B(n1056), .Z(\mult_19/n57 ) );
  XOR2_X1 U7401 ( .A(n1057), .B(n1058), .Z(\mult_19/n56 ) );
  XOR2_X1 U7402 ( .A(n1059), .B(n1060), .Z(\mult_19/n55 ) );
  XOR2_X1 U7403 ( .A(n1061), .B(n1062), .Z(\mult_19/n54 ) );
  XOR2_X1 U7404 ( .A(n1063), .B(n1064), .Z(\mult_19/n53 ) );
  XOR2_X1 U7405 ( .A(n1065), .B(n1066), .Z(\mult_19/n52 ) );
  XOR2_X1 U7406 ( .A(n1067), .B(n1068), .Z(\mult_19/n51 ) );
  XOR2_X1 U7407 ( .A(n1069), .B(n1070), .Z(\mult_19/n50 ) );
  XOR2_X1 U7408 ( .A(n1072), .B(n1073), .Z(\mult_19/n49 ) );
  XOR2_X1 U7409 ( .A(n1074), .B(n1075), .Z(\mult_19/n48 ) );
  XOR2_X1 U7410 ( .A(n1076), .B(n1077), .Z(\mult_19/n47 ) );
  XOR2_X1 U7411 ( .A(n1078), .B(n1079), .Z(\mult_19/n46 ) );
  XOR2_X1 U7412 ( .A(n1080), .B(n1081), .Z(\mult_19/n45 ) );
  XOR2_X1 U7413 ( .A(n1082), .B(n1083), .Z(\mult_19/n44 ) );
  XOR2_X1 U7414 ( .A(n1084), .B(n1085), .Z(\mult_19/n43 ) );
  XOR2_X1 U7415 ( .A(n1086), .B(n1087), .Z(\mult_19/n42 ) );
  XOR2_X1 U7416 ( .A(n1039), .B(n1088), .Z(\mult_19/n41 ) );
  XOR2_X1 U7417 ( .A(n1040), .B(n1089), .Z(\mult_19/n40 ) );
  XOR2_X1 U7418 ( .A(n1041), .B(n1091), .Z(\mult_19/n39 ) );
  XOR2_X1 U7419 ( .A(n1050), .B(n1092), .Z(\mult_19/n38 ) );
  XOR2_X1 U7420 ( .A(n1071), .B(n1093), .Z(\mult_19/n37 ) );
  XOR2_X1 U7421 ( .A(n1090), .B(n1094), .Z(\mult_19/n36 ) );
  XOR2_X1 U7422 ( .A(n1095), .B(n1096), .Z(\mult_19/n35 ) );
  XOR2_X1 U7423 ( .A(n1097), .B(n1098), .Z(\mult_19/n34 ) );
  XOR2_X1 U7424 ( .A(n1100), .B(n1101), .Z(N99) );
  XOR2_X1 U7425 ( .A(n1103), .B(n1104), .Z(N98) );
  XOR2_X1 U7426 ( .A(\mult_20/SUMB[31][1] ), .B(\mult_20/CARRYB[31][0] ), .Z(
        N96) );
  XOR2_X1 U7427 ( .A(n1038), .B(n1108), .Z(N65) );
  XOR2_X1 U7428 ( .A(n1113), .B(n1109), .Z(N62) );
  NAND3_X1 U7429 ( .A1(\mult_19/SUMB[31][30] ), .A2(n488), .A3(
        \mult_19/CARRYB[31][29] ), .ZN(n1112) );
  XOR2_X1 U7430 ( .A(n1111), .B(\mult_19/CARRYB[31][30] ), .Z(n1110) );
  XOR2_X1 U7431 ( .A(n1125), .B(n1121), .Z(N60) );
  NAND3_X1 U7432 ( .A1(\mult_19/SUMB[31][28] ), .A2(n1124), .A3(
        \mult_19/CARRYB[31][27] ), .ZN(n1123) );
  XOR2_X1 U7433 ( .A(\mult_19/CARRYB[31][28] ), .B(\mult_19/SUMB[31][29] ), 
        .Z(n1124) );
  XOR2_X1 U7434 ( .A(n1137), .B(n1133), .Z(N58) );
  NAND3_X1 U7435 ( .A1(\mult_19/SUMB[31][26] ), .A2(n1136), .A3(
        \mult_19/CARRYB[31][25] ), .ZN(n1135) );
  XOR2_X1 U7436 ( .A(\mult_19/CARRYB[31][26] ), .B(\mult_19/SUMB[31][27] ), 
        .Z(n1136) );
  XOR2_X1 U7437 ( .A(n1149), .B(n1145), .Z(N56) );
  NAND3_X1 U7438 ( .A1(\mult_19/SUMB[31][24] ), .A2(n1148), .A3(
        \mult_19/CARRYB[31][23] ), .ZN(n1147) );
  XOR2_X1 U7439 ( .A(\mult_19/CARRYB[31][24] ), .B(\mult_19/SUMB[31][25] ), 
        .Z(n1148) );
  XOR2_X1 U7440 ( .A(n1151), .B(n1156), .Z(N55) );
  NAND3_X1 U7441 ( .A1(\mult_19/SUMB[31][22] ), .A2(n1161), .A3(
        \mult_19/CARRYB[31][21] ), .ZN(n1159) );
  XOR2_X1 U7442 ( .A(\mult_19/CARRYB[31][22] ), .B(\mult_19/SUMB[31][23] ), 
        .Z(n1161) );
  XOR2_X1 U7443 ( .A(n1163), .B(n1167), .Z(N53) );
  XOR2_X1 U7444 ( .A(n1170), .B(n1171), .Z(N52) );
  NAND3_X1 U7445 ( .A1(\mult_19/SUMB[31][20] ), .A2(n1172), .A3(
        \mult_19/CARRYB[31][19] ), .ZN(n1169) );
  XOR2_X1 U7446 ( .A(\mult_19/CARRYB[31][20] ), .B(\mult_19/SUMB[31][21] ), 
        .Z(n1172) );
  XOR2_X1 U7447 ( .A(n1178), .B(n1174), .Z(N51) );
  XOR2_X1 U7448 ( .A(\mult_19/CARRYB[31][19] ), .B(\mult_19/SUMB[31][20] ), 
        .Z(n1177) );
  XOR2_X1 U7449 ( .A(n1179), .B(n1182), .Z(N50) );
  XOR2_X1 U7450 ( .A(\mult_19/CARRYB[31][18] ), .B(\mult_19/SUMB[31][19] ), 
        .Z(n1183) );
  XOR2_X1 U7451 ( .A(n1187), .B(n1184), .Z(N49) );
  NAND3_X1 U7452 ( .A1(\mult_19/SUMB[31][17] ), .A2(n1191), .A3(
        \mult_19/CARRYB[31][16] ), .ZN(n1186) );
  XOR2_X1 U7453 ( .A(\mult_19/CARRYB[31][17] ), .B(\mult_19/SUMB[31][18] ), 
        .Z(n1191) );
  XOR2_X1 U7454 ( .A(n1188), .B(n1192), .Z(N48) );
  XOR2_X1 U7455 ( .A(\mult_19/CARRYB[31][16] ), .B(\mult_19/SUMB[31][17] ), 
        .Z(n1193) );
  XOR2_X1 U7456 ( .A(\mult_19/CARRYB[31][15] ), .B(\mult_19/SUMB[31][16] ), 
        .Z(n1199) );
  XOR2_X1 U7457 ( .A(n1200), .B(n1203), .Z(N46) );
  XOR2_X1 U7458 ( .A(\mult_19/CARRYB[31][14] ), .B(\mult_19/SUMB[31][15] ), 
        .Z(n1204) );
  NAND3_X1 U7459 ( .A1(n502), .A2(n1213), .A3(n1214), .ZN(n1211) );
  XOR2_X1 U7460 ( .A(n1215), .B(n1216), .Z(N45) );
  NAND3_X1 U7461 ( .A1(\mult_19/CARRYB[31][12] ), .A2(n1219), .A3(
        \mult_19/SUMB[31][13] ), .ZN(n1207) );
  XOR2_X1 U7462 ( .A(\mult_19/CARRYB[31][13] ), .B(\mult_19/SUMB[31][14] ), 
        .Z(n1219) );
  XOR2_X1 U7463 ( .A(n1217), .B(n1220), .Z(N44) );
  XOR2_X1 U7464 ( .A(\mult_19/CARRYB[31][12] ), .B(\mult_19/SUMB[31][13] ), 
        .Z(n1221) );
  XOR2_X1 U7465 ( .A(n1223), .B(n1222), .Z(N43) );
  NAND3_X1 U7466 ( .A1(\mult_19/CARRYB[31][10] ), .A2(n1225), .A3(
        \mult_19/SUMB[31][11] ), .ZN(n1212) );
  XOR2_X1 U7467 ( .A(\mult_19/CARRYB[31][11] ), .B(\mult_19/SUMB[31][12] ), 
        .Z(n1225) );
  NAND3_X1 U7469 ( .A1(n1233), .A2(n1234), .A3(n1235), .ZN(n1232) );
  XOR2_X1 U7470 ( .A(n1242), .B(n1243), .Z(N41) );
  XOR2_X1 U7471 ( .A(n1244), .B(n1245), .Z(N40) );
  XOR2_X1 U7472 ( .A(\mult_19/CARRYB[31][8] ), .B(\mult_19/SUMB[31][9] ), .Z(
        n1246) );
  XOR2_X1 U7473 ( .A(n1248), .B(n1247), .Z(N39) );
  NAND3_X1 U7474 ( .A1(\mult_19/CARRYB[31][6] ), .A2(n1250), .A3(
        \mult_19/SUMB[31][7] ), .ZN(n1240) );
  XOR2_X1 U7475 ( .A(\mult_19/CARRYB[31][7] ), .B(\mult_19/SUMB[31][8] ), .Z(
        n1250) );
  XOR2_X1 U7476 ( .A(n1233), .B(n1251), .Z(N38) );
  NAND3_X1 U7477 ( .A1(\mult_19/SUMB[31][5] ), .A2(n1266), .A3(
        \mult_19/CARRYB[31][4] ), .ZN(n1256) );
  XOR2_X1 U7478 ( .A(\mult_19/CARRYB[31][5] ), .B(\mult_19/SUMB[31][6] ), .Z(
        n1266) );
  NAND3_X1 U7479 ( .A1(\mult_19/SUMB[31][4] ), .A2(n1272), .A3(
        \mult_19/CARRYB[31][3] ), .ZN(n1268) );
  XOR2_X1 U7480 ( .A(\mult_19/CARRYB[31][4] ), .B(\mult_19/SUMB[31][5] ), .Z(
        n1272) );
  NAND3_X1 U7481 ( .A1(\mult_19/SUMB[31][3] ), .A2(n1274), .A3(
        \mult_19/CARRYB[31][2] ), .ZN(n1263) );
  XOR2_X1 U7482 ( .A(\mult_19/CARRYB[31][3] ), .B(\mult_19/SUMB[31][4] ), .Z(
        n1274) );
  XOR2_X1 U7483 ( .A(n1260), .B(n1276), .Z(N34) );
  NAND3_X1 U7484 ( .A1(\mult_19/CARRYB[31][0] ), .A2(n1280), .A3(
        \mult_19/SUMB[31][1] ), .ZN(n1260) );
  XOR2_X1 U7485 ( .A(\mult_19/CARRYB[31][1] ), .B(\mult_19/SUMB[31][2] ), .Z(
        n1280) );
  XOR2_X1 U7486 ( .A(\mult_19/SUMB[31][1] ), .B(\mult_19/CARRYB[31][0] ), .Z(
        N32) );
  XOR2_X1 U7488 ( .A(n2171), .B(n1294), .Z(N253) );
  XOR2_X1 U7490 ( .A(\mult_22/CARRYB[63][60] ), .B(\mult_22/SUMB[63][61] ), 
        .Z(n1299) );
  XOR2_X1 U7492 ( .A(\mult_22/CARRYB[63][59] ), .B(\mult_22/SUMB[63][60] ), 
        .Z(n1307) );
  XOR2_X1 U7494 ( .A(\mult_22/CARRYB[63][58] ), .B(\mult_22/SUMB[63][59] ), 
        .Z(n1310) );
  XOR2_X1 U7495 ( .A(n2064), .B(n1315), .Z(N249) );
  XOR2_X1 U7497 ( .A(\mult_22/CARRYB[63][56] ), .B(\mult_22/SUMB[63][57] ), 
        .Z(n1320) );
  NAND3_X1 U7499 ( .A1(\mult_22/CARRYB[63][54] ), .A2(n1328), .A3(
        \mult_22/SUMB[63][55] ), .ZN(n1323) );
  XOR2_X1 U7500 ( .A(\mult_22/CARRYB[63][55] ), .B(\mult_22/SUMB[63][56] ), 
        .Z(n1328) );
  XOR2_X1 U7502 ( .A(\mult_22/CARRYB[63][54] ), .B(\mult_22/SUMB[63][55] ), 
        .Z(n1330) );
  NAND3_X1 U7504 ( .A1(\mult_22/CARRYB[63][52] ), .A2(n1338), .A3(
        \mult_22/SUMB[63][53] ), .ZN(n1333) );
  XOR2_X1 U7505 ( .A(\mult_22/CARRYB[63][53] ), .B(\mult_22/SUMB[63][54] ), 
        .Z(n1338) );
  XOR2_X1 U7506 ( .A(n2179), .B(n1339), .Z(N244) );
  XOR2_X1 U7507 ( .A(\mult_22/CARRYB[63][52] ), .B(\mult_22/SUMB[63][53] ), 
        .Z(n1340) );
  XOR2_X1 U7508 ( .A(n1802), .B(n1344), .Z(N243) );
  NAND3_X1 U7509 ( .A1(\mult_22/CARRYB[63][50] ), .A2(n1348), .A3(
        \mult_22/SUMB[63][51] ), .ZN(n1343) );
  XOR2_X1 U7510 ( .A(\mult_22/CARRYB[63][51] ), .B(\mult_22/SUMB[63][52] ), 
        .Z(n1348) );
  XOR2_X1 U7511 ( .A(n2107), .B(n1349), .Z(N242) );
  XOR2_X1 U7512 ( .A(\mult_22/CARRYB[63][50] ), .B(\mult_22/SUMB[63][51] ), 
        .Z(n1350) );
  XOR2_X1 U7513 ( .A(n1354), .B(n2056), .Z(N241) );
  NAND3_X1 U7514 ( .A1(\mult_22/CARRYB[63][48] ), .A2(n1358), .A3(
        \mult_22/SUMB[63][49] ), .ZN(n1353) );
  XOR2_X1 U7515 ( .A(\mult_22/CARRYB[63][49] ), .B(\mult_22/SUMB[63][50] ), 
        .Z(n1358) );
  XOR2_X1 U7516 ( .A(n2085), .B(n1359), .Z(N240) );
  XOR2_X1 U7517 ( .A(\mult_22/CARRYB[63][48] ), .B(\mult_22/SUMB[63][49] ), 
        .Z(n1360) );
  XOR2_X1 U7518 ( .A(n1364), .B(n2172), .Z(N239) );
  NAND3_X1 U7519 ( .A1(\mult_22/CARRYB[63][46] ), .A2(n1368), .A3(
        \mult_22/SUMB[63][47] ), .ZN(n1363) );
  XOR2_X1 U7520 ( .A(\mult_22/CARRYB[63][47] ), .B(\mult_22/SUMB[63][48] ), 
        .Z(n1368) );
  XOR2_X1 U7521 ( .A(n2181), .B(n1369), .Z(N238) );
  XOR2_X1 U7522 ( .A(\mult_22/CARRYB[63][46] ), .B(\mult_22/SUMB[63][47] ), 
        .Z(n1370) );
  NAND3_X1 U7523 ( .A1(n630), .A2(n628), .A3(n629), .ZN(n1373) );
  XOR2_X1 U7524 ( .A(n1382), .B(n1383), .Z(N237) );
  NAND3_X1 U7525 ( .A1(\mult_22/CARRYB[63][44] ), .A2(n1386), .A3(
        \mult_22/SUMB[63][45] ), .ZN(n1375) );
  XOR2_X1 U7526 ( .A(\mult_22/CARRYB[63][45] ), .B(\mult_22/SUMB[63][46] ), 
        .Z(n1386) );
  XOR2_X1 U7527 ( .A(n1384), .B(n1387), .Z(N236) );
  XOR2_X1 U7528 ( .A(\mult_22/CARRYB[63][44] ), .B(\mult_22/SUMB[63][45] ), 
        .Z(n1388) );
  XOR2_X1 U7529 ( .A(n1390), .B(n1389), .Z(N235) );
  NAND3_X1 U7530 ( .A1(\mult_22/CARRYB[63][42] ), .A2(n1392), .A3(
        \mult_22/SUMB[63][43] ), .ZN(n1381) );
  XOR2_X1 U7531 ( .A(\mult_22/CARRYB[63][43] ), .B(\mult_22/SUMB[63][44] ), 
        .Z(n1392) );
  XOR2_X1 U7532 ( .A(n2232), .B(n1393), .Z(N234) );
  NAND3_X1 U7533 ( .A1(\mult_22/CARRYB[63][41] ), .A2(n1394), .A3(
        \mult_22/SUMB[63][42] ), .ZN(n1380) );
  XOR2_X1 U7534 ( .A(\mult_22/CARRYB[63][42] ), .B(\mult_22/SUMB[63][43] ), 
        .Z(n1394) );
  XOR2_X1 U7536 ( .A(n1405), .B(n1406), .Z(N233) );
  NAND3_X1 U7537 ( .A1(\mult_22/CARRYB[63][40] ), .A2(n1409), .A3(
        \mult_22/SUMB[63][41] ), .ZN(n1397) );
  XOR2_X1 U7538 ( .A(\mult_22/CARRYB[63][41] ), .B(\mult_22/SUMB[63][42] ), 
        .Z(n1409) );
  XOR2_X1 U7539 ( .A(n1407), .B(n1410), .Z(N232) );
  XOR2_X1 U7540 ( .A(\mult_22/CARRYB[63][40] ), .B(\mult_22/SUMB[63][41] ), 
        .Z(n1411) );
  XOR2_X1 U7541 ( .A(n1413), .B(n1412), .Z(N231) );
  NAND3_X1 U7542 ( .A1(\mult_22/CARRYB[63][38] ), .A2(n1415), .A3(
        \mult_22/SUMB[63][39] ), .ZN(n1403) );
  XOR2_X1 U7543 ( .A(\mult_22/CARRYB[63][39] ), .B(\mult_22/SUMB[63][40] ), 
        .Z(n1415) );
  XOR2_X1 U7544 ( .A(n2378), .B(n1416), .Z(N230) );
  NAND3_X1 U7545 ( .A1(\mult_22/CARRYB[63][37] ), .A2(n1417), .A3(
        \mult_22/SUMB[63][38] ), .ZN(n1401) );
  XOR2_X1 U7546 ( .A(\mult_22/CARRYB[63][38] ), .B(\mult_22/SUMB[63][39] ), 
        .Z(n1417) );
  NAND3_X1 U7547 ( .A1(\mult_22/CARRYB[63][36] ), .A2(n1429), .A3(
        \mult_22/SUMB[63][37] ), .ZN(n1421) );
  XOR2_X1 U7548 ( .A(\mult_22/CARRYB[63][37] ), .B(\mult_22/SUMB[63][38] ), 
        .Z(n1429) );
  NAND3_X1 U7549 ( .A1(\mult_22/SUMB[63][36] ), .A2(n1434), .A3(
        \mult_22/CARRYB[63][35] ), .ZN(n1431) );
  XOR2_X1 U7550 ( .A(\mult_22/CARRYB[63][36] ), .B(\mult_22/SUMB[63][37] ), 
        .Z(n1434) );
  NAND3_X1 U7551 ( .A1(\mult_22/CARRYB[63][34] ), .A2(n1437), .A3(
        \mult_22/SUMB[63][35] ), .ZN(n1426) );
  XOR2_X1 U7552 ( .A(\mult_22/CARRYB[63][35] ), .B(\mult_22/SUMB[63][36] ), 
        .Z(n1437) );
  XOR2_X1 U7553 ( .A(n2089), .B(n1440), .Z(N226) );
  NAND3_X1 U7554 ( .A1(\mult_22/SUMB[63][34] ), .A2(n1441), .A3(
        \mult_22/CARRYB[63][33] ), .ZN(n1425) );
  XOR2_X1 U7555 ( .A(\mult_22/CARRYB[63][34] ), .B(\mult_22/SUMB[63][35] ), 
        .Z(n1441) );
  XOR2_X1 U7556 ( .A(n2077), .B(n1445), .Z(N225) );
  NAND3_X1 U7557 ( .A1(\mult_22/CARRYB[63][32] ), .A2(n1449), .A3(
        \mult_22/SUMB[63][33] ), .ZN(n1444) );
  XOR2_X1 U7558 ( .A(\mult_22/CARRYB[63][33] ), .B(\mult_22/SUMB[63][34] ), 
        .Z(n1449) );
  XOR2_X1 U7559 ( .A(n2336), .B(n1450), .Z(N224) );
  XOR2_X1 U7560 ( .A(\mult_22/CARRYB[63][32] ), .B(\mult_22/SUMB[63][33] ), 
        .Z(n1451) );
  XOR2_X1 U7561 ( .A(n2132), .B(n1455), .Z(N223) );
  NAND3_X1 U7562 ( .A1(\mult_22/CARRYB[63][30] ), .A2(n1459), .A3(
        \mult_22/SUMB[63][31] ), .ZN(n1454) );
  XOR2_X1 U7563 ( .A(\mult_22/CARRYB[63][31] ), .B(\mult_22/SUMB[63][32] ), 
        .Z(n1459) );
  XOR2_X1 U7564 ( .A(n2106), .B(n1460), .Z(N222) );
  XOR2_X1 U7565 ( .A(\mult_22/CARRYB[63][30] ), .B(\mult_22/SUMB[63][31] ), 
        .Z(n1461) );
  XOR2_X1 U7567 ( .A(n1473), .B(n1474), .Z(N221) );
  XOR2_X1 U7568 ( .A(n1475), .B(n1477), .Z(N220) );
  XOR2_X1 U7569 ( .A(\mult_22/CARRYB[63][28] ), .B(\mult_22/SUMB[63][29] ), 
        .Z(n1478) );
  XOR2_X1 U7570 ( .A(n1481), .B(n1480), .Z(N219) );
  XOR2_X1 U7571 ( .A(\mult_22/CARRYB[63][27] ), .B(\mult_22/SUMB[63][28] ), 
        .Z(n1483) );
  XOR2_X1 U7572 ( .A(n2365), .B(n1485), .Z(N218) );
  NAND3_X1 U7573 ( .A1(\mult_22/CARRYB[63][25] ), .A2(n1486), .A3(
        \mult_22/SUMB[63][26] ), .ZN(n1468) );
  XOR2_X1 U7574 ( .A(\mult_22/CARRYB[63][26] ), .B(\mult_22/SUMB[63][27] ), 
        .Z(n1486) );
  XOR2_X1 U7576 ( .A(n1499), .B(n1500), .Z(N217) );
  NAND3_X1 U7577 ( .A1(\mult_22/CARRYB[63][24] ), .A2(n1502), .A3(
        \mult_22/SUMB[63][25] ), .ZN(n1489) );
  XOR2_X1 U7578 ( .A(\mult_22/CARRYB[63][25] ), .B(\mult_22/SUMB[63][26] ), 
        .Z(n1502) );
  XOR2_X1 U7579 ( .A(n1501), .B(n1503), .Z(N216) );
  XOR2_X1 U7580 ( .A(\mult_22/CARRYB[63][24] ), .B(\mult_22/SUMB[63][25] ), 
        .Z(n1504) );
  XOR2_X1 U7581 ( .A(n1506), .B(n1505), .Z(N215) );
  NAND3_X1 U7582 ( .A1(\mult_22/CARRYB[63][22] ), .A2(n1508), .A3(
        \mult_22/SUMB[63][23] ), .ZN(n1497) );
  XOR2_X1 U7583 ( .A(\mult_22/CARRYB[63][23] ), .B(\mult_22/SUMB[63][24] ), 
        .Z(n1508) );
  XOR2_X1 U7584 ( .A(n1491), .B(n1509), .Z(N214) );
  XOR2_X1 U7586 ( .A(n1526), .B(n1527), .Z(N213) );
  XOR2_X1 U7587 ( .A(n1528), .B(n1529), .Z(N212) );
  XOR2_X1 U7588 ( .A(\mult_22/CARRYB[63][20] ), .B(\mult_22/SUMB[63][21] ), 
        .Z(n1530) );
  XOR2_X1 U7589 ( .A(n1533), .B(n1532), .Z(N211) );
  XOR2_X1 U7590 ( .A(\mult_22/CARRYB[63][19] ), .B(\mult_22/SUMB[63][20] ), 
        .Z(n1534) );
  XOR2_X1 U7591 ( .A(n2182), .B(n1536), .Z(N210) );
  NAND3_X1 U7592 ( .A1(\mult_22/CARRYB[63][17] ), .A2(n1537), .A3(
        \mult_22/SUMB[63][18] ), .ZN(n1524) );
  XOR2_X1 U7593 ( .A(\mult_22/CARRYB[63][18] ), .B(\mult_22/SUMB[63][19] ), 
        .Z(n1537) );
  XOR2_X1 U7594 ( .A(n1541), .B(n2173), .Z(N209) );
  NAND3_X1 U7595 ( .A1(\mult_22/CARRYB[63][16] ), .A2(n1545), .A3(
        \mult_22/SUMB[63][17] ), .ZN(n1540) );
  XOR2_X1 U7596 ( .A(\mult_22/CARRYB[63][17] ), .B(\mult_22/SUMB[63][18] ), 
        .Z(n1545) );
  XOR2_X1 U7597 ( .A(n2175), .B(n1546), .Z(N208) );
  XOR2_X1 U7598 ( .A(\mult_22/CARRYB[63][16] ), .B(\mult_22/SUMB[63][17] ), 
        .Z(n1547) );
  XOR2_X1 U7599 ( .A(n2084), .B(n1551), .Z(N207) );
  NAND3_X1 U7600 ( .A1(\mult_22/CARRYB[63][14] ), .A2(n1555), .A3(
        \mult_22/SUMB[63][15] ), .ZN(n1550) );
  XOR2_X1 U7601 ( .A(\mult_22/CARRYB[63][15] ), .B(\mult_22/SUMB[63][16] ), 
        .Z(n1555) );
  XOR2_X1 U7602 ( .A(n2082), .B(n1556), .Z(N206) );
  XOR2_X1 U7603 ( .A(\mult_22/CARRYB[63][14] ), .B(\mult_22/SUMB[63][15] ), 
        .Z(n1557) );
  XOR2_X1 U7605 ( .A(n1569), .B(n1570), .Z(N205) );
  XOR2_X1 U7606 ( .A(n1571), .B(n1573), .Z(N204) );
  XOR2_X1 U7607 ( .A(\mult_22/CARRYB[63][12] ), .B(\mult_22/SUMB[63][13] ), 
        .Z(n1574) );
  XOR2_X1 U7608 ( .A(n1577), .B(n1576), .Z(N203) );
  XOR2_X1 U7609 ( .A(\mult_22/CARRYB[63][11] ), .B(\mult_22/SUMB[63][12] ), 
        .Z(n1579) );
  XOR2_X1 U7610 ( .A(n2341), .B(n1581), .Z(N202) );
  NAND3_X1 U7611 ( .A1(\mult_22/CARRYB[63][9] ), .A2(n1582), .A3(
        \mult_22/SUMB[63][10] ), .ZN(n1564) );
  XOR2_X1 U7612 ( .A(\mult_22/CARRYB[63][10] ), .B(\mult_22/SUMB[63][11] ), 
        .Z(n1582) );
  NAND3_X1 U7614 ( .A1(\mult_22/CARRYB[63][8] ), .A2(n1597), .A3(
        \mult_22/SUMB[63][9] ), .ZN(n1585) );
  XOR2_X1 U7615 ( .A(\mult_22/CARRYB[63][9] ), .B(\mult_22/SUMB[63][10] ), .Z(
        n1597) );
  XOR2_X1 U7616 ( .A(n1598), .B(n1599), .Z(N200) );
  XOR2_X1 U7617 ( .A(\mult_22/CARRYB[63][8] ), .B(\mult_22/SUMB[63][9] ), .Z(
        n1600) );
  NAND3_X1 U7618 ( .A1(\mult_22/CARRYB[63][6] ), .A2(n1603), .A3(
        \mult_22/SUMB[63][7] ), .ZN(n1593) );
  XOR2_X1 U7619 ( .A(\mult_22/CARRYB[63][7] ), .B(\mult_22/SUMB[63][8] ), .Z(
        n1603) );
  XOR2_X1 U7620 ( .A(n2366), .B(n1605), .Z(N198) );
  XOR2_X1 U7621 ( .A(n1620), .B(n1621), .Z(N197) );
  XOR2_X1 U7622 ( .A(n1624), .B(n1623), .Z(N196) );
  XOR2_X1 U7623 ( .A(\mult_22/CARRYB[63][4] ), .B(\mult_22/SUMB[63][5] ), .Z(
        n1626) );
  XOR2_X1 U7624 ( .A(n1613), .B(n1631), .Z(N194) );
  NAND3_X1 U7625 ( .A1(n2354), .A2(\mult_22/CARRYB[63][1] ), .A3(
        \mult_22/SUMB[63][2] ), .ZN(n1618) );
  XOR2_X1 U7626 ( .A(n1632), .B(n1633), .Z(N193) );
  XOR2_X1 U7627 ( .A(\mult_22/CARRYB[63][1] ), .B(\mult_22/SUMB[63][2] ), .Z(
        n1633) );
  XOR2_X1 U7628 ( .A(\mult_22/SUMB[63][1] ), .B(\mult_22/CARRYB[63][0] ), .Z(
        N192) );
  XOR2_X1 U7629 ( .A(n907), .B(n1634), .Z(N129) );
  XOR2_X1 U7630 ( .A(n1639), .B(n1635), .Z(N126) );
  NAND3_X1 U7631 ( .A1(\mult_20/SUMB[31][30] ), .A2(n394), .A3(
        \mult_20/CARRYB[31][29] ), .ZN(n1638) );
  XOR2_X1 U7632 ( .A(n1637), .B(\mult_20/CARRYB[31][30] ), .Z(n1636) );
  XOR2_X1 U7633 ( .A(n1651), .B(n1647), .Z(N124) );
  NAND3_X1 U7634 ( .A1(\mult_20/SUMB[31][28] ), .A2(n1650), .A3(
        \mult_20/CARRYB[31][27] ), .ZN(n1649) );
  XOR2_X1 U7635 ( .A(\mult_20/CARRYB[31][28] ), .B(\mult_20/SUMB[31][29] ), 
        .Z(n1650) );
  XOR2_X1 U7636 ( .A(n1663), .B(n1659), .Z(N122) );
  NAND3_X1 U7637 ( .A1(\mult_20/SUMB[31][26] ), .A2(n1662), .A3(
        \mult_20/CARRYB[31][25] ), .ZN(n1661) );
  XOR2_X1 U7638 ( .A(\mult_20/CARRYB[31][26] ), .B(\mult_20/SUMB[31][27] ), 
        .Z(n1662) );
  XOR2_X1 U7639 ( .A(n1675), .B(n1671), .Z(N120) );
  NAND3_X1 U7640 ( .A1(\mult_20/SUMB[31][24] ), .A2(n1674), .A3(
        \mult_20/CARRYB[31][23] ), .ZN(n1673) );
  XOR2_X1 U7641 ( .A(\mult_20/CARRYB[31][24] ), .B(\mult_20/SUMB[31][25] ), 
        .Z(n1674) );
  XOR2_X1 U7642 ( .A(n1677), .B(n1682), .Z(N119) );
  NAND3_X1 U7643 ( .A1(\mult_20/SUMB[31][22] ), .A2(n1687), .A3(
        \mult_20/CARRYB[31][21] ), .ZN(n1685) );
  XOR2_X1 U7644 ( .A(\mult_20/CARRYB[31][22] ), .B(\mult_20/SUMB[31][23] ), 
        .Z(n1687) );
  XOR2_X1 U7645 ( .A(n1689), .B(n1693), .Z(N117) );
  XOR2_X1 U7646 ( .A(n1696), .B(n1697), .Z(N116) );
  NAND3_X1 U7647 ( .A1(\mult_20/SUMB[31][20] ), .A2(n1698), .A3(
        \mult_20/CARRYB[31][19] ), .ZN(n1695) );
  XOR2_X1 U7648 ( .A(\mult_20/CARRYB[31][20] ), .B(\mult_20/SUMB[31][21] ), 
        .Z(n1698) );
  XOR2_X1 U7649 ( .A(n1704), .B(n1700), .Z(N115) );
  XOR2_X1 U7650 ( .A(\mult_20/CARRYB[31][19] ), .B(\mult_20/SUMB[31][20] ), 
        .Z(n1703) );
  XOR2_X1 U7651 ( .A(n1705), .B(n1708), .Z(N114) );
  XOR2_X1 U7652 ( .A(\mult_20/CARRYB[31][18] ), .B(\mult_20/SUMB[31][19] ), 
        .Z(n1709) );
  XOR2_X1 U7653 ( .A(n1713), .B(n1710), .Z(N113) );
  NAND3_X1 U7654 ( .A1(\mult_20/SUMB[31][17] ), .A2(n1717), .A3(
        \mult_20/CARRYB[31][16] ), .ZN(n1712) );
  XOR2_X1 U7655 ( .A(\mult_20/CARRYB[31][17] ), .B(\mult_20/SUMB[31][18] ), 
        .Z(n1717) );
  XOR2_X1 U7656 ( .A(n1714), .B(n1718), .Z(N112) );
  XOR2_X1 U7657 ( .A(\mult_20/CARRYB[31][16] ), .B(\mult_20/SUMB[31][17] ), 
        .Z(n1719) );
  XOR2_X1 U7658 ( .A(\mult_20/CARRYB[31][15] ), .B(\mult_20/SUMB[31][16] ), 
        .Z(n1725) );
  XOR2_X1 U7659 ( .A(n1726), .B(n1729), .Z(N110) );
  XOR2_X1 U7660 ( .A(\mult_20/CARRYB[31][14] ), .B(\mult_20/SUMB[31][15] ), 
        .Z(n1730) );
  NAND3_X1 U7661 ( .A1(n408), .A2(n1739), .A3(n1740), .ZN(n1737) );
  XOR2_X1 U7662 ( .A(n1741), .B(n1742), .Z(N109) );
  NAND3_X1 U7663 ( .A1(\mult_20/CARRYB[31][12] ), .A2(n1745), .A3(
        \mult_20/SUMB[31][13] ), .ZN(n1733) );
  XOR2_X1 U7664 ( .A(\mult_20/CARRYB[31][13] ), .B(\mult_20/SUMB[31][14] ), 
        .Z(n1745) );
  XOR2_X1 U7665 ( .A(n1743), .B(n1746), .Z(N108) );
  XOR2_X1 U7666 ( .A(\mult_20/CARRYB[31][12] ), .B(\mult_20/SUMB[31][13] ), 
        .Z(n1747) );
  XOR2_X1 U7667 ( .A(n1749), .B(n1748), .Z(N107) );
  NAND3_X1 U7668 ( .A1(\mult_20/CARRYB[31][10] ), .A2(n1751), .A3(
        \mult_20/SUMB[31][11] ), .ZN(n1738) );
  XOR2_X1 U7669 ( .A(\mult_20/CARRYB[31][11] ), .B(\mult_20/SUMB[31][12] ), 
        .Z(n1751) );
  NAND3_X1 U7671 ( .A1(n1759), .A2(n1760), .A3(n1761), .ZN(n1758) );
  XOR2_X1 U7672 ( .A(n1768), .B(n1769), .Z(N105) );
  XOR2_X1 U7673 ( .A(n1770), .B(n1771), .Z(N104) );
  XOR2_X1 U7674 ( .A(\mult_20/CARRYB[31][8] ), .B(\mult_20/SUMB[31][9] ), .Z(
        n1772) );
  XOR2_X1 U7675 ( .A(n1774), .B(n1773), .Z(N103) );
  NAND3_X1 U7676 ( .A1(\mult_20/CARRYB[31][6] ), .A2(n1776), .A3(
        \mult_20/SUMB[31][7] ), .ZN(n1766) );
  XOR2_X1 U7677 ( .A(\mult_20/CARRYB[31][7] ), .B(\mult_20/SUMB[31][8] ), .Z(
        n1776) );
  XOR2_X1 U7678 ( .A(n1759), .B(n1777), .Z(N102) );
  XOR2_X1 U7679 ( .A(n1789), .B(n1790), .Z(N101) );
  NAND3_X1 U7680 ( .A1(\mult_20/SUMB[31][5] ), .A2(n1791), .A3(
        \mult_20/CARRYB[31][4] ), .ZN(n1782) );
  XOR2_X1 U7681 ( .A(\mult_20/CARRYB[31][5] ), .B(\mult_20/SUMB[31][6] ), .Z(
        n1791) );
  XOR2_X1 U7682 ( .A(n1794), .B(n1793), .Z(N100) );
  NAND3_X1 U7683 ( .A1(\mult_20/SUMB[31][3] ), .A2(n1795), .A3(
        \mult_20/CARRYB[31][2] ), .ZN(n1788) );
  NAND3_X1 U7684 ( .A1(\mult_20/CARRYB[31][0] ), .A2(n1107), .A3(
        \mult_20/SUMB[31][1] ), .ZN(n1103) );
  XOR2_X1 U7685 ( .A(\mult_20/CARRYB[31][1] ), .B(\mult_20/SUMB[31][2] ), .Z(
        n1107) );
  XOR2_X1 U7686 ( .A(\mult_20/CARRYB[31][2] ), .B(\mult_20/SUMB[31][3] ), .Z(
        n1797) );
  XOR2_X1 U7687 ( .A(\mult_20/CARRYB[31][3] ), .B(\mult_20/SUMB[31][4] ), .Z(
        n1795) );
  NAND3_X1 U7688 ( .A1(\mult_20/SUMB[31][4] ), .A2(n1798), .A3(
        \mult_20/CARRYB[31][3] ), .ZN(n1787) );
  XOR2_X1 U7689 ( .A(\mult_20/CARRYB[31][4] ), .B(\mult_20/SUMB[31][5] ), .Z(
        n1798) );
  XOR2_X1 U7690 ( .A(n1099), .B(n1799), .Z(N1) );
  FA_X1 \mult_22/S0_55  ( .A(\mult_22/ab[1][55] ), .B(1'b0), .CI(
        \mult_22/ab[0][56] ), .CO(\mult_22/CARRYB[1][55] ), .S(
        \mult_22/SUMB[1][55] ) );
  DFF_X1 \reg_mid_0_reg[0]  ( .D(N0), .CK(g_inClk), .Q(reg_mid_0[0]), .QN(
        n2377) );
  DFF_X1 \reg_mid_0_reg[1]  ( .D(N1), .CK(g_inClk), .Q(reg_mid_0[1]), .QN(
        n2373) );
  DFF_X2 \reg_out_reg[127]  ( .D(N255), .CK(g_inClk), .Q(g_outM[127]) );
  DFF_X2 \reg_out_reg[125]  ( .D(N253), .CK(g_inClk), .Q(g_outM[125]) );
  DFF_X2 \reg_out_reg[123]  ( .D(N251), .CK(g_inClk), .Q(g_outM[123]) );
  DFF_X2 \reg_out_reg[121]  ( .D(N249), .CK(g_inClk), .Q(g_outM[121]) );
  DFF_X2 \reg_out_reg[119]  ( .D(N247), .CK(g_inClk), .Q(g_outM[119]) );
  DFF_X2 \reg_out_reg[117]  ( .D(N245), .CK(g_inClk), .Q(g_outM[117]) );
  BUF_X1 U7691 ( .A(n2174), .Z(n1802) );
  AND2_X1 U7692 ( .A1(n1518), .A2(n1517), .ZN(n1803) );
  CLKBUF_X1 U7693 ( .A(n1283), .Z(n1804) );
  CLKBUF_X1 U7694 ( .A(n746), .Z(n2742) );
  NOR2_X1 U7695 ( .A1(n2737), .A2(n2770), .ZN(\mult_22/ab[5][61] ) );
  NOR2_X1 U7696 ( .A1(n2684), .A2(n2769), .ZN(\mult_22/ab[5][51] ) );
  NOR2_X1 U7697 ( .A1(n2658), .A2(n2835), .ZN(\mult_22/ab[16][46] ) );
  NOR2_X1 U7698 ( .A1(n2664), .A2(n2823), .ZN(\mult_22/ab[14][47] ) );
  NOR2_X1 U7699 ( .A1(n2616), .A2(n2852), .ZN(\mult_22/ab[19][39] ) );
  NOR2_X1 U7700 ( .A1(n2557), .A2(n2929), .ZN(\mult_22/ab[32][29] ) );
  BUF_X2 U7701 ( .A(n2111), .Z(n2751) );
  INV_X1 U7702 ( .A(\mult_22/ab[32][29] ), .ZN(n2213) );
  BUF_X1 U7703 ( .A(n1852), .Z(n2852) );
  BUF_X2 U7704 ( .A(n1853), .Z(n2398) );
  CLKBUF_X1 U7705 ( .A(n746), .Z(n2744) );
  AOI21_X1 U7706 ( .B1(\mult_22/CARRYB[63][42] ), .B2(\mult_22/SUMB[63][43] ), 
        .A(n1392), .ZN(n1379) );
  AND2_X1 U7707 ( .A1(\mult_22/SUMB[63][1] ), .A2(\mult_22/CARRYB[63][0] ), 
        .ZN(n1632) );
  AOI21_X1 U7708 ( .B1(\mult_22/CARRYB[63][7] ), .B2(\mult_22/SUMB[63][8] ), 
        .A(n1600), .ZN(n1589) );
  NOR2_X1 U7709 ( .A1(n1574), .A2(n1575), .ZN(n1572) );
  AOI21_X1 U7710 ( .B1(\mult_22/CARRYB[63][17] ), .B2(\mult_22/SUMB[63][18] ), 
        .A(n1537), .ZN(n1520) );
  NOR2_X1 U7711 ( .A1(n1478), .A2(n1479), .ZN(n1476) );
  AOI21_X1 U7712 ( .B1(\mult_22/SUMB[63][34] ), .B2(\mult_22/CARRYB[63][33] ), 
        .A(n1441), .ZN(n1438) );
  BUF_X1 U7713 ( .A(n751), .Z(n2717) );
  BUF_X1 U7714 ( .A(n751), .Z(n2718) );
  BUF_X1 U7715 ( .A(n752), .Z(n2714) );
  BUF_X2 U7716 ( .A(n3512), .Z(n3511) );
  AND2_X1 U7717 ( .A1(n1588), .A2(n583), .ZN(n1830) );
  AND2_X1 U7718 ( .A1(n582), .A2(n580), .ZN(n1831) );
  AND2_X1 U7719 ( .A1(n1492), .A2(n600), .ZN(n1879) );
  AND2_X1 U7720 ( .A1(n2337), .A2(n2338), .ZN(n1880) );
  BUF_X1 U7721 ( .A(n752), .Z(n2713) );
  INV_X1 U7722 ( .A(reg_mid_1[57]), .ZN(n751) );
  AND2_X1 U7723 ( .A1(n617), .A2(n619), .ZN(n1884) );
  AND3_X1 U7724 ( .A1(n613), .A2(n615), .A3(n616), .ZN(n1885) );
  XNOR2_X1 U7725 ( .A(n2057), .B(n2052), .ZN(N245) );
  AND2_X1 U7726 ( .A1(n639), .A2(n1333), .ZN(n2052) );
  XNOR2_X1 U7727 ( .A(n2060), .B(n2053), .ZN(N247) );
  AND2_X1 U7728 ( .A1(n641), .A2(n1323), .ZN(n2053) );
  XNOR2_X1 U7729 ( .A(n2321), .B(n2055), .ZN(N246) );
  OR2_X1 U7730 ( .A1(n1326), .A2(n1327), .ZN(n2055) );
  AOI21_X1 U7731 ( .B1(n2085), .B2(n633), .A(n1356), .ZN(n2056) );
  AOI21_X1 U7732 ( .B1(n2179), .B2(n638), .A(n1336), .ZN(n2057) );
  XNOR2_X1 U7733 ( .A(n2176), .B(n2058), .ZN(N248) );
  OR2_X1 U7734 ( .A1(n1317), .A2(n1318), .ZN(n2058) );
  AOI21_X1 U7735 ( .B1(n2128), .B2(n640), .A(n1326), .ZN(n2060) );
  XNOR2_X1 U7736 ( .A(n2342), .B(n2061), .ZN(N250) );
  OR2_X1 U7737 ( .A1(n1305), .A2(n1306), .ZN(n2061) );
  AOI21_X1 U7738 ( .B1(n2128), .B2(n640), .A(n1326), .ZN(n2160) );
  XNOR2_X1 U7739 ( .A(n2068), .B(n2062), .ZN(N251) );
  AND2_X1 U7740 ( .A1(n1302), .A2(n645), .ZN(n2062) );
  AOI21_X1 U7741 ( .B1(n2176), .B2(n642), .A(n1317), .ZN(n2064) );
  XNOR2_X1 U7742 ( .A(n2170), .B(n2065), .ZN(N252) );
  OR2_X1 U7743 ( .A1(n1296), .A2(n1297), .ZN(n2065) );
  XNOR2_X1 U7744 ( .A(n1804), .B(n2066), .ZN(N254) );
  OR2_X1 U7745 ( .A1(n1284), .A2(n1285), .ZN(n2066) );
  AOI21_X1 U7746 ( .B1(n2105), .B2(n644), .A(n1305), .ZN(n2068) );
  OR2_X1 U7747 ( .A1(n2592), .A2(n2894), .ZN(n2069) );
  INV_X1 U7748 ( .A(n2069), .ZN(n2070) );
  XOR2_X1 U7749 ( .A(\mult_22/CARRYB[13][47] ), .B(\mult_22/ab[14][47] ), .Z(
        n2071) );
  XOR2_X1 U7750 ( .A(\mult_22/SUMB[13][48] ), .B(n2071), .Z(
        \mult_22/SUMB[14][47] ) );
  NAND2_X1 U7751 ( .A1(\mult_22/SUMB[13][48] ), .A2(\mult_22/CARRYB[13][47] ), 
        .ZN(n2072) );
  NAND2_X1 U7752 ( .A1(\mult_22/SUMB[13][48] ), .A2(\mult_22/ab[14][47] ), 
        .ZN(n2073) );
  NAND2_X1 U7753 ( .A1(\mult_22/CARRYB[13][47] ), .A2(\mult_22/ab[14][47] ), 
        .ZN(n2074) );
  NAND3_X1 U7754 ( .A1(n2072), .A2(n2073), .A3(n2074), .ZN(
        \mult_22/CARRYB[14][47] ) );
  CLKBUF_X1 U7755 ( .A(n2142), .Z(n3496) );
  BUF_X1 U7756 ( .A(reg_mid_0[1]), .Z(n2188) );
  XNOR2_X1 U7757 ( .A(\mult_22/CARRYB[25][35] ), .B(n2069), .ZN(n2279) );
  OR3_X1 U7758 ( .A1(n1615), .A2(n2298), .A3(n1613), .ZN(n1612) );
  CLKBUF_X1 U7759 ( .A(reg_mid_0[0]), .Z(n2120) );
  CLKBUF_X1 U7760 ( .A(reg_mid_0[0]), .Z(n2293) );
  XNOR2_X1 U7761 ( .A(\mult_22/SUMB[20][37] ), .B(n951), .ZN(
        \mult_22/SUMB[21][36] ) );
  XNOR2_X1 U7762 ( .A(n2075), .B(n945), .ZN(\mult_22/SUMB[24][32] ) );
  AND2_X1 U7763 ( .A1(reg_mid_0[24]), .A2(reg_mid_1[32]), .ZN(n2075) );
  CLKBUF_X1 U7764 ( .A(n1446), .Z(n2076) );
  AOI21_X1 U7765 ( .B1(n2076), .B2(n610), .A(n1447), .ZN(n2077) );
  CLKBUF_X1 U7766 ( .A(n2142), .Z(n3499) );
  BUF_X1 U7767 ( .A(n3496), .Z(n3498) );
  INV_X1 U7768 ( .A(\mult_22/ab[18][46] ), .ZN(n2277) );
  CLKBUF_X3 U7769 ( .A(n1856), .Z(n2557) );
  INV_X1 U7770 ( .A(\mult_22/ab[21][44] ), .ZN(n2108) );
  OAI211_X1 U7771 ( .C1(n1487), .C2(n1488), .A(n1489), .B(n1490), .ZN(n1471)
         );
  AOI21_X1 U7772 ( .B1(n1516), .B2(n2216), .A(n2078), .ZN(n1490) );
  INV_X1 U7773 ( .A(n2214), .ZN(n2078) );
  OAI211_X1 U7774 ( .C1(n1419), .C2(n1418), .A(n1420), .B(n1421), .ZN(n1404)
         );
  OAI22_X1 U7775 ( .A1(n1464), .A2(n605), .B1(n1463), .B2(n1462), .ZN(n1456)
         );
  OAI22_X1 U7776 ( .A1(n1560), .A2(n585), .B1(n1559), .B2(n1558), .ZN(n2086)
         );
  CLKBUF_X1 U7777 ( .A(n1402), .Z(n2079) );
  CLKBUF_X1 U7778 ( .A(n1469), .Z(n2080) );
  OAI221_X1 U7779 ( .B1(n1371), .B2(n1372), .C1(n2095), .C2(n1373), .A(n1375), 
        .ZN(n2181) );
  CLKBUF_X1 U7780 ( .A(n2086), .Z(n2082) );
  AOI21_X1 U7781 ( .B1(n1446), .B2(n610), .A(n1447), .ZN(n2083) );
  AOI21_X1 U7782 ( .B1(n2082), .B2(n586), .A(n1553), .ZN(n2084) );
  CLKBUF_X1 U7783 ( .A(n1355), .Z(n2085) );
  AOI21_X1 U7784 ( .B1(n2086), .B2(n586), .A(n1553), .ZN(n1549) );
  CLKBUF_X1 U7785 ( .A(n1516), .Z(n2087) );
  OAI211_X1 U7786 ( .C1(n1400), .C2(n1401), .A(n2079), .B(n1403), .ZN(n2088)
         );
  CLKBUF_X1 U7787 ( .A(n1439), .Z(n2089) );
  OR2_X1 U7788 ( .A1(n972), .A2(n709), .ZN(n2090) );
  NAND2_X1 U7789 ( .A1(n2090), .A2(n973), .ZN(\mult_22/CARRYB[22][38] ) );
  INV_X1 U7790 ( .A(n2183), .ZN(n972) );
  XNOR2_X1 U7791 ( .A(\mult_22/CARRYB[3][62] ), .B(n2091), .ZN(
        \mult_22/SUMB[4][62] ) );
  XNOR2_X1 U7792 ( .A(\mult_22/ab[3][63] ), .B(\mult_22/ab[4][62] ), .ZN(n2091) );
  XNOR2_X1 U7793 ( .A(\mult_22/CARRYB[25][40] ), .B(\mult_22/ab[26][40] ), 
        .ZN(n2130) );
  OAI211_X1 U7794 ( .C1(n1467), .C2(n1468), .A(n2080), .B(n1470), .ZN(n2092)
         );
  AOI21_X1 U7795 ( .B1(n2088), .B2(n620), .A(n1399), .ZN(n2093) );
  AOI21_X1 U7796 ( .B1(n2092), .B2(n604), .A(n1466), .ZN(n2094) );
  CLKBUF_X1 U7797 ( .A(n1374), .Z(n2095) );
  CLKBUF_X1 U7798 ( .A(n1586), .Z(n2096) );
  XOR2_X1 U7799 ( .A(\mult_22/SUMB[4][62] ), .B(\mult_22/ab[5][61] ), .Z(n2097) );
  XOR2_X1 U7800 ( .A(\mult_22/CARRYB[4][61] ), .B(n2097), .Z(
        \mult_22/SUMB[5][61] ) );
  NAND2_X1 U7801 ( .A1(\mult_22/CARRYB[4][61] ), .A2(\mult_22/SUMB[4][62] ), 
        .ZN(n2098) );
  NAND2_X1 U7802 ( .A1(\mult_22/CARRYB[4][61] ), .A2(\mult_22/ab[5][61] ), 
        .ZN(n2099) );
  NAND2_X1 U7803 ( .A1(\mult_22/SUMB[4][62] ), .A2(\mult_22/ab[5][61] ), .ZN(
        n2100) );
  NAND3_X1 U7804 ( .A1(n2098), .A2(n2099), .A3(n2100), .ZN(
        \mult_22/CARRYB[5][61] ) );
  OR2_X1 U7805 ( .A1(n2158), .A2(n2142), .ZN(n2101) );
  XNOR2_X1 U7806 ( .A(\mult_22/CARRYB[3][61] ), .B(n2102), .ZN(
        \mult_22/SUMB[4][61] ) );
  XNOR2_X1 U7807 ( .A(\mult_22/SUMB[3][62] ), .B(\mult_22/ab[4][61] ), .ZN(
        n2102) );
  XNOR2_X1 U7808 ( .A(n2103), .B(\mult_22/SUMB[18][42] ), .ZN(
        \mult_22/SUMB[19][41] ) );
  XNOR2_X1 U7809 ( .A(\mult_22/ab[19][41] ), .B(\mult_22/CARRYB[18][41] ), 
        .ZN(n2103) );
  AOI21_X1 U7810 ( .B1(n2085), .B2(n633), .A(n1356), .ZN(n2104) );
  CLKBUF_X1 U7811 ( .A(n1304), .Z(n2105) );
  AOI21_X1 U7812 ( .B1(n1355), .B2(n633), .A(n1356), .ZN(n1352) );
  OAI22_X1 U7813 ( .A1(n1462), .A2(n1463), .B1(n2094), .B2(n605), .ZN(n2106)
         );
  OAI21_X1 U7814 ( .B1(n2104), .B2(n1351), .A(n1353), .ZN(n2107) );
  BUF_X2 U7815 ( .A(reg_mid_0[1]), .Z(n2189) );
  AND2_X1 U7816 ( .A1(n2322), .A2(reg_mid_1[62]), .ZN(n2112) );
  XNOR2_X1 U7817 ( .A(\mult_22/CARRYB[20][44] ), .B(n2108), .ZN(n2123) );
  AND2_X1 U7818 ( .A1(reg_mid_1[61]), .A2(reg_mid_0[2]), .ZN(
        \mult_22/ab[2][61] ) );
  INV_X1 U7819 ( .A(n2357), .ZN(n2295) );
  XNOR2_X1 U7820 ( .A(n931), .B(n2109), .ZN(\mult_22/SUMB[8][50] ) );
  XNOR2_X1 U7821 ( .A(n731), .B(\mult_22/SUMB[7][51] ), .ZN(n2109) );
  XNOR2_X1 U7822 ( .A(n2110), .B(\mult_22/SUMB[18][43] ), .ZN(
        \mult_22/SUMB[19][42] ) );
  XNOR2_X1 U7823 ( .A(\mult_22/ab[19][42] ), .B(\mult_22/CARRYB[18][42] ), 
        .ZN(n2110) );
  XNOR2_X1 U7824 ( .A(n901), .B(n2112), .ZN(\mult_22/n325 ) );
  XOR2_X1 U7825 ( .A(\mult_22/ab[18][43] ), .B(\mult_22/CARRYB[17][43] ), .Z(
        n2113) );
  XOR2_X1 U7826 ( .A(n2113), .B(\mult_22/SUMB[17][44] ), .Z(
        \mult_22/SUMB[18][43] ) );
  NAND2_X1 U7827 ( .A1(\mult_22/ab[18][43] ), .A2(\mult_22/CARRYB[17][43] ), 
        .ZN(n2114) );
  NAND2_X1 U7828 ( .A1(\mult_22/ab[18][43] ), .A2(\mult_22/SUMB[17][44] ), 
        .ZN(n2115) );
  NAND2_X1 U7829 ( .A1(\mult_22/CARRYB[17][43] ), .A2(\mult_22/SUMB[17][44] ), 
        .ZN(n2116) );
  NAND3_X1 U7830 ( .A1(n2114), .A2(n2115), .A3(n2116), .ZN(
        \mult_22/CARRYB[18][43] ) );
  NAND2_X1 U7831 ( .A1(\mult_22/ab[19][42] ), .A2(\mult_22/CARRYB[18][42] ), 
        .ZN(n2117) );
  NAND2_X1 U7832 ( .A1(\mult_22/ab[19][42] ), .A2(\mult_22/SUMB[18][43] ), 
        .ZN(n2118) );
  NAND2_X1 U7833 ( .A1(\mult_22/CARRYB[18][42] ), .A2(\mult_22/SUMB[18][43] ), 
        .ZN(n2119) );
  NAND3_X1 U7834 ( .A1(n2117), .A2(n2118), .A3(n2119), .ZN(
        \mult_22/CARRYB[19][42] ) );
  BUF_X1 U7835 ( .A(reg_mid_0[0]), .Z(n2292) );
  CLKBUF_X1 U7836 ( .A(n1420), .Z(n2121) );
  NAND2_X1 U7837 ( .A1(n1439), .A2(n2122), .ZN(n1420) );
  AND2_X1 U7838 ( .A1(n2379), .A2(n1885), .ZN(n2122) );
  XOR2_X1 U7839 ( .A(\mult_22/SUMB[20][45] ), .B(n2123), .Z(
        \mult_22/SUMB[21][44] ) );
  NAND2_X1 U7840 ( .A1(\mult_22/SUMB[20][45] ), .A2(\mult_22/CARRYB[20][44] ), 
        .ZN(n2124) );
  NAND2_X1 U7841 ( .A1(\mult_22/SUMB[20][45] ), .A2(\mult_22/ab[21][44] ), 
        .ZN(n2125) );
  NAND2_X1 U7842 ( .A1(\mult_22/CARRYB[20][44] ), .A2(\mult_22/ab[21][44] ), 
        .ZN(n2126) );
  NAND3_X1 U7843 ( .A1(n2124), .A2(n2125), .A3(n2126), .ZN(
        \mult_22/CARRYB[21][44] ) );
  AOI21_X1 U7844 ( .B1(n2105), .B2(n644), .A(n1305), .ZN(n2127) );
  AOI21_X1 U7845 ( .B1(n1304), .B2(n644), .A(n1305), .ZN(n1301) );
  CLKBUF_X1 U7846 ( .A(n1325), .Z(n2128) );
  XNOR2_X1 U7847 ( .A(\mult_22/SUMB[15][47] ), .B(n2129), .ZN(
        \mult_22/SUMB[16][46] ) );
  XNOR2_X1 U7848 ( .A(\mult_22/CARRYB[15][46] ), .B(\mult_22/ab[16][46] ), 
        .ZN(n2129) );
  XNOR2_X1 U7849 ( .A(\mult_22/SUMB[25][41] ), .B(n2130), .ZN(
        \mult_22/SUMB[26][40] ) );
  NOR2_X1 U7850 ( .A1(n621), .A2(n2353), .ZN(n2131) );
  AOI21_X1 U7851 ( .B1(n606), .B2(n2106), .A(n1457), .ZN(n2132) );
  BUF_X1 U7852 ( .A(n2377), .Z(n2142) );
  CLKBUF_X3 U7853 ( .A(n1822), .Z(n2720) );
  INV_X1 U7854 ( .A(reg_mid_1[57]), .ZN(n2133) );
  BUF_X4 U7855 ( .A(n751), .Z(n2716) );
  XOR2_X1 U7856 ( .A(\mult_22/CARRYB[8][51] ), .B(\mult_22/ab[9][51] ), .Z(
        n2134) );
  XOR2_X1 U7857 ( .A(\mult_22/SUMB[8][52] ), .B(n2134), .Z(
        \mult_22/SUMB[9][51] ) );
  NAND2_X1 U7858 ( .A1(\mult_22/SUMB[8][52] ), .A2(\mult_22/CARRYB[8][51] ), 
        .ZN(n2135) );
  NAND2_X1 U7859 ( .A1(\mult_22/SUMB[8][52] ), .A2(\mult_22/ab[9][51] ), .ZN(
        n2136) );
  NAND2_X1 U7860 ( .A1(\mult_22/CARRYB[8][51] ), .A2(\mult_22/ab[9][51] ), 
        .ZN(n2137) );
  NAND3_X1 U7861 ( .A1(n2135), .A2(n2136), .A3(n2137), .ZN(
        \mult_22/CARRYB[9][51] ) );
  OR2_X1 U7862 ( .A1(n706), .A2(n946), .ZN(n2138) );
  NAND2_X1 U7863 ( .A1(n2138), .A2(n969), .ZN(\mult_22/CARRYB[23][37] ) );
  BUF_X1 U7864 ( .A(reg_mid_0[1]), .Z(n2187) );
  CLKBUF_X1 U7865 ( .A(n748), .Z(n2732) );
  NOR2_X1 U7866 ( .A1(n903), .A2(n2101), .ZN(\mult_22/n323 ) );
  BUF_X1 U7867 ( .A(n2373), .Z(n2368) );
  INV_X1 U7868 ( .A(n3497), .ZN(n2139) );
  BUF_X2 U7869 ( .A(n2142), .Z(n3497) );
  CLKBUF_X1 U7870 ( .A(n2140), .Z(n2727) );
  NAND2_X1 U7871 ( .A1(reg_mid_1[63]), .A2(n2292), .ZN(n2141) );
  XNOR2_X1 U7872 ( .A(n809), .B(n2143), .ZN(\mult_22/SUMB[1][61] ) );
  AND2_X1 U7873 ( .A1(reg_mid_1[61]), .A2(n2187), .ZN(n2143) );
  OR2_X1 U7874 ( .A1(n2377), .A2(n2193), .ZN(n809) );
  NAND2_X1 U7875 ( .A1(\mult_22/CARRYB[3][62] ), .A2(\mult_22/ab[3][63] ), 
        .ZN(n2144) );
  NAND2_X1 U7876 ( .A1(\mult_22/CARRYB[3][62] ), .A2(\mult_22/ab[4][62] ), 
        .ZN(n2145) );
  NAND2_X1 U7877 ( .A1(\mult_22/ab[3][63] ), .A2(\mult_22/ab[4][62] ), .ZN(
        n2146) );
  NAND3_X1 U7878 ( .A1(n2144), .A2(n2145), .A3(n2146), .ZN(
        \mult_22/CARRYB[4][62] ) );
  INV_X1 U7879 ( .A(reg_mid_0[2]), .ZN(n2147) );
  INV_X1 U7880 ( .A(reg_mid_0[2]), .ZN(n2148) );
  INV_X1 U7881 ( .A(reg_mid_0[2]), .ZN(n2149) );
  INV_X1 U7882 ( .A(reg_mid_0[2]), .ZN(n2150) );
  INV_X1 U7883 ( .A(reg_mid_0[2]), .ZN(n2151) );
  BUF_X1 U7884 ( .A(n2152), .Z(n2153) );
  BUF_X1 U7885 ( .A(n2152), .Z(n2154) );
  BUF_X1 U7886 ( .A(n2152), .Z(n2155) );
  BUF_X1 U7887 ( .A(n2152), .Z(n2156) );
  BUF_X1 U7888 ( .A(n2152), .Z(n2157) );
  FA_X1 U7889 ( .A(\mult_22/ab[63][4] ), .B(\mult_22/CARRYB[62][4] ), .CI(
        \mult_22/SUMB[62][5] ), .S(n2159) );
  AOI21_X1 U7890 ( .B1(n1325), .B2(n640), .A(n1326), .ZN(n1322) );
  XOR2_X1 U7891 ( .A(\mult_22/ab[4][55] ), .B(\mult_22/CARRYB[3][55] ), .Z(
        n2161) );
  XOR2_X1 U7892 ( .A(n2161), .B(\mult_22/SUMB[3][56] ), .Z(
        \mult_22/SUMB[4][55] ) );
  XOR2_X1 U7893 ( .A(\mult_22/ab[5][54] ), .B(\mult_22/CARRYB[4][54] ), .Z(
        n2162) );
  XOR2_X1 U7894 ( .A(n2162), .B(\mult_22/SUMB[4][55] ), .Z(
        \mult_22/SUMB[5][54] ) );
  NAND2_X1 U7895 ( .A1(\mult_22/ab[4][55] ), .A2(\mult_22/CARRYB[3][55] ), 
        .ZN(n2163) );
  NAND2_X1 U7896 ( .A1(\mult_22/ab[4][55] ), .A2(\mult_22/SUMB[3][56] ), .ZN(
        n2164) );
  NAND2_X1 U7897 ( .A1(\mult_22/CARRYB[3][55] ), .A2(\mult_22/SUMB[3][56] ), 
        .ZN(n2165) );
  NAND3_X1 U7898 ( .A1(n2163), .A2(n2164), .A3(n2165), .ZN(
        \mult_22/CARRYB[4][55] ) );
  NAND2_X1 U7899 ( .A1(\mult_22/ab[5][54] ), .A2(\mult_22/CARRYB[4][54] ), 
        .ZN(n2166) );
  NAND2_X1 U7900 ( .A1(\mult_22/ab[5][54] ), .A2(\mult_22/SUMB[4][55] ), .ZN(
        n2167) );
  NAND2_X1 U7901 ( .A1(\mult_22/CARRYB[4][54] ), .A2(\mult_22/SUMB[4][55] ), 
        .ZN(n2168) );
  NAND3_X1 U7902 ( .A1(n2166), .A2(n2167), .A3(n2168), .ZN(
        \mult_22/CARRYB[5][54] ) );
  CLKBUF_X1 U7903 ( .A(n1618), .Z(n2169) );
  OAI21_X1 U7904 ( .B1(n2127), .B2(n1300), .A(n1302), .ZN(n2170) );
  OAI21_X1 U7905 ( .B1(n1301), .B2(n1300), .A(n1302), .ZN(n1295) );
  AOI21_X1 U7906 ( .B1(n2170), .B2(n646), .A(n1296), .ZN(n2171) );
  AOI21_X1 U7907 ( .B1(n2181), .B2(n631), .A(n1366), .ZN(n2172) );
  AOI21_X1 U7908 ( .B1(n2175), .B2(n588), .A(n1543), .ZN(n2173) );
  AOI21_X1 U7909 ( .B1(n2107), .B2(n635), .A(n1346), .ZN(n2174) );
  OAI21_X1 U7910 ( .B1(n2084), .B2(n1548), .A(n1550), .ZN(n2175) );
  OAI21_X1 U7911 ( .B1(n2160), .B2(n1321), .A(n1323), .ZN(n2176) );
  AOI21_X1 U7912 ( .B1(n1345), .B2(n635), .A(n1346), .ZN(n1342) );
  AOI21_X1 U7913 ( .B1(n1542), .B2(n588), .A(n1543), .ZN(n1539) );
  AOI21_X1 U7914 ( .B1(n1398), .B2(n620), .A(n1399), .ZN(n2177) );
  CLKBUF_X1 U7915 ( .A(n2131), .Z(n2178) );
  OAI21_X1 U7916 ( .B1(n2174), .B2(n1341), .A(n1343), .ZN(n2179) );
  AOI21_X1 U7917 ( .B1(n2176), .B2(n642), .A(n1317), .ZN(n2180) );
  OAI21_X1 U7918 ( .B1(n1538), .B2(n2173), .A(n1540), .ZN(n2182) );
  OR2_X2 U7919 ( .A1(n2223), .A2(n712), .ZN(n2183) );
  XNOR2_X1 U7920 ( .A(n2184), .B(\mult_22/SUMB[28][34] ), .ZN(
        \mult_22/SUMB[29][33] ) );
  XNOR2_X1 U7921 ( .A(\mult_22/ab[29][33] ), .B(\mult_22/CARRYB[28][33] ), 
        .ZN(n2184) );
  CLKBUF_X3 U7922 ( .A(n746), .Z(n2185) );
  CLKBUF_X3 U7923 ( .A(n746), .Z(n2186) );
  XNOR2_X1 U7924 ( .A(\mult_22/CARRYB[2][62] ), .B(n2190), .ZN(
        \mult_22/SUMB[3][62] ) );
  XNOR2_X1 U7925 ( .A(\mult_22/ab[2][63] ), .B(\mult_22/ab[3][62] ), .ZN(n2190) );
  NAND3_X1 U7926 ( .A1(n2318), .A2(n2319), .A3(n2320), .ZN(n2191) );
  XNOR2_X1 U7927 ( .A(n903), .B(n2192), .ZN(\mult_22/n196 ) );
  AND2_X1 U7928 ( .A1(reg_mid_0[0]), .A2(reg_mid_1[61]), .ZN(n2192) );
  CLKBUF_X3 U7929 ( .A(n2111), .Z(n2748) );
  BUF_X2 U7930 ( .A(n2140), .Z(n2726) );
  XOR2_X1 U7931 ( .A(\mult_22/ab[18][42] ), .B(\mult_22/CARRYB[17][42] ), .Z(
        n2194) );
  XOR2_X1 U7932 ( .A(n2194), .B(\mult_22/SUMB[17][43] ), .Z(
        \mult_22/SUMB[18][42] ) );
  NAND2_X1 U7933 ( .A1(\mult_22/ab[18][42] ), .A2(\mult_22/CARRYB[17][42] ), 
        .ZN(n2195) );
  NAND2_X1 U7934 ( .A1(\mult_22/ab[18][42] ), .A2(\mult_22/SUMB[17][43] ), 
        .ZN(n2196) );
  NAND2_X1 U7935 ( .A1(\mult_22/CARRYB[17][42] ), .A2(\mult_22/SUMB[17][43] ), 
        .ZN(n2197) );
  NAND3_X1 U7936 ( .A1(n2195), .A2(n2196), .A3(n2197), .ZN(
        \mult_22/CARRYB[18][42] ) );
  NAND2_X1 U7937 ( .A1(\mult_22/ab[19][41] ), .A2(\mult_22/CARRYB[18][41] ), 
        .ZN(n2198) );
  NAND2_X1 U7938 ( .A1(\mult_22/ab[19][41] ), .A2(\mult_22/SUMB[18][42] ), 
        .ZN(n2199) );
  NAND2_X1 U7939 ( .A1(\mult_22/CARRYB[18][41] ), .A2(\mult_22/SUMB[18][42] ), 
        .ZN(n2200) );
  NAND3_X1 U7940 ( .A1(n2198), .A2(n2199), .A3(n2200), .ZN(
        \mult_22/CARRYB[19][41] ) );
  NOR3_X2 U7941 ( .A1(n2257), .A2(n809), .A3(n2158), .ZN(n1800) );
  NAND2_X1 U7942 ( .A1(\mult_22/SUMB[15][47] ), .A2(\mult_22/CARRYB[15][46] ), 
        .ZN(n2201) );
  NAND2_X1 U7943 ( .A1(\mult_22/SUMB[15][47] ), .A2(\mult_22/ab[16][46] ), 
        .ZN(n2202) );
  NAND2_X1 U7944 ( .A1(\mult_22/CARRYB[15][46] ), .A2(\mult_22/ab[16][46] ), 
        .ZN(n2203) );
  NAND3_X1 U7945 ( .A1(n2201), .A2(n2202), .A3(n2203), .ZN(
        \mult_22/CARRYB[16][46] ) );
  XNOR2_X1 U7946 ( .A(\mult_22/SUMB[4][61] ), .B(n2204), .ZN(
        \mult_22/SUMB[5][60] ) );
  XNOR2_X1 U7947 ( .A(\mult_22/CARRYB[4][60] ), .B(\mult_22/ab[5][60] ), .ZN(
        n2204) );
  NAND2_X1 U7948 ( .A1(n2191), .A2(\mult_22/SUMB[3][62] ), .ZN(n2205) );
  NAND2_X1 U7949 ( .A1(\mult_22/CARRYB[3][61] ), .A2(\mult_22/ab[4][61] ), 
        .ZN(n2206) );
  NAND2_X1 U7950 ( .A1(\mult_22/SUMB[3][62] ), .A2(\mult_22/ab[4][61] ), .ZN(
        n2207) );
  NAND3_X1 U7951 ( .A1(n2206), .A2(n2205), .A3(n2207), .ZN(
        \mult_22/CARRYB[4][61] ) );
  XNOR2_X1 U7952 ( .A(n2208), .B(n950), .ZN(\mult_22/SUMB[21][38] ) );
  AND2_X1 U7953 ( .A1(reg_mid_0[21]), .A2(reg_mid_1[38]), .ZN(n2208) );
  XNOR2_X1 U7954 ( .A(\mult_22/SUMB[28][33] ), .B(n2209), .ZN(
        \mult_22/SUMB[29][32] ) );
  XNOR2_X1 U7955 ( .A(\mult_22/CARRYB[28][32] ), .B(\mult_22/ab[29][32] ), 
        .ZN(n2209) );
  XNOR2_X1 U7956 ( .A(\mult_22/SUMB[33][30] ), .B(n2210), .ZN(
        \mult_22/SUMB[34][29] ) );
  XNOR2_X1 U7957 ( .A(\mult_22/CARRYB[33][29] ), .B(\mult_22/ab[34][29] ), 
        .ZN(n2210) );
  XNOR2_X1 U7958 ( .A(n2211), .B(\mult_22/SUMB[3][61] ), .ZN(
        \mult_22/SUMB[4][60] ) );
  XNOR2_X1 U7959 ( .A(\mult_22/CARRYB[3][60] ), .B(\mult_22/ab[4][60] ), .ZN(
        n2211) );
  XNOR2_X1 U7960 ( .A(\mult_22/CARRYB[23][32] ), .B(\mult_22/SUMB[23][33] ), 
        .ZN(n945) );
  XNOR2_X1 U7961 ( .A(n939), .B(n2212), .ZN(\mult_22/SUMB[28][30] ) );
  XNOR2_X1 U7962 ( .A(n693), .B(\mult_22/SUMB[27][31] ), .ZN(n2212) );
  XNOR2_X1 U7963 ( .A(\mult_22/CARRYB[31][29] ), .B(n2213), .ZN(n2332) );
  CLKBUF_X3 U7964 ( .A(n746), .Z(n2745) );
  OR2_X2 U7965 ( .A1(n2368), .A2(n2238), .ZN(n903) );
  OR2_X1 U7966 ( .A1(n2215), .A2(n1880), .ZN(n2214) );
  INV_X1 U7967 ( .A(n1879), .ZN(n2215) );
  AND2_X1 U7968 ( .A1(n1803), .A2(n1879), .ZN(n2216) );
  NAND2_X1 U7969 ( .A1(\mult_22/SUMB[4][61] ), .A2(\mult_22/CARRYB[4][60] ), 
        .ZN(n2217) );
  NAND2_X1 U7970 ( .A1(\mult_22/SUMB[4][61] ), .A2(\mult_22/ab[5][60] ), .ZN(
        n2218) );
  NAND2_X1 U7971 ( .A1(\mult_22/CARRYB[4][60] ), .A2(\mult_22/ab[5][60] ), 
        .ZN(n2219) );
  NAND3_X1 U7972 ( .A1(n2217), .A2(n2218), .A3(n2219), .ZN(
        \mult_22/CARRYB[5][60] ) );
  NAND2_X1 U7973 ( .A1(n1404), .A2(n1884), .ZN(n1402) );
  NAND2_X1 U7974 ( .A1(\mult_22/SUMB[33][30] ), .A2(\mult_22/CARRYB[33][29] ), 
        .ZN(n2220) );
  NAND2_X1 U7975 ( .A1(\mult_22/SUMB[33][30] ), .A2(\mult_22/ab[34][29] ), 
        .ZN(n2221) );
  NAND2_X1 U7976 ( .A1(\mult_22/CARRYB[33][29] ), .A2(\mult_22/ab[34][29] ), 
        .ZN(n2222) );
  NAND3_X1 U7977 ( .A1(n2220), .A2(n2221), .A3(n2222), .ZN(
        \mult_22/CARRYB[34][29] ) );
  AND2_X1 U7978 ( .A1(\mult_22/CARRYB[20][38] ), .A2(\mult_22/SUMB[20][39] ), 
        .ZN(n2223) );
  XNOR2_X1 U7979 ( .A(n2224), .B(\mult_22/SUMB[16][47] ), .ZN(
        \mult_22/SUMB[17][46] ) );
  XNOR2_X1 U7980 ( .A(\mult_22/ab[17][46] ), .B(\mult_22/CARRYB[16][46] ), 
        .ZN(n2224) );
  XNOR2_X1 U7981 ( .A(n2225), .B(\mult_22/SUMB[18][46] ), .ZN(
        \mult_22/SUMB[19][45] ) );
  XNOR2_X1 U7982 ( .A(\mult_22/ab[19][45] ), .B(\mult_22/CARRYB[18][45] ), 
        .ZN(n2225) );
  NAND2_X1 U7983 ( .A1(\mult_22/SUMB[3][61] ), .A2(\mult_22/CARRYB[3][60] ), 
        .ZN(n2226) );
  NAND2_X1 U7984 ( .A1(\mult_22/SUMB[3][61] ), .A2(\mult_22/ab[4][60] ), .ZN(
        n2227) );
  NAND2_X1 U7985 ( .A1(\mult_22/CARRYB[3][60] ), .A2(\mult_22/ab[4][60] ), 
        .ZN(n2228) );
  NAND3_X1 U7986 ( .A1(n2226), .A2(n2227), .A3(n2228), .ZN(
        \mult_22/CARRYB[4][60] ) );
  NAND2_X1 U7987 ( .A1(n1587), .A2(n1830), .ZN(n1586) );
  NAND2_X1 U7988 ( .A1(\mult_22/CARRYB[25][40] ), .A2(\mult_22/SUMB[25][41] ), 
        .ZN(n2229) );
  NAND2_X1 U7989 ( .A1(\mult_22/SUMB[25][41] ), .A2(\mult_22/ab[26][40] ), 
        .ZN(n2230) );
  NAND2_X1 U7990 ( .A1(\mult_22/CARRYB[25][40] ), .A2(\mult_22/ab[26][40] ), 
        .ZN(n2231) );
  NAND3_X1 U7991 ( .A1(n2229), .A2(n2230), .A3(n2231), .ZN(
        \mult_22/CARRYB[26][40] ) );
  NAND2_X1 U7992 ( .A1(n2182), .A2(n1803), .ZN(n1515) );
  OAI21_X1 U7993 ( .B1(n2093), .B2(n1395), .A(n1397), .ZN(n2232) );
  OAI21_X1 U7994 ( .B1(n2177), .B2(n1395), .A(n1397), .ZN(n1376) );
  CLKBUF_X1 U7995 ( .A(n1587), .Z(n2366) );
  XNOR2_X1 U7996 ( .A(\mult_22/SUMB[17][41] ), .B(\mult_22/CARRYB[17][40] ), 
        .ZN(n956) );
  XNOR2_X1 U7997 ( .A(n2233), .B(\mult_22/SUMB[17][46] ), .ZN(
        \mult_22/SUMB[18][45] ) );
  XNOR2_X1 U7998 ( .A(\mult_22/CARRYB[17][45] ), .B(\mult_22/ab[18][45] ), 
        .ZN(n2233) );
  XNOR2_X1 U7999 ( .A(\mult_22/SUMB[25][40] ), .B(n2234), .ZN(
        \mult_22/SUMB[26][39] ) );
  XNOR2_X1 U8000 ( .A(\mult_22/CARRYB[25][39] ), .B(\mult_22/ab[26][39] ), 
        .ZN(n2234) );
  NAND3_X1 U8001 ( .A1(n2307), .A2(n2308), .A3(n2309), .ZN(
        \mult_22/CARRYB[20][38] ) );
  XNOR2_X1 U8002 ( .A(\mult_22/SUMB[23][42] ), .B(n2235), .ZN(
        \mult_22/SUMB[24][41] ) );
  XNOR2_X1 U8003 ( .A(\mult_22/CARRYB[23][41] ), .B(\mult_22/ab[24][41] ), 
        .ZN(n2235) );
  XNOR2_X1 U8004 ( .A(\mult_22/SUMB[10][48] ), .B(n2236), .ZN(
        \mult_22/SUMB[11][47] ) );
  XNOR2_X1 U8005 ( .A(\mult_22/CARRYB[10][47] ), .B(\mult_22/ab[11][47] ), 
        .ZN(n2236) );
  XNOR2_X1 U8006 ( .A(n2237), .B(\mult_22/SUMB[16][43] ), .ZN(
        \mult_22/SUMB[17][42] ) );
  XNOR2_X1 U8007 ( .A(\mult_22/ab[17][42] ), .B(\mult_22/CARRYB[16][42] ), 
        .ZN(n2237) );
  XOR2_X1 U8008 ( .A(\mult_22/CARRYB[30][31] ), .B(\mult_22/ab[31][31] ), .Z(
        n2239) );
  XOR2_X1 U8009 ( .A(\mult_22/SUMB[30][32] ), .B(n2239), .Z(
        \mult_22/SUMB[31][31] ) );
  NAND2_X1 U8010 ( .A1(\mult_22/SUMB[30][32] ), .A2(\mult_22/CARRYB[30][31] ), 
        .ZN(n2240) );
  NAND2_X1 U8011 ( .A1(\mult_22/SUMB[30][32] ), .A2(\mult_22/ab[31][31] ), 
        .ZN(n2241) );
  NAND2_X1 U8012 ( .A1(\mult_22/CARRYB[30][31] ), .A2(\mult_22/ab[31][31] ), 
        .ZN(n2242) );
  NAND3_X1 U8013 ( .A1(n2240), .A2(n2241), .A3(n2242), .ZN(
        \mult_22/CARRYB[31][31] ) );
  XOR2_X1 U8014 ( .A(\mult_22/ab[30][32] ), .B(\mult_22/CARRYB[29][32] ), .Z(
        n2243) );
  XOR2_X1 U8015 ( .A(n2243), .B(\mult_22/SUMB[29][33] ), .Z(
        \mult_22/SUMB[30][32] ) );
  NAND2_X1 U8016 ( .A1(\mult_22/ab[29][33] ), .A2(\mult_22/CARRYB[28][33] ), 
        .ZN(n2244) );
  NAND2_X1 U8017 ( .A1(\mult_22/ab[29][33] ), .A2(\mult_22/SUMB[28][34] ), 
        .ZN(n2245) );
  NAND2_X1 U8018 ( .A1(\mult_22/CARRYB[28][33] ), .A2(\mult_22/SUMB[28][34] ), 
        .ZN(n2246) );
  NAND3_X1 U8019 ( .A1(n2244), .A2(n2245), .A3(n2246), .ZN(
        \mult_22/CARRYB[29][33] ) );
  NAND2_X1 U8020 ( .A1(\mult_22/ab[30][32] ), .A2(\mult_22/CARRYB[29][32] ), 
        .ZN(n2247) );
  NAND2_X1 U8021 ( .A1(\mult_22/ab[30][32] ), .A2(\mult_22/SUMB[29][33] ), 
        .ZN(n2248) );
  NAND2_X1 U8022 ( .A1(\mult_22/CARRYB[29][32] ), .A2(\mult_22/SUMB[29][33] ), 
        .ZN(n2249) );
  NAND3_X1 U8023 ( .A1(n2247), .A2(n2248), .A3(n2249), .ZN(
        \mult_22/CARRYB[30][32] ) );
  XOR2_X1 U8024 ( .A(\mult_22/ab[16][43] ), .B(\mult_22/CARRYB[15][43] ), .Z(
        n2250) );
  XOR2_X1 U8025 ( .A(n2250), .B(\mult_22/SUMB[15][44] ), .Z(
        \mult_22/SUMB[16][43] ) );
  NAND2_X1 U8026 ( .A1(\mult_22/ab[16][43] ), .A2(\mult_22/CARRYB[15][43] ), 
        .ZN(n2251) );
  NAND2_X1 U8027 ( .A1(\mult_22/ab[16][43] ), .A2(\mult_22/SUMB[15][44] ), 
        .ZN(n2252) );
  NAND2_X1 U8028 ( .A1(\mult_22/CARRYB[15][43] ), .A2(\mult_22/SUMB[15][44] ), 
        .ZN(n2253) );
  NAND3_X1 U8029 ( .A1(n2251), .A2(n2252), .A3(n2253), .ZN(
        \mult_22/CARRYB[16][43] ) );
  NAND2_X1 U8030 ( .A1(\mult_22/ab[17][42] ), .A2(\mult_22/CARRYB[16][42] ), 
        .ZN(n2254) );
  NAND2_X1 U8031 ( .A1(\mult_22/ab[17][42] ), .A2(\mult_22/SUMB[16][43] ), 
        .ZN(n2255) );
  NAND2_X1 U8032 ( .A1(\mult_22/CARRYB[16][42] ), .A2(\mult_22/SUMB[16][43] ), 
        .ZN(n2256) );
  NAND3_X1 U8033 ( .A1(n2254), .A2(n2255), .A3(n2256), .ZN(
        \mult_22/CARRYB[17][42] ) );
  INV_X1 U8034 ( .A(n2187), .ZN(n2257) );
  NAND2_X1 U8035 ( .A1(\mult_22/SUMB[23][42] ), .A2(\mult_22/CARRYB[23][41] ), 
        .ZN(n2258) );
  NAND2_X1 U8036 ( .A1(\mult_22/SUMB[23][42] ), .A2(\mult_22/ab[24][41] ), 
        .ZN(n2259) );
  NAND2_X1 U8037 ( .A1(\mult_22/CARRYB[23][41] ), .A2(\mult_22/ab[24][41] ), 
        .ZN(n2260) );
  NAND3_X1 U8038 ( .A1(n2258), .A2(n2259), .A3(n2260), .ZN(
        \mult_22/CARRYB[24][41] ) );
  XNOR2_X1 U8039 ( .A(\mult_22/SUMB[2][62] ), .B(n2261), .ZN(
        \mult_22/SUMB[3][61] ) );
  XNOR2_X1 U8040 ( .A(\mult_22/CARRYB[2][61] ), .B(\mult_22/ab[3][61] ), .ZN(
        n2261) );
  NAND2_X1 U8041 ( .A1(\mult_22/SUMB[25][40] ), .A2(\mult_22/CARRYB[25][39] ), 
        .ZN(n2262) );
  NAND2_X1 U8042 ( .A1(\mult_22/SUMB[25][40] ), .A2(\mult_22/ab[26][39] ), 
        .ZN(n2263) );
  NAND2_X1 U8043 ( .A1(\mult_22/CARRYB[25][39] ), .A2(\mult_22/ab[26][39] ), 
        .ZN(n2264) );
  NAND3_X1 U8044 ( .A1(n2262), .A2(n2263), .A3(n2264), .ZN(
        \mult_22/CARRYB[26][39] ) );
  NAND2_X1 U8045 ( .A1(\mult_22/CARRYB[2][62] ), .A2(\mult_22/ab[2][63] ), 
        .ZN(n2265) );
  NAND2_X1 U8046 ( .A1(\mult_22/CARRYB[2][62] ), .A2(\mult_22/ab[3][62] ), 
        .ZN(n2266) );
  NAND2_X1 U8047 ( .A1(\mult_22/ab[2][63] ), .A2(\mult_22/ab[3][62] ), .ZN(
        n2267) );
  NAND3_X1 U8048 ( .A1(n2265), .A2(n2266), .A3(n2267), .ZN(
        \mult_22/CARRYB[3][62] ) );
  XNOR2_X1 U8049 ( .A(n958), .B(n2268), .ZN(\mult_22/SUMB[11][46] ) );
  AND2_X1 U8050 ( .A1(reg_mid_0[11]), .A2(reg_mid_1[46]), .ZN(n2268) );
  NAND2_X1 U8051 ( .A1(\mult_22/ab[17][46] ), .A2(\mult_22/CARRYB[16][46] ), 
        .ZN(n2269) );
  NAND2_X1 U8052 ( .A1(\mult_22/ab[17][46] ), .A2(\mult_22/SUMB[16][47] ), 
        .ZN(n2270) );
  NAND2_X1 U8053 ( .A1(\mult_22/CARRYB[16][46] ), .A2(\mult_22/SUMB[16][47] ), 
        .ZN(n2271) );
  NAND3_X1 U8054 ( .A1(n2269), .A2(n2270), .A3(n2271), .ZN(
        \mult_22/CARRYB[17][46] ) );
  NAND2_X1 U8055 ( .A1(\mult_22/ab[18][45] ), .A2(\mult_22/CARRYB[17][45] ), 
        .ZN(n2272) );
  NAND2_X1 U8056 ( .A1(\mult_22/ab[18][45] ), .A2(\mult_22/SUMB[17][46] ), 
        .ZN(n2273) );
  NAND2_X1 U8057 ( .A1(\mult_22/CARRYB[17][45] ), .A2(\mult_22/SUMB[17][46] ), 
        .ZN(n2274) );
  NAND3_X1 U8058 ( .A1(n2272), .A2(n2273), .A3(n2274), .ZN(
        \mult_22/CARRYB[18][45] ) );
  XNOR2_X1 U8059 ( .A(n935), .B(n2275), .ZN(\mult_22/SUMB[3][56] ) );
  XNOR2_X1 U8060 ( .A(n740), .B(\mult_22/SUMB[2][57] ), .ZN(n2275) );
  XNOR2_X1 U8061 ( .A(\mult_22/SUMB[8][51] ), .B(n2276), .ZN(
        \mult_22/SUMB[9][50] ) );
  XNOR2_X1 U8062 ( .A(\mult_22/CARRYB[8][50] ), .B(\mult_22/ab[9][50] ), .ZN(
        n2276) );
  XNOR2_X1 U8063 ( .A(n2277), .B(\mult_22/CARRYB[17][46] ), .ZN(n2311) );
  XNOR2_X1 U8064 ( .A(n2278), .B(\mult_22/SUMB[19][45] ), .ZN(
        \mult_22/SUMB[20][44] ) );
  XNOR2_X1 U8065 ( .A(\mult_22/ab[20][44] ), .B(\mult_22/CARRYB[19][44] ), 
        .ZN(n2278) );
  NAND2_X1 U8066 ( .A1(n1567), .A2(n1831), .ZN(n1565) );
  XOR2_X1 U8067 ( .A(\mult_22/SUMB[25][36] ), .B(n2279), .Z(
        \mult_22/SUMB[26][35] ) );
  NAND2_X1 U8068 ( .A1(\mult_22/SUMB[25][36] ), .A2(\mult_22/CARRYB[25][35] ), 
        .ZN(n2280) );
  NAND2_X1 U8069 ( .A1(\mult_22/SUMB[25][36] ), .A2(n2070), .ZN(n2281) );
  NAND2_X1 U8070 ( .A1(\mult_22/CARRYB[25][35] ), .A2(n2070), .ZN(n2282) );
  NAND3_X1 U8071 ( .A1(n2280), .A2(n2281), .A3(n2282), .ZN(
        \mult_22/CARRYB[26][35] ) );
  NAND2_X1 U8072 ( .A1(\mult_22/SUMB[10][48] ), .A2(\mult_22/CARRYB[10][47] ), 
        .ZN(n2283) );
  NAND2_X1 U8073 ( .A1(\mult_22/SUMB[10][48] ), .A2(\mult_22/ab[11][47] ), 
        .ZN(n2284) );
  NAND2_X1 U8074 ( .A1(\mult_22/CARRYB[10][47] ), .A2(\mult_22/ab[11][47] ), 
        .ZN(n2285) );
  NAND3_X1 U8075 ( .A1(n2283), .A2(n2284), .A3(n2285), .ZN(
        \mult_22/CARRYB[11][47] ) );
  XNOR2_X1 U8076 ( .A(n887), .B(n2286), .ZN(\mult_22/n322 ) );
  AND2_X1 U8077 ( .A1(reg_mid_1[57]), .A2(reg_mid_0[0]), .ZN(n2286) );
  AND2_X1 U8078 ( .A1(n2159), .A2(\mult_22/CARRYB[63][3] ), .ZN(n2287) );
  NAND2_X1 U8079 ( .A1(\mult_22/SUMB[28][33] ), .A2(\mult_22/CARRYB[28][32] ), 
        .ZN(n2288) );
  NAND2_X1 U8080 ( .A1(\mult_22/SUMB[28][33] ), .A2(\mult_22/ab[29][32] ), 
        .ZN(n2289) );
  NAND2_X1 U8081 ( .A1(\mult_22/CARRYB[28][32] ), .A2(\mult_22/ab[29][32] ), 
        .ZN(n2290) );
  NAND3_X1 U8082 ( .A1(n2288), .A2(n2289), .A3(n2290), .ZN(
        \mult_22/CARRYB[29][32] ) );
  CLKBUF_X3 U8083 ( .A(n2158), .Z(n2741) );
  BUF_X2 U8084 ( .A(n2158), .Z(n2739) );
  XNOR2_X1 U8085 ( .A(n2291), .B(\mult_22/SUMB[20][44] ), .ZN(
        \mult_22/SUMB[21][43] ) );
  XNOR2_X1 U8086 ( .A(\mult_22/ab[21][43] ), .B(\mult_22/CARRYB[20][43] ), 
        .ZN(n2291) );
  NAND2_X1 U8087 ( .A1(n1515), .A2(n1880), .ZN(n1491) );
  XNOR2_X1 U8088 ( .A(n2294), .B(\mult_22/SUMB[2][56] ), .ZN(
        \mult_22/SUMB[3][55] ) );
  XNOR2_X1 U8089 ( .A(\mult_22/ab[3][55] ), .B(\mult_22/CARRYB[2][55] ), .ZN(
        n2294) );
  XNOR2_X1 U8090 ( .A(n2296), .B(n2295), .ZN(\mult_22/SUMB[4][52] ) );
  XNOR2_X1 U8091 ( .A(\mult_22/SUMB[3][53] ), .B(n737), .ZN(n2296) );
  XNOR2_X1 U8092 ( .A(n2297), .B(\mult_22/CARRYB[25][34] ), .ZN(n942) );
  AND2_X1 U8093 ( .A1(reg_mid_0[26]), .A2(reg_mid_1[34]), .ZN(n2297) );
  OR2_X1 U8094 ( .A1(n1608), .A2(n1614), .ZN(n2298) );
  XOR2_X1 U8095 ( .A(\mult_22/ab[2][56] ), .B(\mult_22/n59 ), .Z(n2299) );
  XOR2_X1 U8096 ( .A(n2299), .B(\mult_22/n159 ), .Z(\mult_22/SUMB[2][56] ) );
  NAND2_X1 U8097 ( .A1(\mult_22/ab[2][56] ), .A2(\mult_22/n59 ), .ZN(n2300) );
  NAND2_X1 U8098 ( .A1(\mult_22/ab[2][56] ), .A2(\mult_22/n159 ), .ZN(n2301)
         );
  NAND2_X1 U8099 ( .A1(\mult_22/n59 ), .A2(\mult_22/n159 ), .ZN(n2302) );
  NAND3_X1 U8100 ( .A1(n2300), .A2(n2301), .A3(n2302), .ZN(
        \mult_22/CARRYB[2][56] ) );
  NAND2_X1 U8101 ( .A1(\mult_22/ab[3][55] ), .A2(\mult_22/CARRYB[2][55] ), 
        .ZN(n2303) );
  NAND2_X1 U8102 ( .A1(\mult_22/ab[3][55] ), .A2(\mult_22/SUMB[2][56] ), .ZN(
        n2304) );
  NAND2_X1 U8103 ( .A1(\mult_22/CARRYB[2][55] ), .A2(\mult_22/SUMB[2][56] ), 
        .ZN(n2305) );
  NAND3_X1 U8104 ( .A1(n2303), .A2(n2304), .A3(n2305), .ZN(
        \mult_22/CARRYB[3][55] ) );
  XOR2_X1 U8105 ( .A(\mult_22/CARRYB[19][38] ), .B(\mult_22/ab[20][38] ), .Z(
        n2306) );
  XOR2_X1 U8106 ( .A(\mult_22/SUMB[19][39] ), .B(n2306), .Z(
        \mult_22/SUMB[20][38] ) );
  NAND2_X1 U8107 ( .A1(\mult_22/SUMB[19][39] ), .A2(\mult_22/CARRYB[19][38] ), 
        .ZN(n2307) );
  NAND2_X1 U8108 ( .A1(\mult_22/SUMB[19][39] ), .A2(\mult_22/ab[20][38] ), 
        .ZN(n2308) );
  NAND2_X1 U8109 ( .A1(\mult_22/CARRYB[19][38] ), .A2(\mult_22/ab[20][38] ), 
        .ZN(n2309) );
  AOI21_X1 U8110 ( .B1(n2179), .B2(n638), .A(n1336), .ZN(n2310) );
  NOR2_X1 U8111 ( .A1(n2353), .A2(n621), .ZN(n1614) );
  AOI21_X1 U8112 ( .B1(n1335), .B2(n638), .A(n1336), .ZN(n1332) );
  XOR2_X1 U8113 ( .A(n2311), .B(\mult_22/SUMB[17][47] ), .Z(
        \mult_22/SUMB[18][46] ) );
  NAND2_X1 U8114 ( .A1(\mult_22/ab[18][46] ), .A2(\mult_22/CARRYB[17][46] ), 
        .ZN(n2312) );
  NAND2_X1 U8115 ( .A1(\mult_22/ab[18][46] ), .A2(\mult_22/SUMB[17][47] ), 
        .ZN(n2313) );
  NAND2_X1 U8116 ( .A1(\mult_22/CARRYB[17][46] ), .A2(\mult_22/SUMB[17][47] ), 
        .ZN(n2314) );
  NAND3_X1 U8117 ( .A1(n2312), .A2(n2313), .A3(n2314), .ZN(
        \mult_22/CARRYB[18][46] ) );
  NAND2_X1 U8118 ( .A1(\mult_22/ab[19][45] ), .A2(\mult_22/CARRYB[18][45] ), 
        .ZN(n2315) );
  NAND2_X1 U8119 ( .A1(\mult_22/ab[19][45] ), .A2(\mult_22/SUMB[18][46] ), 
        .ZN(n2316) );
  NAND2_X1 U8120 ( .A1(\mult_22/CARRYB[18][45] ), .A2(\mult_22/SUMB[18][46] ), 
        .ZN(n2317) );
  NAND3_X1 U8121 ( .A1(n2315), .A2(n2316), .A3(n2317), .ZN(
        \mult_22/CARRYB[19][45] ) );
  NAND2_X1 U8122 ( .A1(\mult_22/SUMB[2][62] ), .A2(\mult_22/CARRYB[2][61] ), 
        .ZN(n2318) );
  NAND2_X1 U8123 ( .A1(\mult_22/SUMB[2][62] ), .A2(\mult_22/ab[3][61] ), .ZN(
        n2319) );
  NAND2_X1 U8124 ( .A1(\mult_22/CARRYB[2][61] ), .A2(\mult_22/ab[3][61] ), 
        .ZN(n2320) );
  NAND3_X1 U8125 ( .A1(n2318), .A2(n2319), .A3(n2320), .ZN(
        \mult_22/CARRYB[3][61] ) );
  OAI21_X1 U8126 ( .B1(n2310), .B2(n1331), .A(n1333), .ZN(n2321) );
  INV_X1 U8127 ( .A(n2373), .ZN(n2322) );
  NAND2_X1 U8128 ( .A1(\mult_22/ab[20][44] ), .A2(\mult_22/CARRYB[19][44] ), 
        .ZN(n2323) );
  NAND2_X1 U8129 ( .A1(\mult_22/ab[20][44] ), .A2(\mult_22/SUMB[19][45] ), 
        .ZN(n2324) );
  NAND2_X1 U8130 ( .A1(\mult_22/CARRYB[19][44] ), .A2(\mult_22/SUMB[19][45] ), 
        .ZN(n2325) );
  NAND3_X1 U8131 ( .A1(n2323), .A2(n2324), .A3(n2325), .ZN(
        \mult_22/CARRYB[20][44] ) );
  NAND2_X1 U8132 ( .A1(\mult_22/ab[21][43] ), .A2(\mult_22/CARRYB[20][43] ), 
        .ZN(n2326) );
  NAND2_X1 U8133 ( .A1(\mult_22/ab[21][43] ), .A2(\mult_22/SUMB[20][44] ), 
        .ZN(n2327) );
  NAND2_X1 U8134 ( .A1(\mult_22/CARRYB[20][43] ), .A2(\mult_22/SUMB[20][44] ), 
        .ZN(n2328) );
  NAND3_X1 U8135 ( .A1(n2326), .A2(n2327), .A3(n2328), .ZN(
        \mult_22/CARRYB[21][43] ) );
  NAND2_X1 U8136 ( .A1(\mult_22/SUMB[8][51] ), .A2(\mult_22/CARRYB[8][50] ), 
        .ZN(n2329) );
  NAND2_X1 U8137 ( .A1(\mult_22/SUMB[8][51] ), .A2(\mult_22/ab[9][50] ), .ZN(
        n2330) );
  NAND2_X1 U8138 ( .A1(\mult_22/CARRYB[8][50] ), .A2(\mult_22/ab[9][50] ), 
        .ZN(n2331) );
  NAND3_X1 U8139 ( .A1(n2329), .A2(n2330), .A3(n2331), .ZN(
        \mult_22/CARRYB[9][50] ) );
  XOR2_X1 U8140 ( .A(\mult_22/SUMB[31][30] ), .B(n2332), .Z(
        \mult_22/SUMB[32][29] ) );
  NAND2_X1 U8141 ( .A1(\mult_22/SUMB[31][30] ), .A2(\mult_22/CARRYB[31][29] ), 
        .ZN(n2333) );
  NAND2_X1 U8142 ( .A1(\mult_22/SUMB[31][30] ), .A2(\mult_22/ab[32][29] ), 
        .ZN(n2334) );
  NAND2_X1 U8143 ( .A1(\mult_22/CARRYB[31][29] ), .A2(\mult_22/ab[32][29] ), 
        .ZN(n2335) );
  NAND3_X1 U8144 ( .A1(n2333), .A2(n2334), .A3(n2335), .ZN(
        \mult_22/CARRYB[32][29] ) );
  OAI21_X1 U8145 ( .B1(n1452), .B2(n2132), .A(n1454), .ZN(n2336) );
  OR2_X1 U8146 ( .A1(n595), .A2(n1512), .ZN(n2337) );
  OR2_X1 U8147 ( .A1(n1513), .A2(n1514), .ZN(n2338) );
  OR2_X1 U8148 ( .A1(n1609), .A2(n1608), .ZN(n2339) );
  OR2_X1 U8149 ( .A1(n1610), .A2(n1611), .ZN(n2340) );
  NAND3_X1 U8150 ( .A1(n2339), .A2(n1612), .A3(n2340), .ZN(n1587) );
  OAI211_X1 U8151 ( .C1(n1583), .C2(n1584), .A(n2096), .B(n1585), .ZN(n2341)
         );
  OAI22_X1 U8152 ( .A1(n2180), .A2(n643), .B1(n1312), .B2(n1313), .ZN(n2342)
         );
  XNOR2_X1 U8153 ( .A(n2183), .B(\mult_22/SUMB[21][39] ), .ZN(n2347) );
  XNOR2_X1 U8154 ( .A(\mult_22/CARRYB[32][28] ), .B(\mult_22/SUMB[32][29] ), 
        .ZN(n938) );
  XNOR2_X1 U8155 ( .A(n2343), .B(n938), .ZN(\mult_22/SUMB[33][28] ) );
  AND2_X1 U8156 ( .A1(reg_mid_0[33]), .A2(reg_mid_1[28]), .ZN(n2343) );
  CLKBUF_X1 U8157 ( .A(n1869), .Z(n2845) );
  CLKBUF_X1 U8158 ( .A(n1852), .Z(n2850) );
  NOR2_X2 U8159 ( .A1(n1534), .A2(n1535), .ZN(n1521) );
  XOR2_X1 U8160 ( .A(n1427), .B(n2344), .Z(N229) );
  NAND2_X1 U8161 ( .A1(n616), .A2(n1421), .ZN(n2344) );
  XOR2_X1 U8162 ( .A(n1595), .B(n2345), .Z(N201) );
  NAND2_X1 U8163 ( .A1(n1585), .A2(n583), .ZN(n2345) );
  BUF_X2 U8164 ( .A(n1821), .Z(n2684) );
  CLKBUF_X3 U8165 ( .A(n1881), .Z(n2692) );
  BUF_X2 U8166 ( .A(n1881), .Z(n2691) );
  BUF_X2 U8167 ( .A(n754), .Z(n2703) );
  CLKBUF_X1 U8168 ( .A(n1822), .Z(n2721) );
  BUF_X2 U8169 ( .A(n753), .Z(n2709) );
  CLKBUF_X1 U8170 ( .A(n754), .Z(n2701) );
  BUF_X2 U8171 ( .A(n2360), .Z(n2666) );
  BUF_X2 U8172 ( .A(n2361), .Z(n2660) );
  BUF_X2 U8173 ( .A(n1813), .Z(n2642) );
  BUF_X2 U8174 ( .A(n1818), .Z(n2630) );
  CLKBUF_X3 U8175 ( .A(n1810), .Z(n2757) );
  BUF_X2 U8176 ( .A(n1810), .Z(n2758) );
  CLKBUF_X1 U8177 ( .A(n1809), .Z(n2696) );
  CLKBUF_X1 U8178 ( .A(n1837), .Z(n2459) );
  CLKBUF_X1 U8179 ( .A(n1861), .Z(n2447) );
  CLKBUF_X1 U8180 ( .A(n1844), .Z(n2435) );
  CLKBUF_X1 U8181 ( .A(n1863), .Z(n2453) );
  CLKBUF_X1 U8182 ( .A(n1845), .Z(n2429) );
  CLKBUF_X1 U8183 ( .A(n1843), .Z(n2465) );
  CLKBUF_X1 U8184 ( .A(n1832), .Z(n2423) );
  CLKBUF_X1 U8185 ( .A(n1835), .Z(n2471) );
  CLKBUF_X1 U8186 ( .A(n2362), .Z(n2652) );
  CLKBUF_X1 U8187 ( .A(n1847), .Z(n2411) );
  CLKBUF_X1 U8188 ( .A(n1846), .Z(n2417) );
  CLKBUF_X1 U8189 ( .A(n1821), .Z(n2685) );
  CLKBUF_X1 U8190 ( .A(n1836), .Z(n2477) );
  CLKBUF_X1 U8191 ( .A(n1825), .Z(n2640) );
  CLKBUF_X1 U8192 ( .A(n1824), .Z(n2624) );
  CLKBUF_X1 U8193 ( .A(n1874), .Z(n2443) );
  CLKBUF_X1 U8194 ( .A(n1842), .Z(n2483) );
  CLKBUF_X1 U8195 ( .A(n1824), .Z(n2628) );
  CLKBUF_X1 U8196 ( .A(n1841), .Z(n2489) );
  CLKBUF_X1 U8197 ( .A(n1873), .Z(n2528) );
  CLKBUF_X1 U8198 ( .A(n1840), .Z(n2495) );
  CLKBUF_X1 U8199 ( .A(n1883), .Z(n2576) );
  CLKBUF_X1 U8200 ( .A(n1839), .Z(n2501) );
  CLKBUF_X1 U8201 ( .A(n1826), .Z(n2676) );
  CLKBUF_X1 U8202 ( .A(n1838), .Z(n2507) );
  CLKBUF_X1 U8203 ( .A(n1833), .Z(n2519) );
  CLKBUF_X1 U8204 ( .A(n1825), .Z(n2636) );
  CLKBUF_X1 U8205 ( .A(n1834), .Z(n2513) );
  CLKBUF_X1 U8206 ( .A(n1864), .Z(n2531) );
  CLKBUF_X1 U8207 ( .A(n1816), .Z(n2567) );
  CLKBUF_X1 U8208 ( .A(n1862), .Z(n2537) );
  CLKBUF_X1 U8209 ( .A(n1865), .Z(n2543) );
  CLKBUF_X1 U8210 ( .A(n1823), .Z(n2561) );
  CLKBUF_X1 U8211 ( .A(n1873), .Z(n2527) );
  CLKBUF_X1 U8212 ( .A(n1856), .Z(n2555) );
  CLKBUF_X1 U8213 ( .A(n1868), .Z(n2549) );
  CLKBUF_X1 U8214 ( .A(n1817), .Z(n2578) );
  CLKBUF_X1 U8215 ( .A(n2158), .Z(n2737) );
  CLKBUF_X1 U8216 ( .A(n746), .Z(n2743) );
  CLKBUF_X1 U8217 ( .A(n2140), .Z(n2728) );
  CLKBUF_X1 U8218 ( .A(n748), .Z(n2734) );
  CLKBUF_X1 U8219 ( .A(n1822), .Z(n2722) );
  CLKBUF_X1 U8220 ( .A(n753), .Z(n2707) );
  CLKBUF_X1 U8221 ( .A(n2140), .Z(n2729) );
  CLKBUF_X1 U8222 ( .A(n748), .Z(n2735) );
  CLKBUF_X1 U8223 ( .A(n1822), .Z(n2723) );
  CLKBUF_X1 U8224 ( .A(n1826), .Z(n2675) );
  CLKBUF_X1 U8225 ( .A(n2362), .Z(n2648) );
  CLKBUF_X1 U8226 ( .A(n2111), .Z(n2750) );
  CLKBUF_X1 U8227 ( .A(n1813), .Z(n2643) );
  CLKBUF_X1 U8228 ( .A(n2361), .Z(n2661) );
  CLKBUF_X1 U8229 ( .A(n1812), .Z(n2619) );
  CLKBUF_X1 U8230 ( .A(n1818), .Z(n2631) );
  CLKBUF_X1 U8231 ( .A(n2363), .Z(n2655) );
  CLKBUF_X1 U8232 ( .A(n1824), .Z(n2627) );
  CLKBUF_X1 U8233 ( .A(n1883), .Z(n2575) );
  CLKBUF_X1 U8234 ( .A(n2111), .Z(n2749) );
  CLKBUF_X1 U8235 ( .A(n1825), .Z(n2639) );
  CLKBUF_X1 U8236 ( .A(n2359), .Z(n2679) );
  CLKBUF_X1 U8237 ( .A(n2362), .Z(n2651) );
  CLKBUF_X1 U8238 ( .A(n1820), .Z(n2613) );
  CLKBUF_X1 U8239 ( .A(n2360), .Z(n2667) );
  CLKBUF_X1 U8240 ( .A(n1881), .Z(n2694) );
  CLKBUF_X1 U8241 ( .A(n1819), .Z(n2584) );
  CLKBUF_X1 U8242 ( .A(n2140), .Z(n2725) );
  CLKBUF_X1 U8243 ( .A(n1826), .Z(n2672) );
  CLKBUF_X1 U8244 ( .A(n1822), .Z(n2719) );
  CLKBUF_X1 U8245 ( .A(n1881), .Z(n2690) );
  CLKBUF_X1 U8246 ( .A(n748), .Z(n2731) );
  CLKBUF_X1 U8247 ( .A(n1811), .Z(n2590) );
  CLKBUF_X1 U8248 ( .A(n1882), .Z(n2608) );
  CLKBUF_X1 U8249 ( .A(n1815), .Z(n2596) );
  CLKBUF_X1 U8250 ( .A(n1814), .Z(n2602) );
  BUF_X2 U8251 ( .A(n1845), .Z(n2428) );
  BUF_X2 U8252 ( .A(n1846), .Z(n2416) );
  BUF_X2 U8253 ( .A(n1832), .Z(n2422) );
  BUF_X2 U8254 ( .A(n1844), .Z(n2434) );
  BUF_X2 U8255 ( .A(n1838), .Z(n2506) );
  BUF_X2 U8256 ( .A(n1843), .Z(n2464) );
  BUF_X2 U8257 ( .A(n1839), .Z(n2500) );
  BUF_X2 U8258 ( .A(n1835), .Z(n2470) );
  BUF_X2 U8259 ( .A(n1836), .Z(n2476) );
  BUF_X2 U8260 ( .A(n1834), .Z(n2512) );
  CLKBUF_X3 U8261 ( .A(n1854), .Z(n2392) );
  BUF_X2 U8262 ( .A(n1840), .Z(n2494) );
  BUF_X2 U8263 ( .A(n1842), .Z(n2482) );
  BUF_X2 U8264 ( .A(n1841), .Z(n2488) );
  BUF_X2 U8265 ( .A(n1820), .Z(n2612) );
  BUF_X2 U8266 ( .A(n1882), .Z(n2607) );
  BUF_X2 U8267 ( .A(n1833), .Z(n2518) );
  BUF_X2 U8268 ( .A(n1814), .Z(n2601) );
  BUF_X2 U8269 ( .A(n1812), .Z(n2618) );
  BUF_X2 U8270 ( .A(n1815), .Z(n2595) );
  BUF_X2 U8271 ( .A(n1811), .Z(n2589) );
  BUF_X2 U8272 ( .A(n1819), .Z(n2583) );
  BUF_X2 U8273 ( .A(n1847), .Z(n2410) );
  BUF_X2 U8274 ( .A(n1837), .Z(n2458) );
  CLKBUF_X3 U8275 ( .A(n1855), .Z(n2386) );
  BUF_X2 U8276 ( .A(n1816), .Z(n2566) );
  BUF_X2 U8277 ( .A(n1817), .Z(n2577) );
  CLKBUF_X1 U8278 ( .A(n1829), .Z(n2768) );
  CLKBUF_X1 U8279 ( .A(n1810), .Z(n2756) );
  CLKBUF_X1 U8280 ( .A(n1827), .Z(n2762) );
  CLKBUF_X1 U8281 ( .A(n1828), .Z(n2774) );
  CLKBUF_X1 U8282 ( .A(n1878), .Z(n2780) );
  CLKBUF_X1 U8283 ( .A(n1829), .Z(n2766) );
  CLKBUF_X1 U8284 ( .A(n1810), .Z(n2755) );
  CLKBUF_X1 U8285 ( .A(n1810), .Z(n2754) );
  CLKBUF_X1 U8286 ( .A(n1827), .Z(n2760) );
  CLKBUF_X1 U8287 ( .A(n1827), .Z(n2761) );
  CLKBUF_X1 U8288 ( .A(n1829), .Z(n2767) );
  CLKBUF_X1 U8289 ( .A(n1828), .Z(n2772) );
  CLKBUF_X1 U8290 ( .A(n1828), .Z(n2773) );
  CLKBUF_X1 U8291 ( .A(n1877), .Z(n2786) );
  CLKBUF_X1 U8292 ( .A(n1878), .Z(n2779) );
  CLKBUF_X1 U8293 ( .A(n1877), .Z(n2785) );
  CLKBUF_X1 U8294 ( .A(n753), .Z(n2706) );
  CLKBUF_X1 U8295 ( .A(n1820), .Z(n2616) );
  CLKBUF_X1 U8296 ( .A(n1874), .Z(n2444) );
  CLKBUF_X1 U8297 ( .A(n1875), .Z(n2408) );
  CLKBUF_X1 U8298 ( .A(n1812), .Z(n2622) );
  CLKBUF_X1 U8299 ( .A(n1882), .Z(n2611) );
  CLKBUF_X1 U8300 ( .A(n1818), .Z(n2634) );
  CLKBUF_X1 U8301 ( .A(n1876), .Z(n2384) );
  CLKBUF_X1 U8302 ( .A(n1853), .Z(n2399) );
  CLKBUF_X1 U8303 ( .A(n1875), .Z(n2407) );
  CLKBUF_X1 U8304 ( .A(n1855), .Z(n2387) );
  CLKBUF_X1 U8305 ( .A(n1854), .Z(n2393) );
  CLKBUF_X1 U8306 ( .A(n1813), .Z(n2646) );
  CLKBUF_X1 U8307 ( .A(n1876), .Z(n2383) );
  CLKBUF_X1 U8308 ( .A(n1847), .Z(n2414) );
  CLKBUF_X1 U8309 ( .A(n1855), .Z(n2390) );
  CLKBUF_X1 U8310 ( .A(n753), .Z(n2710) );
  CLKBUF_X1 U8311 ( .A(n1854), .Z(n2396) );
  CLKBUF_X1 U8312 ( .A(n746), .Z(n2746) );
  CLKBUF_X1 U8313 ( .A(n2111), .Z(n2752) );
  CLKBUF_X1 U8314 ( .A(n1819), .Z(n2587) );
  CLKBUF_X1 U8315 ( .A(n1811), .Z(n2593) );
  CLKBUF_X1 U8316 ( .A(n2363), .Z(n2658) );
  CLKBUF_X1 U8317 ( .A(n1823), .Z(n2564) );
  CLKBUF_X1 U8318 ( .A(n1814), .Z(n2605) );
  CLKBUF_X1 U8319 ( .A(n1815), .Z(n2599) );
  CLKBUF_X1 U8320 ( .A(n1868), .Z(n2552) );
  CLKBUF_X1 U8321 ( .A(n1817), .Z(n2581) );
  CLKBUF_X1 U8322 ( .A(n2360), .Z(n2670) );
  CLKBUF_X1 U8323 ( .A(n1856), .Z(n2558) );
  CLKBUF_X1 U8324 ( .A(n1816), .Z(n2570) );
  CLKBUF_X1 U8325 ( .A(n1840), .Z(n2498) );
  CLKBUF_X1 U8326 ( .A(n1839), .Z(n2504) );
  CLKBUF_X1 U8327 ( .A(n1838), .Z(n2510) );
  CLKBUF_X1 U8328 ( .A(n1834), .Z(n2516) );
  CLKBUF_X1 U8329 ( .A(n1833), .Z(n2522) );
  CLKBUF_X1 U8330 ( .A(n1864), .Z(n2534) );
  CLKBUF_X1 U8331 ( .A(n1862), .Z(n2540) );
  CLKBUF_X1 U8332 ( .A(n1865), .Z(n2546) );
  CLKBUF_X1 U8333 ( .A(n2361), .Z(n2664) );
  CLKBUF_X1 U8334 ( .A(n2359), .Z(n2682) );
  CLKBUF_X1 U8335 ( .A(n754), .Z(n2704) );
  CLKBUF_X1 U8336 ( .A(n2158), .Z(n2740) );
  CLKBUF_X1 U8337 ( .A(n1821), .Z(n2688) );
  CLKBUF_X1 U8338 ( .A(n1883), .Z(n2572) );
  CLKBUF_X1 U8339 ( .A(n1873), .Z(n2524) );
  CLKBUF_X1 U8340 ( .A(n1844), .Z(n2438) );
  CLKBUF_X1 U8341 ( .A(n1841), .Z(n2492) );
  CLKBUF_X1 U8342 ( .A(n1842), .Z(n2486) );
  CLKBUF_X1 U8343 ( .A(n1836), .Z(n2480) );
  CLKBUF_X1 U8344 ( .A(n1835), .Z(n2474) );
  CLKBUF_X1 U8345 ( .A(n1843), .Z(n2468) );
  CLKBUF_X1 U8346 ( .A(n1863), .Z(n2456) );
  CLKBUF_X1 U8347 ( .A(n1861), .Z(n2450) );
  CLKBUF_X1 U8348 ( .A(n1837), .Z(n2462) );
  CLKBUF_X1 U8349 ( .A(n1853), .Z(n2402) );
  CLKBUF_X1 U8350 ( .A(n1845), .Z(n2432) );
  CLKBUF_X1 U8351 ( .A(n1832), .Z(n2426) );
  CLKBUF_X1 U8352 ( .A(n1846), .Z(n2420) );
  CLKBUF_X1 U8353 ( .A(n1874), .Z(n2440) );
  CLKBUF_X1 U8354 ( .A(n1875), .Z(n2404) );
  CLKBUF_X1 U8355 ( .A(n1876), .Z(n2380) );
  BUF_X2 U8356 ( .A(n1849), .Z(n2823) );
  BUF_X2 U8357 ( .A(n1850), .Z(n2817) );
  BUF_X2 U8358 ( .A(n1848), .Z(n2829) );
  BUF_X2 U8359 ( .A(n1851), .Z(n2811) );
  CLKBUF_X1 U8360 ( .A(n1867), .Z(n2832) );
  CLKBUF_X1 U8361 ( .A(n1852), .Z(n2851) );
  CLKBUF_X1 U8362 ( .A(n1869), .Z(n2844) );
  CLKBUF_X1 U8363 ( .A(n1870), .Z(n2838) );
  CLKBUF_X1 U8364 ( .A(n1878), .Z(n2778) );
  CLKBUF_X1 U8365 ( .A(n1866), .Z(n2790) );
  CLKBUF_X1 U8366 ( .A(n1866), .Z(n2791) );
  CLKBUF_X1 U8367 ( .A(n1872), .Z(n2797) );
  CLKBUF_X1 U8368 ( .A(n1871), .Z(n2803) );
  CLKBUF_X1 U8369 ( .A(n1851), .Z(n2809) );
  CLKBUF_X1 U8370 ( .A(n1850), .Z(n2815) );
  CLKBUF_X1 U8371 ( .A(n1849), .Z(n2821) );
  CLKBUF_X1 U8372 ( .A(n1848), .Z(n2827) );
  CLKBUF_X1 U8373 ( .A(n1867), .Z(n2833) );
  CLKBUF_X1 U8374 ( .A(n1870), .Z(n2839) );
  CLKBUF_X1 U8375 ( .A(n1877), .Z(n2784) );
  CLKBUF_X1 U8376 ( .A(n1872), .Z(n2796) );
  CLKBUF_X1 U8377 ( .A(n1871), .Z(n2802) );
  CLKBUF_X1 U8378 ( .A(n1851), .Z(n2808) );
  CLKBUF_X1 U8379 ( .A(n1850), .Z(n2814) );
  CLKBUF_X1 U8380 ( .A(n1849), .Z(n2820) );
  CLKBUF_X1 U8381 ( .A(n1848), .Z(n2826) );
  CLKBUF_X1 U8382 ( .A(n1881), .Z(n2693) );
  XNOR2_X1 U8383 ( .A(n2347), .B(n2346), .ZN(n946) );
  NAND2_X1 U8384 ( .A1(reg_mid_0[22]), .A2(reg_mid_1[38]), .ZN(n2346) );
  NOR2_X1 U8385 ( .A1(n649), .A2(n636), .ZN(n1608) );
  INV_X1 U8386 ( .A(n1300), .ZN(n645) );
  INV_X1 U8387 ( .A(n1622), .ZN(n622) );
  INV_X1 U8388 ( .A(n1604), .ZN(n647) );
  AND2_X1 U8389 ( .A1(n601), .A2(n603), .ZN(n2348) );
  INV_X1 U8390 ( .A(n1594), .ZN(n648) );
  INV_X1 U8391 ( .A(n1519), .ZN(n593) );
  INV_X1 U8392 ( .A(n1507), .ZN(n596) );
  INV_X1 U8393 ( .A(n1563), .ZN(n580) );
  INV_X1 U8394 ( .A(n1572), .ZN(n584) );
  INV_X1 U8395 ( .A(n1498), .ZN(n597) );
  AOI21_X1 U8396 ( .B1(n607), .B2(n1625), .A(n608), .ZN(n1623) );
  INV_X1 U8397 ( .A(n1619), .ZN(n608) );
  AOI21_X1 U8398 ( .B1(n601), .B2(n2365), .A(n602), .ZN(n1480) );
  OAI21_X1 U8399 ( .B1(n1521), .B2(n1532), .A(n1525), .ZN(n1528) );
  OAI21_X1 U8400 ( .B1(n1563), .B2(n1576), .A(n1566), .ZN(n1571) );
  OAI21_X1 U8401 ( .B1(n1467), .B2(n1480), .A(n1470), .ZN(n1475) );
  NAND2_X1 U8402 ( .A1(n1566), .A2(n580), .ZN(n1577) );
  AOI21_X1 U8403 ( .B1(n636), .B2(n649), .A(n1608), .ZN(n1621) );
  OAI21_X1 U8404 ( .B1(n1622), .B2(n1623), .A(n1617), .ZN(n1620) );
  NOR2_X1 U8405 ( .A1(n596), .A2(n1498), .ZN(n1509) );
  NOR2_X1 U8406 ( .A1(n647), .A2(n1594), .ZN(n1605) );
  NAND2_X1 U8407 ( .A1(n622), .A2(n1617), .ZN(n1624) );
  NAND2_X1 U8408 ( .A1(n1470), .A2(n603), .ZN(n1481) );
  NAND2_X1 U8409 ( .A1(n1525), .A2(n592), .ZN(n1533) );
  INV_X1 U8410 ( .A(n1521), .ZN(n592) );
  NOR2_X1 U8411 ( .A1(n1466), .A2(n1476), .ZN(n1477) );
  NOR2_X1 U8412 ( .A1(n1562), .A2(n1572), .ZN(n1573) );
  NOR2_X1 U8413 ( .A1(n1523), .A2(n1519), .ZN(n1529) );
  INV_X1 U8414 ( .A(n2178), .ZN(n607) );
  XNOR2_X1 U8415 ( .A(n1628), .B(n1625), .ZN(N195) );
  NAND2_X1 U8416 ( .A1(n1619), .A2(n607), .ZN(n1628) );
  INV_X1 U8417 ( .A(n1476), .ZN(n604) );
  OAI21_X1 U8418 ( .B1(n1720), .B2(n1721), .A(n1722), .ZN(n1714) );
  OAI21_X1 U8419 ( .B1(n1194), .B2(n1195), .A(n1196), .ZN(n1188) );
  INV_X1 U8420 ( .A(n1775), .ZN(n413) );
  INV_X1 U8421 ( .A(n1249), .ZN(n507) );
  INV_X1 U8422 ( .A(n1275), .ZN(n513) );
  INV_X1 U8423 ( .A(n1785), .ZN(n420) );
  INV_X1 U8424 ( .A(n1750), .ZN(n409) );
  INV_X1 U8425 ( .A(n1224), .ZN(n503) );
  AOI21_X1 U8426 ( .B1(n1258), .B2(n514), .A(n1275), .ZN(n1270) );
  AOI21_X1 U8427 ( .B1(n1739), .B2(n1740), .A(n1750), .ZN(n1748) );
  AOI21_X1 U8428 ( .B1(n1213), .B2(n1214), .A(n1224), .ZN(n1222) );
  AOI21_X1 U8429 ( .B1(n418), .B2(n1100), .A(n419), .ZN(n1793) );
  AOI21_X1 U8430 ( .B1(n1759), .B2(n1775), .A(n1767), .ZN(n1773) );
  AOI21_X1 U8431 ( .B1(n1233), .B2(n1249), .A(n1241), .ZN(n1247) );
  XNOR2_X1 U8432 ( .A(n1740), .B(n2349), .ZN(N106) );
  NAND2_X1 U8433 ( .A1(n1739), .A2(n409), .ZN(n2349) );
  XNOR2_X1 U8434 ( .A(n1214), .B(n2350), .ZN(N42) );
  NAND2_X1 U8435 ( .A1(n1213), .A2(n503), .ZN(n2350) );
  NOR2_X1 U8436 ( .A1(n413), .A2(n1767), .ZN(n1777) );
  NOR2_X1 U8437 ( .A1(n507), .A2(n1241), .ZN(n1251) );
  XNOR2_X1 U8438 ( .A(n1720), .B(n1723), .ZN(N111) );
  NOR2_X1 U8439 ( .A1(n1721), .A2(n404), .ZN(n1723) );
  INV_X1 U8440 ( .A(n1722), .ZN(n404) );
  XNOR2_X1 U8441 ( .A(n1194), .B(n1197), .ZN(N47) );
  NOR2_X1 U8442 ( .A1(n1195), .A2(n498), .ZN(n1197) );
  INV_X1 U8443 ( .A(n1196), .ZN(n498) );
  INV_X1 U8444 ( .A(n1293), .ZN(n650) );
  AOI21_X1 U8445 ( .B1(n1591), .B2(n654), .A(n1592), .ZN(n1584) );
  OAI21_X1 U8446 ( .B1(n1590), .B2(n648), .A(n1593), .ZN(n1591) );
  INV_X1 U8447 ( .A(n1314), .ZN(n643) );
  INV_X1 U8448 ( .A(n1544), .ZN(n588) );
  INV_X1 U8449 ( .A(n1517), .ZN(n595) );
  AOI21_X1 U8450 ( .B1(n1522), .B2(n593), .A(n1523), .ZN(n1512) );
  INV_X1 U8451 ( .A(n1617), .ZN(n623) );
  INV_X1 U8452 ( .A(n1318), .ZN(n642) );
  INV_X1 U8453 ( .A(n1297), .ZN(n646) );
  INV_X1 U8454 ( .A(n1357), .ZN(n633) );
  INV_X1 U8455 ( .A(n1448), .ZN(n610) );
  INV_X1 U8456 ( .A(n1347), .ZN(n635) );
  INV_X1 U8457 ( .A(n1337), .ZN(n638) );
  INV_X1 U8458 ( .A(n1367), .ZN(n631) );
  INV_X1 U8459 ( .A(n1306), .ZN(n644) );
  INV_X1 U8460 ( .A(n1554), .ZN(n586) );
  INV_X1 U8461 ( .A(n1458), .ZN(n606) );
  NOR2_X1 U8462 ( .A1(n1606), .A2(n1607), .ZN(n1594) );
  AOI21_X1 U8463 ( .B1(n1495), .B2(n599), .A(n1496), .ZN(n1488) );
  OAI21_X1 U8464 ( .B1(n1494), .B2(n597), .A(n1497), .ZN(n1495) );
  OAI21_X1 U8465 ( .B1(n1539), .B2(n1538), .A(n1540), .ZN(n1516) );
  NOR2_X1 U8466 ( .A1(n1626), .A2(n2287), .ZN(n1622) );
  NOR3_X1 U8467 ( .A1(n1589), .A2(n647), .A3(n1590), .ZN(n1588) );
  INV_X1 U8468 ( .A(n1472), .ZN(n605) );
  INV_X1 U8469 ( .A(n1568), .ZN(n585) );
  OAI21_X1 U8470 ( .B1(n1291), .B2(n1292), .A(n1293), .ZN(n1294) );
  OAI21_X1 U8471 ( .B1(n1312), .B2(n1313), .A(n1314), .ZN(n1315) );
  NAND2_X1 U8472 ( .A1(n2287), .A2(n1626), .ZN(n1617) );
  NAND2_X1 U8473 ( .A1(n621), .A2(n2353), .ZN(n1619) );
  OAI21_X1 U8474 ( .B1(n2131), .B2(n1618), .A(n1619), .ZN(n1616) );
  NAND2_X1 U8475 ( .A1(n1632), .A2(n1633), .ZN(n1613) );
  INV_X1 U8476 ( .A(n1589), .ZN(n654) );
  NAND2_X1 U8477 ( .A1(n1607), .A2(n1606), .ZN(n1604) );
  INV_X1 U8478 ( .A(n1610), .ZN(n649) );
  INV_X1 U8479 ( .A(n1438), .ZN(n2379) );
  INV_X1 U8480 ( .A(n1611), .ZN(n636) );
  AOI21_X1 U8481 ( .B1(n1377), .B2(n629), .A(n1378), .ZN(n1372) );
  INV_X1 U8482 ( .A(n1583), .ZN(n583) );
  OAI21_X1 U8483 ( .B1(n1424), .B2(n1433), .A(n1426), .ZN(n1430) );
  NOR2_X1 U8484 ( .A1(n1510), .A2(n1511), .ZN(n1498) );
  OAI21_X1 U8485 ( .B1(n1379), .B2(n1389), .A(n1381), .ZN(n1384) );
  OAI21_X1 U8486 ( .B1(n1400), .B2(n1412), .A(n1403), .ZN(n1407) );
  NOR3_X1 U8487 ( .A1(n1493), .A2(n596), .A3(n1494), .ZN(n1492) );
  NOR3_X1 U8488 ( .A1(n1519), .A2(n1520), .A3(n1521), .ZN(n1518) );
  NOR2_X1 U8489 ( .A1(n612), .A2(n1438), .ZN(n1440) );
  NAND2_X1 U8490 ( .A1(n632), .A2(n1363), .ZN(n1364) );
  INV_X1 U8491 ( .A(n1361), .ZN(n632) );
  NAND2_X1 U8492 ( .A1(n628), .A2(n1381), .ZN(n1390) );
  NAND2_X1 U8493 ( .A1(n619), .A2(n1403), .ZN(n1413) );
  NAND2_X1 U8494 ( .A1(n625), .A2(n1397), .ZN(n1405) );
  AOI21_X1 U8495 ( .B1(n1407), .B2(n620), .A(n1399), .ZN(n1406) );
  INV_X1 U8496 ( .A(n1395), .ZN(n625) );
  NAND2_X1 U8497 ( .A1(n637), .A2(n1343), .ZN(n1344) );
  INV_X1 U8498 ( .A(n1341), .ZN(n637) );
  NAND2_X1 U8499 ( .A1(n634), .A2(n1353), .ZN(n1354) );
  INV_X1 U8500 ( .A(n1351), .ZN(n634) );
  NAND2_X1 U8501 ( .A1(n630), .A2(n1375), .ZN(n1382) );
  AOI21_X1 U8502 ( .B1(n1384), .B2(n629), .A(n1378), .ZN(n1383) );
  NAND2_X1 U8503 ( .A1(n611), .A2(n1444), .ZN(n1445) );
  INV_X1 U8504 ( .A(n1442), .ZN(n611) );
  NOR2_X1 U8505 ( .A1(n1336), .A2(n1337), .ZN(n1339) );
  NOR2_X1 U8506 ( .A1(n1346), .A2(n1347), .ZN(n1349) );
  NOR2_X1 U8507 ( .A1(n1356), .A2(n1357), .ZN(n1359) );
  NOR2_X1 U8508 ( .A1(n1378), .A2(n1385), .ZN(n1387) );
  NOR2_X1 U8509 ( .A1(n1366), .A2(n1367), .ZN(n1369) );
  NOR2_X1 U8510 ( .A1(n627), .A2(n1391), .ZN(n1393) );
  NOR2_X1 U8511 ( .A1(n1399), .A2(n1408), .ZN(n1410) );
  NOR2_X1 U8512 ( .A1(n618), .A2(n1414), .ZN(n1416) );
  OAI21_X1 U8513 ( .B1(n1521), .B2(n1524), .A(n1525), .ZN(n1522) );
  NAND2_X1 U8514 ( .A1(n1535), .A2(n1534), .ZN(n1525) );
  AND2_X1 U8515 ( .A1(n1531), .A2(n1530), .ZN(n1523) );
  NAND2_X1 U8516 ( .A1(n1513), .A2(n1514), .ZN(n1517) );
  NAND2_X1 U8517 ( .A1(n1580), .A2(n1579), .ZN(n1566) );
  NAND2_X1 U8518 ( .A1(n1484), .A2(n1483), .ZN(n1470) );
  AND2_X1 U8519 ( .A1(n1575), .A2(n1574), .ZN(n1562) );
  XNOR2_X1 U8520 ( .A(n1432), .B(n1430), .ZN(N228) );
  NAND2_X1 U8521 ( .A1(n615), .A2(n1431), .ZN(n1432) );
  NAND2_X1 U8522 ( .A1(n1558), .A2(n1559), .ZN(n1568) );
  XOR2_X1 U8523 ( .A(n1433), .B(n2351), .Z(N227) );
  NAND2_X1 U8524 ( .A1(n613), .A2(n1426), .ZN(n2351) );
  AOI21_X1 U8525 ( .B1(n615), .B2(n1430), .A(n614), .ZN(n1427) );
  INV_X1 U8526 ( .A(n1493), .ZN(n599) );
  NAND2_X1 U8527 ( .A1(n1511), .A2(n1510), .ZN(n1507) );
  INV_X1 U8528 ( .A(n1487), .ZN(n600) );
  INV_X1 U8529 ( .A(n1578), .ZN(n582) );
  INV_X1 U8530 ( .A(n1520), .ZN(n590) );
  OAI21_X1 U8531 ( .B1(n1590), .B2(n1601), .A(n1593), .ZN(n1598) );
  OAI21_X1 U8532 ( .B1(n1494), .B2(n1505), .A(n1497), .ZN(n1501) );
  AOI21_X1 U8533 ( .B1(n654), .B2(n1598), .A(n1592), .ZN(n1595) );
  AOI21_X1 U8534 ( .B1(n1423), .B2(n615), .A(n614), .ZN(n1418) );
  OAI21_X1 U8535 ( .B1(n1424), .B2(n1425), .A(n1426), .ZN(n1423) );
  NOR2_X1 U8536 ( .A1(n1307), .A2(n1308), .ZN(n1300) );
  OAI21_X1 U8537 ( .B1(n1462), .B2(n1463), .A(n1472), .ZN(n1473) );
  AOI21_X1 U8538 ( .B1(n1475), .B2(n604), .A(n1466), .ZN(n1474) );
  OAI21_X1 U8539 ( .B1(n1513), .B2(n1514), .A(n1517), .ZN(n1526) );
  AOI21_X1 U8540 ( .B1(n1528), .B2(n593), .A(n1523), .ZN(n1527) );
  OAI21_X1 U8541 ( .B1(n1558), .B2(n1559), .A(n1568), .ZN(n1569) );
  AOI21_X1 U8542 ( .B1(n1571), .B2(n584), .A(n1562), .ZN(n1570) );
  NAND2_X1 U8543 ( .A1(n598), .A2(n1497), .ZN(n1506) );
  INV_X1 U8544 ( .A(n1494), .ZN(n598) );
  NAND2_X1 U8545 ( .A1(n589), .A2(n1540), .ZN(n1541) );
  INV_X1 U8546 ( .A(n1538), .ZN(n589) );
  NAND2_X1 U8547 ( .A1(n609), .A2(n1454), .ZN(n1455) );
  INV_X1 U8548 ( .A(n1452), .ZN(n609) );
  NAND2_X1 U8549 ( .A1(n600), .A2(n1489), .ZN(n1499) );
  AOI21_X1 U8550 ( .B1(n1501), .B2(n599), .A(n1496), .ZN(n1500) );
  NAND2_X1 U8551 ( .A1(n587), .A2(n1550), .ZN(n1551) );
  INV_X1 U8552 ( .A(n1548), .ZN(n587) );
  NOR2_X1 U8553 ( .A1(n602), .A2(n1482), .ZN(n1485) );
  NOR2_X1 U8554 ( .A1(n1448), .A2(n1447), .ZN(n1450) );
  NOR2_X1 U8555 ( .A1(n1458), .A2(n1457), .ZN(n1460) );
  NOR2_X1 U8556 ( .A1(n1544), .A2(n1543), .ZN(n1546) );
  NOR2_X1 U8557 ( .A1(n1554), .A2(n1553), .ZN(n1556) );
  NOR2_X1 U8558 ( .A1(n581), .A2(n1578), .ZN(n1581) );
  NOR2_X1 U8559 ( .A1(n1493), .A2(n1496), .ZN(n1503) );
  NOR2_X1 U8560 ( .A1(n1589), .A2(n1592), .ZN(n1599) );
  NOR2_X1 U8561 ( .A1(n591), .A2(n1520), .ZN(n1536) );
  OAI21_X1 U8562 ( .B1(n1379), .B2(n1380), .A(n1381), .ZN(n1377) );
  XNOR2_X1 U8563 ( .A(n1601), .B(n1602), .ZN(N199) );
  NOR2_X1 U8564 ( .A1(n653), .A2(n1590), .ZN(n1602) );
  INV_X1 U8565 ( .A(n1593), .ZN(n653) );
  NAND2_X1 U8566 ( .A1(n1312), .A2(n1313), .ZN(n1314) );
  NAND2_X1 U8567 ( .A1(n1462), .A2(n1463), .ZN(n1472) );
  INV_X1 U8568 ( .A(n1385), .ZN(n629) );
  INV_X1 U8569 ( .A(n1431), .ZN(n614) );
  INV_X1 U8570 ( .A(n1468), .ZN(n602) );
  INV_X1 U8571 ( .A(n1425), .ZN(n612) );
  INV_X1 U8572 ( .A(n1380), .ZN(n627) );
  INV_X1 U8573 ( .A(n1524), .ZN(n591) );
  INV_X1 U8574 ( .A(n1401), .ZN(n618) );
  INV_X1 U8575 ( .A(n1564), .ZN(n581) );
  INV_X1 U8576 ( .A(n1379), .ZN(n628) );
  INV_X1 U8577 ( .A(n1408), .ZN(n620) );
  INV_X1 U8578 ( .A(n1400), .ZN(n619) );
  INV_X1 U8579 ( .A(n1424), .ZN(n613) );
  INV_X1 U8580 ( .A(n1371), .ZN(n630) );
  INV_X1 U8581 ( .A(n1391), .ZN(n626) );
  INV_X1 U8582 ( .A(n1419), .ZN(n616) );
  INV_X1 U8583 ( .A(n1414), .ZN(n617) );
  NAND2_X1 U8584 ( .A1(n1291), .A2(n1292), .ZN(n1293) );
  NAND2_X1 U8585 ( .A1(n1308), .A2(n1307), .ZN(n1302) );
  OAI221_X1 U8586 ( .B1(n410), .B2(n1755), .C1(n1756), .C2(n1757), .A(n1758), 
        .ZN(n1740) );
  INV_X1 U8587 ( .A(n1760), .ZN(n410) );
  AOI21_X1 U8588 ( .B1(n1764), .B2(n411), .A(n1765), .ZN(n1755) );
  OAI221_X1 U8589 ( .B1(n504), .B2(n1229), .C1(n1230), .C2(n1231), .A(n1232), 
        .ZN(n1214) );
  INV_X1 U8590 ( .A(n1234), .ZN(n504) );
  AOI21_X1 U8591 ( .B1(n1238), .B2(n505), .A(n1239), .ZN(n1229) );
  NOR2_X1 U8592 ( .A1(n1778), .A2(n1779), .ZN(n1767) );
  NOR2_X1 U8593 ( .A1(n1252), .A2(n1253), .ZN(n1241) );
  OAI211_X1 U8594 ( .C1(n1780), .C2(n1781), .A(n1782), .B(n1783), .ZN(n1759)
         );
  AOI21_X1 U8595 ( .B1(n1786), .B2(n417), .A(n416), .ZN(n1781) );
  NAND4_X1 U8596 ( .A1(n420), .A2(n418), .A3(n417), .A4(n1784), .ZN(n1783) );
  INV_X1 U8597 ( .A(n1787), .ZN(n416) );
  OAI211_X1 U8598 ( .C1(n1254), .C2(n1255), .A(n1256), .B(n1257), .ZN(n1233)
         );
  NAND4_X1 U8599 ( .A1(n512), .A2(n1258), .A3(n511), .A4(n1259), .ZN(n1257) );
  AOI21_X1 U8600 ( .B1(n1261), .B2(n511), .A(n510), .ZN(n1255) );
  NOR2_X1 U8601 ( .A1(n1254), .A2(n1260), .ZN(n1259) );
  AOI21_X1 U8602 ( .B1(n1726), .B2(n405), .A(n1727), .ZN(n1720) );
  INV_X1 U8603 ( .A(n1728), .ZN(n405) );
  AOI21_X1 U8604 ( .B1(n1200), .B2(n499), .A(n1201), .ZN(n1194) );
  INV_X1 U8605 ( .A(n1202), .ZN(n499) );
  AOI21_X1 U8606 ( .B1(n1688), .B2(n1689), .A(n1690), .ZN(n1683) );
  NAND2_X1 U8607 ( .A1(n1691), .A2(n1692), .ZN(n1688) );
  AOI21_X1 U8608 ( .B1(n1162), .B2(n1163), .A(n1164), .ZN(n1157) );
  NAND2_X1 U8609 ( .A1(n1165), .A2(n1166), .ZN(n1162) );
  AOI21_X1 U8610 ( .B1(n1705), .B2(n401), .A(n1706), .ZN(n1700) );
  INV_X1 U8611 ( .A(n1707), .ZN(n401) );
  AOI21_X1 U8612 ( .B1(n1179), .B2(n495), .A(n1180), .ZN(n1174) );
  INV_X1 U8613 ( .A(n1181), .ZN(n495) );
  AOI21_X1 U8614 ( .B1(n403), .B2(n1714), .A(n1715), .ZN(n1710) );
  INV_X1 U8615 ( .A(n1716), .ZN(n403) );
  AOI21_X1 U8616 ( .B1(n497), .B2(n1188), .A(n1189), .ZN(n1184) );
  INV_X1 U8617 ( .A(n1190), .ZN(n497) );
  AOI21_X1 U8618 ( .B1(n1676), .B2(n1677), .A(n1678), .ZN(n1671) );
  NAND2_X1 U8619 ( .A1(n1679), .A2(n1680), .ZN(n1676) );
  AOI21_X1 U8620 ( .B1(n1150), .B2(n1151), .A(n1152), .ZN(n1145) );
  NAND2_X1 U8621 ( .A1(n1153), .A2(n1154), .ZN(n1150) );
  OAI21_X1 U8622 ( .B1(n400), .B2(n1694), .A(n1695), .ZN(n1689) );
  INV_X1 U8623 ( .A(n1696), .ZN(n400) );
  OAI21_X1 U8624 ( .B1(n494), .B2(n1168), .A(n1169), .ZN(n1163) );
  INV_X1 U8625 ( .A(n1170), .ZN(n494) );
  OAI21_X1 U8626 ( .B1(n1683), .B2(n1684), .A(n1685), .ZN(n1677) );
  OAI21_X1 U8627 ( .B1(n1157), .B2(n1158), .A(n1159), .ZN(n1151) );
  OAI21_X1 U8628 ( .B1(n1699), .B2(n1700), .A(n1701), .ZN(n1696) );
  NOR2_X1 U8629 ( .A1(n1702), .A2(n1703), .ZN(n1699) );
  OAI21_X1 U8630 ( .B1(n1173), .B2(n1174), .A(n1175), .ZN(n1170) );
  NOR2_X1 U8631 ( .A1(n1176), .A2(n1177), .ZN(n1173) );
  OAI21_X1 U8632 ( .B1(n1710), .B2(n1711), .A(n1712), .ZN(n1705) );
  OAI21_X1 U8633 ( .B1(n1184), .B2(n1185), .A(n1186), .ZN(n1179) );
  OAI21_X1 U8634 ( .B1(n1731), .B2(n1732), .A(n1733), .ZN(n1726) );
  AOI21_X1 U8635 ( .B1(n1734), .B2(n407), .A(n1735), .ZN(n1732) );
  OAI211_X1 U8636 ( .C1(n1736), .C2(n409), .A(n1737), .B(n1738), .ZN(n1734) );
  OAI21_X1 U8637 ( .B1(n1205), .B2(n1206), .A(n1207), .ZN(n1200) );
  AOI21_X1 U8638 ( .B1(n1208), .B2(n501), .A(n1209), .ZN(n1206) );
  OAI211_X1 U8639 ( .C1(n1210), .C2(n503), .A(n1211), .B(n1212), .ZN(n1208) );
  NOR2_X1 U8640 ( .A1(n1797), .A2(n1796), .ZN(n1785) );
  NOR2_X1 U8641 ( .A1(n1753), .A2(n1754), .ZN(n1750) );
  NOR2_X1 U8642 ( .A1(n1227), .A2(n1228), .ZN(n1224) );
  NOR2_X1 U8643 ( .A1(n1278), .A2(n1277), .ZN(n1275) );
  NOR2_X1 U8644 ( .A1(n1640), .A2(n1641), .ZN(n1635) );
  AOI21_X1 U8645 ( .B1(n1642), .B2(n1643), .A(n395), .ZN(n1640) );
  NOR2_X1 U8646 ( .A1(n1114), .A2(n1115), .ZN(n1109) );
  AOI21_X1 U8647 ( .B1(n1116), .B2(n1117), .A(n489), .ZN(n1114) );
  NOR3_X1 U8648 ( .A1(n1762), .A2(n413), .A3(n1763), .ZN(n1761) );
  NOR3_X1 U8649 ( .A1(n1236), .A2(n507), .A3(n1237), .ZN(n1235) );
  NOR2_X1 U8650 ( .A1(n1664), .A2(n1665), .ZN(n1659) );
  AOI21_X1 U8651 ( .B1(n1666), .B2(n1667), .A(n397), .ZN(n1664) );
  NOR2_X1 U8652 ( .A1(n1138), .A2(n1139), .ZN(n1133) );
  AOI21_X1 U8653 ( .B1(n1140), .B2(n1141), .A(n491), .ZN(n1138) );
  NOR2_X1 U8654 ( .A1(n1652), .A2(n1653), .ZN(n1647) );
  AOI21_X1 U8655 ( .B1(n1654), .B2(n1655), .A(n396), .ZN(n1652) );
  NOR2_X1 U8656 ( .A1(n1126), .A2(n1127), .ZN(n1121) );
  AOI21_X1 U8657 ( .B1(n1128), .B2(n1129), .A(n490), .ZN(n1126) );
  NOR2_X1 U8658 ( .A1(n1780), .A2(n1103), .ZN(n1784) );
  OAI21_X1 U8659 ( .B1(n1763), .B2(n414), .A(n1766), .ZN(n1764) );
  INV_X1 U8660 ( .A(n1767), .ZN(n414) );
  OAI21_X1 U8661 ( .B1(n1237), .B2(n508), .A(n1240), .ZN(n1238) );
  INV_X1 U8662 ( .A(n1241), .ZN(n508) );
  NAND2_X1 U8663 ( .A1(n1796), .A2(n1797), .ZN(n1105) );
  OAI21_X1 U8664 ( .B1(n1102), .B2(n1105), .A(n1788), .ZN(n1786) );
  OAI21_X1 U8665 ( .B1(n1262), .B2(n513), .A(n1263), .ZN(n1261) );
  NAND2_X1 U8666 ( .A1(n1277), .A2(n1278), .ZN(n1258) );
  NAND2_X1 U8667 ( .A1(n1756), .A2(n1757), .ZN(n1760) );
  NAND2_X1 U8668 ( .A1(n1230), .A2(n1231), .ZN(n1234) );
  INV_X1 U8669 ( .A(n1792), .ZN(n417) );
  XNOR2_X1 U8670 ( .A(n397), .B(n1669), .ZN(N121) );
  AOI21_X1 U8671 ( .B1(n1667), .B2(n1666), .A(n1665), .ZN(n1669) );
  XNOR2_X1 U8672 ( .A(n396), .B(n1657), .ZN(N123) );
  AOI21_X1 U8673 ( .B1(n1655), .B2(n1654), .A(n1653), .ZN(n1657) );
  XNOR2_X1 U8674 ( .A(n395), .B(n1645), .ZN(N125) );
  AOI21_X1 U8675 ( .B1(n1643), .B2(n1642), .A(n1641), .ZN(n1645) );
  XNOR2_X1 U8676 ( .A(n491), .B(n1143), .ZN(N57) );
  AOI21_X1 U8677 ( .B1(n1141), .B2(n1140), .A(n1139), .ZN(n1143) );
  XNOR2_X1 U8678 ( .A(n490), .B(n1131), .ZN(N59) );
  AOI21_X1 U8679 ( .B1(n1129), .B2(n1128), .A(n1127), .ZN(n1131) );
  XNOR2_X1 U8680 ( .A(n489), .B(n1119), .ZN(N61) );
  AOI21_X1 U8681 ( .B1(n1117), .B2(n1116), .A(n1115), .ZN(n1119) );
  NAND2_X1 U8682 ( .A1(n1754), .A2(n1753), .ZN(n1739) );
  NAND2_X1 U8683 ( .A1(n1228), .A2(n1227), .ZN(n1213) );
  NAND2_X1 U8684 ( .A1(n1779), .A2(n1778), .ZN(n1775) );
  NAND2_X1 U8685 ( .A1(n1253), .A2(n1252), .ZN(n1249) );
  INV_X1 U8686 ( .A(n1268), .ZN(n510) );
  INV_X1 U8687 ( .A(n1762), .ZN(n411) );
  INV_X1 U8688 ( .A(n1236), .ZN(n505) );
  INV_X1 U8689 ( .A(n1102), .ZN(n418) );
  INV_X1 U8690 ( .A(n1744), .ZN(n407) );
  INV_X1 U8691 ( .A(n1218), .ZN(n501) );
  INV_X1 U8692 ( .A(n1262), .ZN(n512) );
  INV_X1 U8693 ( .A(n1736), .ZN(n408) );
  INV_X1 U8694 ( .A(n1210), .ZN(n502) );
  OAI21_X1 U8695 ( .B1(n1262), .B2(n1270), .A(n1263), .ZN(n1267) );
  OAI21_X1 U8696 ( .B1(n1785), .B2(n1103), .A(n1105), .ZN(n1100) );
  OAI21_X1 U8697 ( .B1(n1763), .B2(n1773), .A(n1766), .ZN(n1770) );
  OAI21_X1 U8698 ( .B1(n1237), .B2(n1247), .A(n1240), .ZN(n1244) );
  NOR2_X1 U8699 ( .A1(n1725), .A2(n1724), .ZN(n1721) );
  NOR2_X1 U8700 ( .A1(n1199), .A2(n1198), .ZN(n1195) );
  OAI21_X1 U8701 ( .B1(n1736), .B2(n1748), .A(n1738), .ZN(n1743) );
  OAI21_X1 U8702 ( .B1(n1210), .B2(n1222), .A(n1212), .ZN(n1217) );
  NOR2_X1 U8703 ( .A1(n1679), .A2(n1680), .ZN(n1678) );
  NOR2_X1 U8704 ( .A1(n1153), .A2(n1154), .ZN(n1152) );
  NOR2_X1 U8705 ( .A1(n1691), .A2(n1692), .ZN(n1690) );
  NOR2_X1 U8706 ( .A1(n1165), .A2(n1166), .ZN(n1164) );
  XNOR2_X1 U8707 ( .A(n1264), .B(n1265), .ZN(N37) );
  NOR2_X1 U8708 ( .A1(n509), .A2(n1254), .ZN(n1265) );
  AOI21_X1 U8709 ( .B1(n511), .B2(n1267), .A(n510), .ZN(n1264) );
  INV_X1 U8710 ( .A(n1256), .ZN(n509) );
  NAND2_X1 U8711 ( .A1(n513), .A2(n1258), .ZN(n1276) );
  NOR2_X1 U8712 ( .A1(n415), .A2(n1780), .ZN(n1790) );
  OAI21_X1 U8713 ( .B1(n1792), .B2(n1793), .A(n1787), .ZN(n1789) );
  INV_X1 U8714 ( .A(n1782), .ZN(n415) );
  NAND2_X1 U8715 ( .A1(n412), .A2(n1766), .ZN(n1774) );
  INV_X1 U8716 ( .A(n1763), .ZN(n412) );
  NAND2_X1 U8717 ( .A1(n408), .A2(n1738), .ZN(n1749) );
  NAND2_X1 U8718 ( .A1(n506), .A2(n1240), .ZN(n1248) );
  INV_X1 U8719 ( .A(n1237), .ZN(n506) );
  NAND2_X1 U8720 ( .A1(n502), .A2(n1212), .ZN(n1223) );
  NAND2_X1 U8721 ( .A1(n1787), .A2(n417), .ZN(n1794) );
  NAND2_X1 U8722 ( .A1(n402), .A2(n1712), .ZN(n1713) );
  INV_X1 U8723 ( .A(n1711), .ZN(n402) );
  NAND2_X1 U8724 ( .A1(n496), .A2(n1186), .ZN(n1187) );
  INV_X1 U8725 ( .A(n1185), .ZN(n496) );
  OAI21_X1 U8726 ( .B1(n1702), .B2(n1703), .A(n1701), .ZN(n1704) );
  OAI21_X1 U8727 ( .B1(n1176), .B2(n1177), .A(n1175), .ZN(n1178) );
  NOR2_X1 U8728 ( .A1(n1744), .A2(n1735), .ZN(n1746) );
  NOR2_X1 U8729 ( .A1(n1728), .A2(n1727), .ZN(n1729) );
  NOR2_X1 U8730 ( .A1(n1716), .A2(n1715), .ZN(n1718) );
  NOR2_X1 U8731 ( .A1(n1707), .A2(n1706), .ZN(n1708) );
  NOR2_X1 U8732 ( .A1(n1694), .A2(n399), .ZN(n1697) );
  INV_X1 U8733 ( .A(n1695), .ZN(n399) );
  NOR2_X1 U8734 ( .A1(n1218), .A2(n1209), .ZN(n1220) );
  NOR2_X1 U8735 ( .A1(n1202), .A2(n1201), .ZN(n1203) );
  NOR2_X1 U8736 ( .A1(n1190), .A2(n1189), .ZN(n1192) );
  NOR2_X1 U8737 ( .A1(n1181), .A2(n1180), .ZN(n1182) );
  NOR2_X1 U8738 ( .A1(n1168), .A2(n493), .ZN(n1171) );
  INV_X1 U8739 ( .A(n1169), .ZN(n493) );
  NOR2_X1 U8740 ( .A1(n1762), .A2(n1765), .ZN(n1771) );
  NOR2_X1 U8741 ( .A1(n1236), .A2(n1239), .ZN(n1245) );
  NOR2_X1 U8742 ( .A1(n419), .A2(n1102), .ZN(n1101) );
  AOI21_X1 U8743 ( .B1(n1692), .B2(n1691), .A(n1690), .ZN(n1693) );
  AOI21_X1 U8744 ( .B1(n1680), .B2(n1679), .A(n1678), .ZN(n1682) );
  AOI21_X1 U8745 ( .B1(n1166), .B2(n1165), .A(n1164), .ZN(n1167) );
  AOI21_X1 U8746 ( .B1(n1154), .B2(n1153), .A(n1152), .ZN(n1156) );
  OAI21_X1 U8747 ( .B1(n1756), .B2(n1757), .A(n1760), .ZN(n1768) );
  AOI21_X1 U8748 ( .B1(n1770), .B2(n411), .A(n1765), .ZN(n1769) );
  NAND2_X1 U8749 ( .A1(n406), .A2(n1733), .ZN(n1741) );
  AOI21_X1 U8750 ( .B1(n1743), .B2(n407), .A(n1735), .ZN(n1742) );
  INV_X1 U8751 ( .A(n1731), .ZN(n406) );
  OAI21_X1 U8752 ( .B1(n1230), .B2(n1231), .A(n1234), .ZN(n1242) );
  AOI21_X1 U8753 ( .B1(n1244), .B2(n505), .A(n1239), .ZN(n1243) );
  NAND2_X1 U8754 ( .A1(n500), .A2(n1207), .ZN(n1215) );
  AOI21_X1 U8755 ( .B1(n1217), .B2(n501), .A(n1209), .ZN(n1216) );
  INV_X1 U8756 ( .A(n1205), .ZN(n500) );
  NAND2_X1 U8757 ( .A1(n1702), .A2(n1703), .ZN(n1701) );
  NAND2_X1 U8758 ( .A1(n1176), .A2(n1177), .ZN(n1175) );
  INV_X1 U8759 ( .A(n1260), .ZN(n514) );
  XNOR2_X1 U8760 ( .A(n1683), .B(n1686), .ZN(N118) );
  NOR2_X1 U8761 ( .A1(n1684), .A2(n398), .ZN(n1686) );
  INV_X1 U8762 ( .A(n1685), .ZN(n398) );
  XNOR2_X1 U8763 ( .A(n1157), .B(n1160), .ZN(N54) );
  NOR2_X1 U8764 ( .A1(n1158), .A2(n492), .ZN(n1160) );
  INV_X1 U8765 ( .A(n1159), .ZN(n492) );
  XOR2_X1 U8766 ( .A(n1270), .B(n2352), .Z(N35) );
  NAND2_X1 U8767 ( .A1(n1263), .A2(n512), .ZN(n2352) );
  NAND2_X1 U8768 ( .A1(n1724), .A2(n1725), .ZN(n1722) );
  NAND2_X1 U8769 ( .A1(n1198), .A2(n1199), .ZN(n1196) );
  XNOR2_X1 U8770 ( .A(n1269), .B(n1267), .ZN(N36) );
  NAND2_X1 U8771 ( .A1(n1268), .A2(n511), .ZN(n1269) );
  INV_X1 U8772 ( .A(n1788), .ZN(n419) );
  NAND2_X1 U8773 ( .A1(n420), .A2(n1105), .ZN(n1104) );
  NOR2_X1 U8774 ( .A1(n1666), .A2(n1667), .ZN(n1665) );
  NOR2_X1 U8775 ( .A1(n1140), .A2(n1141), .ZN(n1139) );
  NOR2_X1 U8776 ( .A1(n1654), .A2(n1655), .ZN(n1653) );
  NOR2_X1 U8777 ( .A1(n1128), .A2(n1129), .ZN(n1127) );
  NOR2_X1 U8778 ( .A1(n1642), .A2(n1643), .ZN(n1641) );
  NOR2_X1 U8779 ( .A1(n1116), .A2(n1117), .ZN(n1115) );
  INV_X1 U8780 ( .A(n1327), .ZN(n640) );
  XNOR2_X1 U8781 ( .A(\mult_22/CARRYB[63][6] ), .B(\mult_22/SUMB[63][7] ), 
        .ZN(n1607) );
  AOI21_X1 U8782 ( .B1(\mult_22/CARRYB[63][8] ), .B2(\mult_22/SUMB[63][9] ), 
        .A(n1597), .ZN(n1583) );
  XNOR2_X1 U8783 ( .A(\mult_22/CARRYB[63][5] ), .B(\mult_22/SUMB[63][6] ), 
        .ZN(n1610) );
  AND3_X1 U8784 ( .A1(\mult_22/CARRYB[63][7] ), .A2(n1600), .A3(
        \mult_22/SUMB[63][8] ), .ZN(n1592) );
  NAND2_X1 U8785 ( .A1(\mult_22/SUMB[63][6] ), .A2(\mult_22/CARRYB[63][5] ), 
        .ZN(n1606) );
  NAND2_X1 U8786 ( .A1(\mult_22/SUMB[63][4] ), .A2(\mult_22/CARRYB[63][3] ), 
        .ZN(n1627) );
  INV_X1 U8787 ( .A(\mult_22/CARRYB[25][34] ), .ZN(n698) );
  NAND2_X1 U8788 ( .A1(\mult_22/CARRYB[63][4] ), .A2(\mult_22/SUMB[63][5] ), 
        .ZN(n1611) );
  INV_X1 U8789 ( .A(\mult_22/CARRYB[23][32] ), .ZN(n703) );
  INV_X1 U8790 ( .A(\mult_22/CARRYB[27][30] ), .ZN(n693) );
  INV_X1 U8791 ( .A(n1630), .ZN(n621) );
  OAI21_X1 U8792 ( .B1(\mult_22/CARRYB[63][3] ), .B2(n2159), .A(n1627), .ZN(
        n1630) );
  INV_X1 U8793 ( .A(\mult_22/CARRYB[32][28] ), .ZN(n686) );
  INV_X1 U8794 ( .A(\mult_22/SUMB[20][37] ), .ZN(n713) );
  AND2_X1 U8795 ( .A1(\mult_22/SUMB[63][3] ), .A2(\mult_22/CARRYB[63][2] ), 
        .ZN(n2353) );
  INV_X1 U8796 ( .A(\mult_22/SUMB[21][39] ), .ZN(n709) );
  INV_X1 U8797 ( .A(\mult_22/SUMB[10][47] ), .ZN(n727) );
  XOR2_X1 U8798 ( .A(\mult_22/SUMB[63][3] ), .B(\mult_22/CARRYB[63][2] ), .Z(
        n2354) );
  AOI21_X1 U8799 ( .B1(\mult_22/CARRYB[63][22] ), .B2(\mult_22/SUMB[63][23] ), 
        .A(n1508), .ZN(n1494) );
  AOI21_X1 U8800 ( .B1(\mult_22/CARRYB[63][23] ), .B2(\mult_22/SUMB[63][24] ), 
        .A(n1504), .ZN(n1493) );
  XNOR2_X1 U8801 ( .A(\mult_22/CARRYB[63][13] ), .B(\mult_22/SUMB[63][14] ), 
        .ZN(n1558) );
  XNOR2_X1 U8802 ( .A(\mult_22/CARRYB[63][21] ), .B(\mult_22/SUMB[63][22] ), 
        .ZN(n1513) );
  AOI21_X1 U8803 ( .B1(\mult_22/CARRYB[63][13] ), .B2(\mult_22/SUMB[63][14] ), 
        .A(n1557), .ZN(n1554) );
  AOI21_X1 U8804 ( .B1(\mult_22/CARRYB[63][9] ), .B2(\mult_22/SUMB[63][10] ), 
        .A(n1582), .ZN(n1578) );
  AOI21_X1 U8805 ( .B1(\mult_22/CARRYB[63][15] ), .B2(\mult_22/SUMB[63][16] ), 
        .A(n1547), .ZN(n1544) );
  AOI21_X1 U8806 ( .B1(\mult_22/CARRYB[63][16] ), .B2(\mult_22/SUMB[63][17] ), 
        .A(n1545), .ZN(n1538) );
  XNOR2_X1 U8807 ( .A(\mult_22/CARRYB[63][22] ), .B(\mult_22/SUMB[63][23] ), 
        .ZN(n1511) );
  AOI21_X1 U8808 ( .B1(\mult_22/CARRYB[63][25] ), .B2(\mult_22/SUMB[63][26] ), 
        .A(n1486), .ZN(n1482) );
  AOI21_X1 U8809 ( .B1(\mult_22/CARRYB[63][14] ), .B2(\mult_22/SUMB[63][15] ), 
        .A(n1555), .ZN(n1548) );
  AOI21_X1 U8810 ( .B1(\mult_22/CARRYB[63][24] ), .B2(\mult_22/SUMB[63][25] ), 
        .A(n1502), .ZN(n1487) );
  INV_X1 U8811 ( .A(n1321), .ZN(n641) );
  INV_X1 U8812 ( .A(n1331), .ZN(n639) );
  AND3_X1 U8813 ( .A1(\mult_22/CARRYB[63][23] ), .A2(n1504), .A3(
        \mult_22/SUMB[63][24] ), .ZN(n1496) );
  NAND2_X1 U8814 ( .A1(\mult_22/CARRYB[63][20] ), .A2(\mult_22/SUMB[63][21] ), 
        .ZN(n1514) );
  NAND2_X1 U8815 ( .A1(\mult_22/SUMB[63][13] ), .A2(\mult_22/CARRYB[63][12] ), 
        .ZN(n1559) );
  NAND2_X1 U8816 ( .A1(\mult_22/SUMB[63][22] ), .A2(\mult_22/CARRYB[63][21] ), 
        .ZN(n1510) );
  AND3_X1 U8817 ( .A1(\mult_22/CARRYB[63][15] ), .A2(n1547), .A3(
        \mult_22/SUMB[63][16] ), .ZN(n1543) );
  AND3_X1 U8818 ( .A1(\mult_22/CARRYB[63][13] ), .A2(n1557), .A3(
        \mult_22/SUMB[63][14] ), .ZN(n1553) );
  AND2_X1 U8819 ( .A1(\mult_22/SUMB[63][11] ), .A2(\mult_22/CARRYB[63][10] ), 
        .ZN(n1580) );
  AND2_X1 U8820 ( .A1(\mult_22/SUMB[63][27] ), .A2(\mult_22/CARRYB[63][26] ), 
        .ZN(n1484) );
  AND2_X1 U8821 ( .A1(\mult_22/CARRYB[63][18] ), .A2(\mult_22/SUMB[63][19] ), 
        .ZN(n1535) );
  AND2_X1 U8822 ( .A1(\mult_22/SUMB[63][12] ), .A2(\mult_22/CARRYB[63][11] ), 
        .ZN(n1575) );
  AND2_X1 U8823 ( .A1(\mult_22/CARRYB[63][19] ), .A2(\mult_22/SUMB[63][20] ), 
        .ZN(n1531) );
  AOI21_X1 U8824 ( .B1(\mult_22/CARRYB[63][34] ), .B2(\mult_22/SUMB[63][35] ), 
        .A(n1437), .ZN(n1424) );
  XNOR2_X1 U8825 ( .A(\mult_22/CARRYB[63][57] ), .B(\mult_22/SUMB[63][58] ), 
        .ZN(n1312) );
  XNOR2_X1 U8826 ( .A(\mult_22/CARRYB[63][29] ), .B(\mult_22/SUMB[63][30] ), 
        .ZN(n1462) );
  AOI21_X1 U8827 ( .B1(\mult_22/CARRYB[63][36] ), .B2(\mult_22/SUMB[63][37] ), 
        .A(n1429), .ZN(n1419) );
  AOI21_X1 U8828 ( .B1(\mult_22/SUMB[63][58] ), .B2(\mult_22/CARRYB[63][57] ), 
        .A(n1310), .ZN(n1306) );
  AOI21_X1 U8829 ( .B1(\mult_22/CARRYB[63][29] ), .B2(\mult_22/SUMB[63][30] ), 
        .A(n1461), .ZN(n1458) );
  AOI21_X1 U8830 ( .B1(\mult_22/CARRYB[63][47] ), .B2(\mult_22/SUMB[63][48] ), 
        .A(n1360), .ZN(n1357) );
  AOI21_X1 U8831 ( .B1(\mult_22/CARRYB[63][43] ), .B2(\mult_22/SUMB[63][44] ), 
        .A(n1388), .ZN(n1385) );
  AOI21_X1 U8832 ( .B1(\mult_22/CARRYB[63][39] ), .B2(\mult_22/SUMB[63][40] ), 
        .A(n1411), .ZN(n1408) );
  AOI21_X1 U8833 ( .B1(\mult_22/CARRYB[63][45] ), .B2(\mult_22/SUMB[63][46] ), 
        .A(n1370), .ZN(n1367) );
  AOI21_X1 U8834 ( .B1(\mult_22/CARRYB[63][51] ), .B2(\mult_22/SUMB[63][52] ), 
        .A(n1340), .ZN(n1337) );
  AOI21_X1 U8835 ( .B1(\mult_22/CARRYB[63][55] ), .B2(\mult_22/SUMB[63][56] ), 
        .A(n1320), .ZN(n1318) );
  AOI21_X1 U8836 ( .B1(\mult_22/CARRYB[63][37] ), .B2(\mult_22/SUMB[63][38] ), 
        .A(n1417), .ZN(n1414) );
  AOI21_X1 U8837 ( .B1(\mult_22/CARRYB[63][41] ), .B2(\mult_22/SUMB[63][42] ), 
        .A(n1394), .ZN(n1391) );
  AOI21_X1 U8838 ( .B1(\mult_22/SUMB[63][50] ), .B2(\mult_22/CARRYB[63][49] ), 
        .A(n1350), .ZN(n1347) );
  AOI21_X1 U8839 ( .B1(\mult_22/CARRYB[63][40] ), .B2(\mult_22/SUMB[63][41] ), 
        .A(n1409), .ZN(n1395) );
  AOI21_X1 U8840 ( .B1(\mult_22/CARRYB[63][31] ), .B2(\mult_22/SUMB[63][32] ), 
        .A(n1451), .ZN(n1448) );
  AOI21_X1 U8841 ( .B1(\mult_22/CARRYB[63][46] ), .B2(\mult_22/SUMB[63][47] ), 
        .A(n1368), .ZN(n1361) );
  AOI21_X1 U8842 ( .B1(\mult_22/CARRYB[63][32] ), .B2(\mult_22/SUMB[63][33] ), 
        .A(n1449), .ZN(n1442) );
  AOI21_X1 U8843 ( .B1(\mult_22/CARRYB[63][30] ), .B2(\mult_22/SUMB[63][31] ), 
        .A(n1459), .ZN(n1452) );
  AOI21_X1 U8844 ( .B1(\mult_22/CARRYB[63][48] ), .B2(\mult_22/SUMB[63][49] ), 
        .A(n1358), .ZN(n1351) );
  AOI21_X1 U8845 ( .B1(\mult_22/CARRYB[63][50] ), .B2(\mult_22/SUMB[63][51] ), 
        .A(n1348), .ZN(n1341) );
  AOI21_X1 U8846 ( .B1(\mult_22/CARRYB[63][44] ), .B2(\mult_22/SUMB[63][45] ), 
        .A(n1386), .ZN(n1371) );
  AND3_X1 U8847 ( .A1(\mult_22/CARRYB[63][43] ), .A2(n1388), .A3(
        \mult_22/SUMB[63][44] ), .ZN(n1378) );
  INV_X1 U8848 ( .A(n1435), .ZN(n615) );
  AOI21_X1 U8849 ( .B1(\mult_22/SUMB[63][36] ), .B2(\mult_22/CARRYB[63][35] ), 
        .A(n1434), .ZN(n1435) );
  NAND2_X1 U8850 ( .A1(\mult_22/SUMB[63][57] ), .A2(\mult_22/CARRYB[63][56] ), 
        .ZN(n1313) );
  NAND2_X1 U8851 ( .A1(\mult_22/SUMB[63][29] ), .A2(\mult_22/CARRYB[63][28] ), 
        .ZN(n1463) );
  AND3_X1 U8852 ( .A1(\mult_22/CARRYB[63][39] ), .A2(n1411), .A3(
        \mult_22/SUMB[63][40] ), .ZN(n1399) );
  AND3_X1 U8853 ( .A1(\mult_22/CARRYB[63][31] ), .A2(n1451), .A3(
        \mult_22/SUMB[63][32] ), .ZN(n1447) );
  AND3_X1 U8854 ( .A1(\mult_22/CARRYB[63][29] ), .A2(n1461), .A3(
        \mult_22/SUMB[63][30] ), .ZN(n1457) );
  AND3_X1 U8855 ( .A1(\mult_22/CARRYB[63][45] ), .A2(n1370), .A3(
        \mult_22/SUMB[63][46] ), .ZN(n1366) );
  AND3_X1 U8856 ( .A1(\mult_22/CARRYB[63][47] ), .A2(n1360), .A3(
        \mult_22/SUMB[63][48] ), .ZN(n1356) );
  AND3_X1 U8857 ( .A1(\mult_22/SUMB[63][50] ), .A2(n1350), .A3(
        \mult_22/CARRYB[63][49] ), .ZN(n1346) );
  AND3_X1 U8858 ( .A1(\mult_22/CARRYB[63][51] ), .A2(n1340), .A3(
        \mult_22/SUMB[63][52] ), .ZN(n1336) );
  AND3_X1 U8859 ( .A1(\mult_22/CARRYB[63][55] ), .A2(n1320), .A3(
        \mult_22/SUMB[63][56] ), .ZN(n1317) );
  AND3_X1 U8860 ( .A1(\mult_22/SUMB[63][58] ), .A2(n1310), .A3(
        \mult_22/CARRYB[63][57] ), .ZN(n1305) );
  AND2_X1 U8861 ( .A1(\mult_22/SUMB[63][28] ), .A2(\mult_22/CARRYB[63][27] ), 
        .ZN(n1479) );
  XNOR2_X1 U8862 ( .A(\mult_22/CARRYB[63][61] ), .B(\mult_22/SUMB[63][62] ), 
        .ZN(n1291) );
  AOI21_X1 U8863 ( .B1(\mult_22/CARRYB[63][59] ), .B2(\mult_22/SUMB[63][60] ), 
        .A(n1299), .ZN(n1297) );
  NAND2_X1 U8864 ( .A1(\mult_22/SUMB[63][61] ), .A2(\mult_22/CARRYB[63][60] ), 
        .ZN(n1292) );
  INV_X1 U8865 ( .A(\mult_22/CARRYB[63][62] ), .ZN(n652) );
  AND3_X1 U8866 ( .A1(\mult_22/CARRYB[63][59] ), .A2(n1299), .A3(
        \mult_22/SUMB[63][60] ), .ZN(n1296) );
  AND2_X1 U8867 ( .A1(\mult_22/SUMB[63][59] ), .A2(\mult_22/CARRYB[63][58] ), 
        .ZN(n1308) );
  AOI21_X1 U8868 ( .B1(\mult_20/CARRYB[31][6] ), .B2(\mult_20/SUMB[31][7] ), 
        .A(n1776), .ZN(n1763) );
  AOI21_X1 U8869 ( .B1(\mult_19/CARRYB[31][6] ), .B2(\mult_19/SUMB[31][7] ), 
        .A(n1250), .ZN(n1237) );
  AOI21_X1 U8870 ( .B1(\mult_20/CARRYB[31][7] ), .B2(\mult_20/SUMB[31][8] ), 
        .A(n1772), .ZN(n1762) );
  AOI21_X1 U8871 ( .B1(\mult_19/CARRYB[31][7] ), .B2(\mult_19/SUMB[31][8] ), 
        .A(n1246), .ZN(n1236) );
  AOI21_X1 U8872 ( .B1(\mult_20/SUMB[31][3] ), .B2(\mult_20/CARRYB[31][2] ), 
        .A(n1795), .ZN(n1102) );
  AOI21_X1 U8873 ( .B1(\mult_20/SUMB[31][5] ), .B2(\mult_20/CARRYB[31][4] ), 
        .A(n1791), .ZN(n1780) );
  AOI21_X1 U8874 ( .B1(\mult_19/SUMB[31][5] ), .B2(\mult_19/CARRYB[31][4] ), 
        .A(n1266), .ZN(n1254) );
  AOI21_X1 U8875 ( .B1(\mult_19/SUMB[31][3] ), .B2(\mult_19/CARRYB[31][2] ), 
        .A(n1274), .ZN(n1262) );
  AOI21_X1 U8876 ( .B1(\mult_20/CARRYB[31][10] ), .B2(\mult_20/SUMB[31][11] ), 
        .A(n1751), .ZN(n1736) );
  AOI21_X1 U8877 ( .B1(\mult_19/CARRYB[31][10] ), .B2(\mult_19/SUMB[31][11] ), 
        .A(n1225), .ZN(n1210) );
  XNOR2_X1 U8878 ( .A(\mult_20/CARRYB[31][9] ), .B(\mult_20/SUMB[31][10] ), 
        .ZN(n1756) );
  XNOR2_X1 U8879 ( .A(\mult_19/CARRYB[31][9] ), .B(\mult_19/SUMB[31][10] ), 
        .ZN(n1230) );
  AOI21_X1 U8880 ( .B1(\mult_20/CARRYB[31][11] ), .B2(\mult_20/SUMB[31][12] ), 
        .A(n1747), .ZN(n1744) );
  AOI21_X1 U8881 ( .B1(\mult_19/CARRYB[31][11] ), .B2(\mult_19/SUMB[31][12] ), 
        .A(n1221), .ZN(n1218) );
  AOI21_X1 U8882 ( .B1(\mult_20/SUMB[31][4] ), .B2(\mult_20/CARRYB[31][3] ), 
        .A(n1798), .ZN(n1792) );
  XNOR2_X1 U8883 ( .A(\mult_19/CARRYB[31][2] ), .B(\mult_19/SUMB[31][3] ), 
        .ZN(n1277) );
  XNOR2_X1 U8884 ( .A(\mult_20/CARRYB[31][10] ), .B(\mult_20/SUMB[31][11] ), 
        .ZN(n1754) );
  XNOR2_X1 U8885 ( .A(\mult_19/CARRYB[31][10] ), .B(\mult_19/SUMB[31][11] ), 
        .ZN(n1228) );
  XNOR2_X1 U8886 ( .A(\mult_20/CARRYB[31][6] ), .B(\mult_20/SUMB[31][7] ), 
        .ZN(n1779) );
  XNOR2_X1 U8887 ( .A(\mult_19/CARRYB[31][6] ), .B(\mult_19/SUMB[31][7] ), 
        .ZN(n1253) );
  OAI21_X1 U8888 ( .B1(n1681), .B2(n1674), .A(n1673), .ZN(n1675) );
  AND2_X1 U8889 ( .A1(\mult_20/SUMB[31][24] ), .A2(\mult_20/CARRYB[31][23] ), 
        .ZN(n1681) );
  OAI21_X1 U8890 ( .B1(n1668), .B2(n1662), .A(n1661), .ZN(n1663) );
  AND2_X1 U8891 ( .A1(\mult_20/SUMB[31][26] ), .A2(\mult_20/CARRYB[31][25] ), 
        .ZN(n1668) );
  OAI21_X1 U8892 ( .B1(n1656), .B2(n1650), .A(n1649), .ZN(n1651) );
  AND2_X1 U8893 ( .A1(\mult_20/SUMB[31][28] ), .A2(\mult_20/CARRYB[31][27] ), 
        .ZN(n1656) );
  OAI21_X1 U8894 ( .B1(n1155), .B2(n1148), .A(n1147), .ZN(n1149) );
  AND2_X1 U8895 ( .A1(\mult_19/SUMB[31][24] ), .A2(\mult_19/CARRYB[31][23] ), 
        .ZN(n1155) );
  OAI21_X1 U8896 ( .B1(n1142), .B2(n1136), .A(n1135), .ZN(n1137) );
  AND2_X1 U8897 ( .A1(\mult_19/SUMB[31][26] ), .A2(\mult_19/CARRYB[31][25] ), 
        .ZN(n1142) );
  OAI21_X1 U8898 ( .B1(n1130), .B2(n1124), .A(n1123), .ZN(n1125) );
  AND2_X1 U8899 ( .A1(\mult_19/SUMB[31][28] ), .A2(\mult_19/CARRYB[31][27] ), 
        .ZN(n1130) );
  NAND2_X1 U8900 ( .A1(n1638), .A2(n393), .ZN(n1639) );
  INV_X1 U8901 ( .A(n1644), .ZN(n393) );
  AOI21_X1 U8902 ( .B1(\mult_20/SUMB[31][30] ), .B2(\mult_20/CARRYB[31][29] ), 
        .A(n394), .ZN(n1644) );
  NAND2_X1 U8903 ( .A1(n1112), .A2(n487), .ZN(n1113) );
  INV_X1 U8904 ( .A(n1118), .ZN(n487) );
  AOI21_X1 U8905 ( .B1(\mult_19/SUMB[31][30] ), .B2(\mult_19/CARRYB[31][29] ), 
        .A(n488), .ZN(n1118) );
  INV_X1 U8906 ( .A(n1271), .ZN(n511) );
  AOI21_X1 U8907 ( .B1(\mult_19/SUMB[31][4] ), .B2(\mult_19/CARRYB[31][3] ), 
        .A(n1272), .ZN(n1271) );
  INV_X1 U8908 ( .A(n1658), .ZN(n396) );
  OAI21_X1 U8909 ( .B1(n1659), .B2(n1660), .A(n1661), .ZN(n1658) );
  AOI21_X1 U8910 ( .B1(\mult_20/CARRYB[31][25] ), .B2(\mult_20/SUMB[31][26] ), 
        .A(n1662), .ZN(n1660) );
  INV_X1 U8911 ( .A(n1132), .ZN(n490) );
  OAI21_X1 U8912 ( .B1(n1133), .B2(n1134), .A(n1135), .ZN(n1132) );
  AOI21_X1 U8913 ( .B1(\mult_19/CARRYB[31][25] ), .B2(\mult_19/SUMB[31][26] ), 
        .A(n1136), .ZN(n1134) );
  INV_X1 U8914 ( .A(n1646), .ZN(n395) );
  OAI21_X1 U8915 ( .B1(n1647), .B2(n1648), .A(n1649), .ZN(n1646) );
  AOI21_X1 U8916 ( .B1(\mult_20/CARRYB[31][27] ), .B2(\mult_20/SUMB[31][28] ), 
        .A(n1650), .ZN(n1648) );
  INV_X1 U8917 ( .A(n1120), .ZN(n489) );
  OAI21_X1 U8918 ( .B1(n1121), .B2(n1122), .A(n1123), .ZN(n1120) );
  AOI21_X1 U8919 ( .B1(\mult_19/CARRYB[31][27] ), .B2(\mult_19/SUMB[31][28] ), 
        .A(n1124), .ZN(n1122) );
  NAND2_X1 U8920 ( .A1(\mult_20/SUMB[31][9] ), .A2(\mult_20/CARRYB[31][8] ), 
        .ZN(n1757) );
  NAND2_X1 U8921 ( .A1(\mult_19/SUMB[31][9] ), .A2(\mult_19/CARRYB[31][8] ), 
        .ZN(n1231) );
  AND3_X1 U8922 ( .A1(\mult_20/CARRYB[31][11] ), .A2(n1747), .A3(
        \mult_20/SUMB[31][12] ), .ZN(n1735) );
  AND3_X1 U8923 ( .A1(\mult_19/CARRYB[31][11] ), .A2(n1221), .A3(
        \mult_19/SUMB[31][12] ), .ZN(n1209) );
  AND3_X1 U8924 ( .A1(\mult_20/CARRYB[31][7] ), .A2(n1772), .A3(
        \mult_20/SUMB[31][8] ), .ZN(n1765) );
  AND3_X1 U8925 ( .A1(\mult_19/CARRYB[31][7] ), .A2(n1246), .A3(
        \mult_19/SUMB[31][8] ), .ZN(n1239) );
  NAND2_X1 U8926 ( .A1(\mult_20/SUMB[31][10] ), .A2(\mult_20/CARRYB[31][9] ), 
        .ZN(n1753) );
  NAND2_X1 U8927 ( .A1(\mult_19/SUMB[31][10] ), .A2(\mult_19/CARRYB[31][9] ), 
        .ZN(n1227) );
  NAND2_X1 U8928 ( .A1(\mult_20/SUMB[31][6] ), .A2(\mult_20/CARRYB[31][5] ), 
        .ZN(n1778) );
  NAND2_X1 U8929 ( .A1(\mult_19/SUMB[31][2] ), .A2(\mult_19/CARRYB[31][1] ), 
        .ZN(n1278) );
  NAND2_X1 U8930 ( .A1(\mult_19/SUMB[31][6] ), .A2(\mult_19/CARRYB[31][5] ), 
        .ZN(n1252) );
  AND2_X1 U8931 ( .A1(\mult_20/SUMB[31][2] ), .A2(\mult_20/CARRYB[31][1] ), 
        .ZN(n1796) );
  INV_X1 U8932 ( .A(n1670), .ZN(n397) );
  OAI21_X1 U8933 ( .B1(n1671), .B2(n1672), .A(n1673), .ZN(n1670) );
  AOI21_X1 U8934 ( .B1(\mult_20/CARRYB[31][23] ), .B2(\mult_20/SUMB[31][24] ), 
        .A(n1674), .ZN(n1672) );
  INV_X1 U8935 ( .A(n1144), .ZN(n491) );
  OAI21_X1 U8936 ( .B1(n1145), .B2(n1146), .A(n1147), .ZN(n1144) );
  AOI21_X1 U8937 ( .B1(\mult_19/CARRYB[31][23] ), .B2(\mult_19/SUMB[31][24] ), 
        .A(n1148), .ZN(n1146) );
  XNOR2_X1 U8938 ( .A(\mult_20/CARRYB[31][23] ), .B(\mult_20/SUMB[31][24] ), 
        .ZN(n1680) );
  XNOR2_X1 U8939 ( .A(\mult_19/CARRYB[31][23] ), .B(\mult_19/SUMB[31][24] ), 
        .ZN(n1154) );
  XNOR2_X1 U8940 ( .A(\mult_20/CARRYB[31][21] ), .B(\mult_20/SUMB[31][22] ), 
        .ZN(n1692) );
  XNOR2_X1 U8941 ( .A(\mult_19/CARRYB[31][21] ), .B(\mult_19/SUMB[31][22] ), 
        .ZN(n1166) );
  AOI21_X1 U8942 ( .B1(\mult_20/CARRYB[31][21] ), .B2(\mult_20/SUMB[31][22] ), 
        .A(n1687), .ZN(n1684) );
  AOI21_X1 U8943 ( .B1(\mult_19/CARRYB[31][21] ), .B2(\mult_19/SUMB[31][22] ), 
        .A(n1161), .ZN(n1158) );
  AOI21_X1 U8944 ( .B1(\mult_20/CARRYB[31][19] ), .B2(\mult_20/SUMB[31][20] ), 
        .A(n1698), .ZN(n1694) );
  AOI21_X1 U8945 ( .B1(\mult_19/CARRYB[31][19] ), .B2(\mult_19/SUMB[31][20] ), 
        .A(n1172), .ZN(n1168) );
  AOI21_X1 U8946 ( .B1(\mult_20/SUMB[31][17] ), .B2(\mult_20/CARRYB[31][16] ), 
        .A(n1717), .ZN(n1711) );
  AOI21_X1 U8947 ( .B1(\mult_19/SUMB[31][17] ), .B2(\mult_19/CARRYB[31][16] ), 
        .A(n1191), .ZN(n1185) );
  AOI21_X1 U8948 ( .B1(\mult_20/CARRYB[31][13] ), .B2(\mult_20/SUMB[31][14] ), 
        .A(n1730), .ZN(n1728) );
  AOI21_X1 U8949 ( .B1(\mult_19/CARRYB[31][13] ), .B2(\mult_19/SUMB[31][14] ), 
        .A(n1204), .ZN(n1202) );
  AOI21_X1 U8950 ( .B1(\mult_20/CARRYB[31][15] ), .B2(\mult_20/SUMB[31][16] ), 
        .A(n1719), .ZN(n1716) );
  AOI21_X1 U8951 ( .B1(\mult_19/CARRYB[31][15] ), .B2(\mult_19/SUMB[31][16] ), 
        .A(n1193), .ZN(n1190) );
  AOI21_X1 U8952 ( .B1(\mult_20/CARRYB[31][17] ), .B2(\mult_20/SUMB[31][18] ), 
        .A(n1709), .ZN(n1707) );
  AOI21_X1 U8953 ( .B1(\mult_19/CARRYB[31][17] ), .B2(\mult_19/SUMB[31][18] ), 
        .A(n1183), .ZN(n1181) );
  AOI21_X1 U8954 ( .B1(\mult_20/CARRYB[31][12] ), .B2(\mult_20/SUMB[31][13] ), 
        .A(n1745), .ZN(n1731) );
  AOI21_X1 U8955 ( .B1(\mult_19/CARRYB[31][12] ), .B2(\mult_19/SUMB[31][13] ), 
        .A(n1219), .ZN(n1205) );
  NAND2_X1 U8956 ( .A1(\mult_20/SUMB[31][21] ), .A2(\mult_20/CARRYB[31][20] ), 
        .ZN(n1691) );
  NAND2_X1 U8957 ( .A1(\mult_19/SUMB[31][21] ), .A2(\mult_19/CARRYB[31][20] ), 
        .ZN(n1165) );
  NAND2_X1 U8958 ( .A1(\mult_20/SUMB[31][23] ), .A2(\mult_20/CARRYB[31][22] ), 
        .ZN(n1679) );
  NAND2_X1 U8959 ( .A1(\mult_19/SUMB[31][23] ), .A2(\mult_19/CARRYB[31][22] ), 
        .ZN(n1153) );
  AND2_X1 U8960 ( .A1(\mult_20/SUMB[31][19] ), .A2(\mult_20/CARRYB[31][18] ), 
        .ZN(n1702) );
  AND2_X1 U8961 ( .A1(\mult_19/SUMB[31][19] ), .A2(\mult_19/CARRYB[31][18] ), 
        .ZN(n1176) );
  AND3_X1 U8962 ( .A1(\mult_20/CARRYB[31][15] ), .A2(n1719), .A3(
        \mult_20/SUMB[31][16] ), .ZN(n1715) );
  AND3_X1 U8963 ( .A1(\mult_19/CARRYB[31][15] ), .A2(n1193), .A3(
        \mult_19/SUMB[31][16] ), .ZN(n1189) );
  AND3_X1 U8964 ( .A1(\mult_20/CARRYB[31][13] ), .A2(n1730), .A3(
        \mult_20/SUMB[31][14] ), .ZN(n1727) );
  AND3_X1 U8965 ( .A1(\mult_19/CARRYB[31][13] ), .A2(n1204), .A3(
        \mult_19/SUMB[31][14] ), .ZN(n1201) );
  AND3_X1 U8966 ( .A1(\mult_20/SUMB[31][18] ), .A2(n1709), .A3(
        \mult_20/CARRYB[31][17] ), .ZN(n1706) );
  AND3_X1 U8967 ( .A1(\mult_19/SUMB[31][18] ), .A2(n1183), .A3(
        \mult_19/CARRYB[31][17] ), .ZN(n1180) );
  AND2_X1 U8968 ( .A1(\mult_20/CARRYB[31][14] ), .A2(\mult_20/SUMB[31][15] ), 
        .ZN(n1724) );
  AND2_X1 U8969 ( .A1(\mult_19/CARRYB[31][14] ), .A2(\mult_19/SUMB[31][15] ), 
        .ZN(n1198) );
  XNOR2_X1 U8970 ( .A(\mult_20/CARRYB[31][25] ), .B(\mult_20/SUMB[31][26] ), 
        .ZN(n1667) );
  XNOR2_X1 U8971 ( .A(\mult_19/CARRYB[31][25] ), .B(\mult_19/SUMB[31][26] ), 
        .ZN(n1141) );
  XNOR2_X1 U8972 ( .A(\mult_20/CARRYB[31][27] ), .B(\mult_20/SUMB[31][28] ), 
        .ZN(n1655) );
  XNOR2_X1 U8973 ( .A(\mult_19/CARRYB[31][27] ), .B(\mult_19/SUMB[31][28] ), 
        .ZN(n1129) );
  XNOR2_X1 U8974 ( .A(\mult_20/CARRYB[31][29] ), .B(\mult_20/SUMB[31][30] ), 
        .ZN(n1643) );
  XNOR2_X1 U8975 ( .A(\mult_19/CARRYB[31][29] ), .B(\mult_19/SUMB[31][30] ), 
        .ZN(n1117) );
  NAND2_X1 U8976 ( .A1(\mult_20/SUMB[31][25] ), .A2(\mult_20/CARRYB[31][24] ), 
        .ZN(n1666) );
  NAND2_X1 U8977 ( .A1(\mult_19/SUMB[31][25] ), .A2(\mult_19/CARRYB[31][24] ), 
        .ZN(n1140) );
  NAND2_X1 U8978 ( .A1(\mult_20/SUMB[31][27] ), .A2(\mult_20/CARRYB[31][26] ), 
        .ZN(n1654) );
  NAND2_X1 U8979 ( .A1(\mult_19/SUMB[31][27] ), .A2(\mult_19/CARRYB[31][26] ), 
        .ZN(n1128) );
  NAND2_X1 U8980 ( .A1(\mult_20/SUMB[31][29] ), .A2(\mult_20/CARRYB[31][28] ), 
        .ZN(n1642) );
  NAND2_X1 U8981 ( .A1(\mult_19/SUMB[31][29] ), .A2(\mult_19/CARRYB[31][28] ), 
        .ZN(n1116) );
  NOR2_X1 U8982 ( .A1(n514), .A2(n1279), .ZN(N33) );
  AOI21_X1 U8983 ( .B1(\mult_19/SUMB[31][1] ), .B2(\mult_19/CARRYB[31][0] ), 
        .A(n1280), .ZN(n1279) );
  NOR2_X1 U8984 ( .A1(n421), .A2(n1106), .ZN(N97) );
  AOI21_X1 U8985 ( .B1(\mult_20/SUMB[31][1] ), .B2(\mult_20/CARRYB[31][0] ), 
        .A(n1107), .ZN(n1106) );
  INV_X1 U8986 ( .A(n1103), .ZN(n421) );
  INV_X1 U8987 ( .A(n3498), .ZN(n3493) );
  INV_X1 U8988 ( .A(n3511), .ZN(n3502) );
  NOR2_X1 U8989 ( .A1(n2422), .A2(n3119), .ZN(\mult_22/ab[63][7] ) );
  NOR2_X1 U8990 ( .A1(n2684), .A2(n2781), .ZN(\mult_22/ab[7][51] ) );
  NOR2_X1 U8991 ( .A1(n2581), .A2(n2876), .ZN(\mult_22/ab[23][33] ) );
  NOR2_X1 U8992 ( .A1(n2569), .A2(n2900), .ZN(\mult_22/ab[27][31] ) );
  NOR2_X1 U8993 ( .A1(n2398), .A2(n3116), .ZN(\mult_22/ab[63][3] ) );
  NOR2_X1 U8994 ( .A1(n2428), .A2(n3119), .ZN(\mult_22/ab[63][8] ) );
  NOR2_X1 U8995 ( .A1(n2434), .A2(n3119), .ZN(\mult_22/ab[63][9] ) );
  NOR2_X1 U8996 ( .A1(n2444), .A2(n3114), .ZN(\mult_22/ab[63][10] ) );
  NOR2_X1 U8997 ( .A1(n2416), .A2(n3118), .ZN(\mult_22/ab[63][6] ) );
  NOR2_X1 U8998 ( .A1(n2665), .A2(n2799), .ZN(\mult_22/ab[10][47] ) );
  NOR2_X1 U8999 ( .A1(n2392), .A2(n3115), .ZN(\mult_22/ab[63][2] ) );
  NOR2_X1 U9000 ( .A1(n2408), .A2(n3117), .ZN(\mult_22/ab[63][4] ) );
  NOR2_X1 U9001 ( .A1(n2624), .A2(n2840), .ZN(\mult_22/ab[17][41] ) );
  NOR2_X1 U9002 ( .A1(n2573), .A2(n2876), .ZN(\mult_22/ab[23][32] ) );
  NOR2_X1 U9003 ( .A1(n2563), .A2(n2899), .ZN(\mult_22/ab[27][30] ) );
  NOR2_X1 U9004 ( .A1(n2410), .A2(n3118), .ZN(\mult_22/ab[63][5] ) );
  NOR2_X1 U9005 ( .A1(n2386), .A2(n3114), .ZN(\mult_22/ab[63][1] ) );
  NOR2_X1 U9006 ( .A1(n2616), .A2(n2864), .ZN(\mult_22/ab[21][39] ) );
  NOR2_X1 U9007 ( .A1(n2551), .A2(n2929), .ZN(\mult_22/ab[32][28] ) );
  NOR2_X1 U9008 ( .A1(n2678), .A2(n2781), .ZN(\mult_22/ab[7][50] ) );
  NOR2_X1 U9009 ( .A1(n2384), .A2(n3114), .ZN(\mult_22/ab[63][0] ) );
  INV_X1 U9010 ( .A(n1285), .ZN(n651) );
  NOR2_X1 U9011 ( .A1(n2743), .A2(n2758), .ZN(\mult_22/ab[3][62] ) );
  NOR2_X1 U9012 ( .A1(n2408), .A2(n3105), .ZN(\mult_22/ab[61][4] ) );
  NOR2_X1 U9013 ( .A1(n2398), .A2(n3110), .ZN(\mult_22/ab[62][3] ) );
  NOR2_X1 U9014 ( .A1(n2416), .A2(n3095), .ZN(\mult_22/ab[59][6] ) );
  NOR2_X1 U9015 ( .A1(n2429), .A2(n3083), .ZN(\mult_22/ab[57][8] ) );
  NOR2_X1 U9016 ( .A1(n2444), .A2(n3066), .ZN(\mult_22/ab[55][10] ) );
  NOR2_X1 U9017 ( .A1(n2453), .A2(n3054), .ZN(\mult_22/ab[53][12] ) );
  NOR2_X1 U9018 ( .A1(n2465), .A2(n3030), .ZN(\mult_22/ab[49][14] ) );
  NOR2_X1 U9019 ( .A1(n2622), .A2(n2840), .ZN(\mult_22/ab[17][40] ) );
  NOR2_X1 U9020 ( .A1(n2186), .A2(n2776), .ZN(\mult_22/ab[6][62] ) );
  NOR2_X1 U9021 ( .A1(n2748), .A2(n2770), .ZN(\mult_22/ab[5][63] ) );
  NOR2_X1 U9022 ( .A1(n2185), .A2(n2782), .ZN(\mult_22/ab[7][62] ) );
  NOR2_X1 U9023 ( .A1(n2748), .A2(n2776), .ZN(\mult_22/ab[6][63] ) );
  NOR2_X1 U9024 ( .A1(n2748), .A2(n2782), .ZN(\mult_22/ab[7][63] ) );
  NOR2_X1 U9025 ( .A1(n2185), .A2(n2788), .ZN(\mult_22/ab[8][62] ) );
  NOR2_X1 U9026 ( .A1(n2185), .A2(n2794), .ZN(\mult_22/ab[9][62] ) );
  NOR2_X1 U9027 ( .A1(n2748), .A2(n2788), .ZN(\mult_22/ab[8][63] ) );
  NOR2_X1 U9028 ( .A1(n2745), .A2(n2800), .ZN(\mult_22/ab[10][62] ) );
  NOR2_X1 U9029 ( .A1(n2750), .A2(n2794), .ZN(\mult_22/ab[9][63] ) );
  NOR2_X1 U9030 ( .A1(n2750), .A2(n2758), .ZN(\mult_22/ab[3][63] ) );
  NOR2_X1 U9031 ( .A1(n2186), .A2(n2764), .ZN(\mult_22/ab[4][62] ) );
  NOR2_X1 U9032 ( .A1(n2186), .A2(n2770), .ZN(\mult_22/ab[5][62] ) );
  NOR2_X1 U9033 ( .A1(n2749), .A2(n2764), .ZN(\mult_22/ab[4][63] ) );
  NOR2_X1 U9034 ( .A1(n2739), .A2(n2764), .ZN(\mult_22/ab[4][61] ) );
  NOR2_X1 U9035 ( .A1(n2410), .A2(n3112), .ZN(\mult_22/ab[62][5] ) );
  NOR2_X1 U9036 ( .A1(n2416), .A2(n3113), .ZN(\mult_22/ab[62][6] ) );
  NOR2_X1 U9037 ( .A1(n2428), .A2(n3113), .ZN(\mult_22/ab[62][8] ) );
  NOR2_X1 U9038 ( .A1(n2408), .A2(n3111), .ZN(\mult_22/ab[62][4] ) );
  NOR2_X1 U9039 ( .A1(n2434), .A2(n3113), .ZN(\mult_22/ab[62][9] ) );
  NOR2_X1 U9040 ( .A1(n2422), .A2(n3113), .ZN(\mult_22/ab[62][7] ) );
  NOR2_X1 U9041 ( .A1(n2410), .A2(n3106), .ZN(\mult_22/ab[61][5] ) );
  NOR2_X1 U9042 ( .A1(n2416), .A2(n3107), .ZN(\mult_22/ab[61][6] ) );
  NOR2_X1 U9043 ( .A1(n2422), .A2(n3107), .ZN(\mult_22/ab[61][7] ) );
  NOR2_X1 U9044 ( .A1(n2428), .A2(n3107), .ZN(\mult_22/ab[61][8] ) );
  NOR2_X1 U9045 ( .A1(n2434), .A2(n3107), .ZN(\mult_22/ab[61][9] ) );
  NOR2_X1 U9046 ( .A1(n2444), .A2(n3108), .ZN(\mult_22/ab[62][10] ) );
  NOR2_X1 U9047 ( .A1(n2416), .A2(n3101), .ZN(\mult_22/ab[60][6] ) );
  NOR2_X1 U9048 ( .A1(n2444), .A2(n3102), .ZN(\mult_22/ab[61][10] ) );
  NOR2_X1 U9049 ( .A1(n2422), .A2(n3101), .ZN(\mult_22/ab[60][7] ) );
  NOR2_X1 U9050 ( .A1(n2410), .A2(n3100), .ZN(\mult_22/ab[60][5] ) );
  NOR2_X1 U9051 ( .A1(n2446), .A2(n3108), .ZN(\mult_22/ab[62][11] ) );
  NOR2_X1 U9052 ( .A1(n2428), .A2(n3101), .ZN(\mult_22/ab[60][8] ) );
  NOR2_X1 U9053 ( .A1(n2434), .A2(n3101), .ZN(\mult_22/ab[60][9] ) );
  NOR2_X1 U9054 ( .A1(n2444), .A2(n3096), .ZN(\mult_22/ab[60][10] ) );
  NOR2_X1 U9055 ( .A1(n2446), .A2(n3102), .ZN(\mult_22/ab[61][11] ) );
  NOR2_X1 U9056 ( .A1(n2422), .A2(n3095), .ZN(\mult_22/ab[59][7] ) );
  NOR2_X1 U9057 ( .A1(n2452), .A2(n3102), .ZN(\mult_22/ab[61][12] ) );
  NOR2_X1 U9058 ( .A1(n2428), .A2(n3095), .ZN(\mult_22/ab[59][8] ) );
  NOR2_X1 U9059 ( .A1(n2446), .A2(n3096), .ZN(\mult_22/ab[60][11] ) );
  NOR2_X1 U9060 ( .A1(n2434), .A2(n3095), .ZN(\mult_22/ab[59][9] ) );
  NOR2_X1 U9061 ( .A1(n2444), .A2(n3090), .ZN(\mult_22/ab[59][10] ) );
  NOR2_X1 U9062 ( .A1(n2410), .A2(n3094), .ZN(\mult_22/ab[59][5] ) );
  NOR2_X1 U9063 ( .A1(n2446), .A2(n3090), .ZN(\mult_22/ab[59][11] ) );
  NOR2_X1 U9064 ( .A1(n2422), .A2(n3089), .ZN(\mult_22/ab[58][7] ) );
  NOR2_X1 U9065 ( .A1(n2428), .A2(n3089), .ZN(\mult_22/ab[58][8] ) );
  NOR2_X1 U9066 ( .A1(n2452), .A2(n3096), .ZN(\mult_22/ab[60][12] ) );
  NOR2_X1 U9067 ( .A1(n2458), .A2(n3096), .ZN(\mult_22/ab[60][13] ) );
  NOR2_X1 U9068 ( .A1(n2434), .A2(n3089), .ZN(\mult_22/ab[58][9] ) );
  NOR2_X1 U9069 ( .A1(n2444), .A2(n3084), .ZN(\mult_22/ab[58][10] ) );
  NOR2_X1 U9070 ( .A1(n2446), .A2(n3084), .ZN(\mult_22/ab[58][11] ) );
  NOR2_X1 U9071 ( .A1(n2452), .A2(n3090), .ZN(\mult_22/ab[59][12] ) );
  NOR2_X1 U9072 ( .A1(n2423), .A2(n3083), .ZN(\mult_22/ab[57][7] ) );
  NOR2_X1 U9073 ( .A1(n2411), .A2(n3088), .ZN(\mult_22/ab[58][5] ) );
  NOR2_X1 U9074 ( .A1(n2435), .A2(n3083), .ZN(\mult_22/ab[57][9] ) );
  NOR2_X1 U9075 ( .A1(n2444), .A2(n3078), .ZN(\mult_22/ab[57][10] ) );
  NOR2_X1 U9076 ( .A1(n2458), .A2(n3090), .ZN(\mult_22/ab[59][13] ) );
  NOR2_X1 U9077 ( .A1(n2447), .A2(n3078), .ZN(\mult_22/ab[57][11] ) );
  NOR2_X1 U9078 ( .A1(n2452), .A2(n3084), .ZN(\mult_22/ab[58][12] ) );
  NOR2_X1 U9079 ( .A1(n2464), .A2(n3090), .ZN(\mult_22/ab[59][14] ) );
  NOR2_X1 U9080 ( .A1(n2622), .A2(n2858), .ZN(\mult_22/ab[20][40] ) );
  NOR2_X1 U9081 ( .A1(n2435), .A2(n3077), .ZN(\mult_22/ab[56][9] ) );
  NOR2_X1 U9082 ( .A1(n2453), .A2(n3078), .ZN(\mult_22/ab[57][12] ) );
  NOR2_X1 U9083 ( .A1(n2444), .A2(n3072), .ZN(\mult_22/ab[56][10] ) );
  NOR2_X1 U9084 ( .A1(n2447), .A2(n3072), .ZN(\mult_22/ab[56][11] ) );
  NOR2_X1 U9085 ( .A1(n2459), .A2(n3084), .ZN(\mult_22/ab[58][13] ) );
  NOR2_X1 U9086 ( .A1(n2423), .A2(n3077), .ZN(\mult_22/ab[56][7] ) );
  NOR2_X1 U9087 ( .A1(n2464), .A2(n3084), .ZN(\mult_22/ab[58][14] ) );
  NOR2_X1 U9088 ( .A1(n2453), .A2(n3072), .ZN(\mult_22/ab[56][12] ) );
  NOR2_X1 U9089 ( .A1(n2411), .A2(n3082), .ZN(\mult_22/ab[57][5] ) );
  NOR2_X1 U9090 ( .A1(n2435), .A2(n3071), .ZN(\mult_22/ab[55][9] ) );
  NOR2_X1 U9091 ( .A1(n2459), .A2(n3078), .ZN(\mult_22/ab[57][13] ) );
  NOR2_X1 U9092 ( .A1(n2447), .A2(n3066), .ZN(\mult_22/ab[55][11] ) );
  NOR2_X1 U9093 ( .A1(n2470), .A2(n3084), .ZN(\mult_22/ab[58][15] ) );
  NOR2_X1 U9094 ( .A1(n2453), .A2(n3066), .ZN(\mult_22/ab[55][12] ) );
  NOR2_X1 U9095 ( .A1(n2459), .A2(n3072), .ZN(\mult_22/ab[56][13] ) );
  NOR2_X1 U9096 ( .A1(n2423), .A2(n3071), .ZN(\mult_22/ab[55][7] ) );
  NOR2_X1 U9097 ( .A1(n2465), .A2(n3078), .ZN(\mult_22/ab[57][14] ) );
  NOR2_X1 U9098 ( .A1(n2435), .A2(n3065), .ZN(\mult_22/ab[54][9] ) );
  NOR2_X1 U9099 ( .A1(n2447), .A2(n3060), .ZN(\mult_22/ab[54][11] ) );
  NOR2_X1 U9100 ( .A1(n2459), .A2(n3066), .ZN(\mult_22/ab[55][13] ) );
  NOR2_X1 U9101 ( .A1(n2453), .A2(n3060), .ZN(\mult_22/ab[54][12] ) );
  NOR2_X1 U9102 ( .A1(n2471), .A2(n3078), .ZN(\mult_22/ab[57][15] ) );
  NOR2_X1 U9103 ( .A1(n2465), .A2(n3072), .ZN(\mult_22/ab[56][14] ) );
  NOR2_X1 U9104 ( .A1(n2411), .A2(n3076), .ZN(\mult_22/ab[56][5] ) );
  NOR2_X1 U9105 ( .A1(n2459), .A2(n3060), .ZN(\mult_22/ab[54][13] ) );
  NOR2_X1 U9106 ( .A1(n2447), .A2(n3054), .ZN(\mult_22/ab[53][11] ) );
  NOR2_X1 U9107 ( .A1(n2423), .A2(n3065), .ZN(\mult_22/ab[54][7] ) );
  NOR2_X1 U9108 ( .A1(n2465), .A2(n3066), .ZN(\mult_22/ab[55][14] ) );
  NOR2_X1 U9109 ( .A1(n2435), .A2(n3059), .ZN(\mult_22/ab[53][9] ) );
  NOR2_X1 U9110 ( .A1(n2471), .A2(n3072), .ZN(\mult_22/ab[56][15] ) );
  NOR2_X1 U9111 ( .A1(n2477), .A2(n3078), .ZN(\mult_22/ab[57][16] ) );
  NOR2_X1 U9112 ( .A1(n2459), .A2(n3054), .ZN(\mult_22/ab[53][13] ) );
  NOR2_X1 U9113 ( .A1(n2624), .A2(n2846), .ZN(\mult_22/ab[18][41] ) );
  NOR2_X1 U9114 ( .A1(n2465), .A2(n3060), .ZN(\mult_22/ab[54][14] ) );
  NOR2_X1 U9115 ( .A1(n2624), .A2(n2852), .ZN(\mult_22/ab[19][41] ) );
  NOR2_X1 U9116 ( .A1(n2471), .A2(n3066), .ZN(\mult_22/ab[55][15] ) );
  NOR2_X1 U9117 ( .A1(n2477), .A2(n3072), .ZN(\mult_22/ab[56][16] ) );
  NOR2_X1 U9118 ( .A1(n2447), .A2(n3048), .ZN(\mult_22/ab[52][11] ) );
  NOR2_X1 U9119 ( .A1(n2453), .A2(n3048), .ZN(\mult_22/ab[52][12] ) );
  NOR2_X1 U9120 ( .A1(n2465), .A2(n3054), .ZN(\mult_22/ab[53][14] ) );
  NOR2_X1 U9121 ( .A1(n2435), .A2(n3053), .ZN(\mult_22/ab[52][9] ) );
  NOR2_X1 U9122 ( .A1(n2459), .A2(n3048), .ZN(\mult_22/ab[52][13] ) );
  NOR2_X1 U9123 ( .A1(n2471), .A2(n3060), .ZN(\mult_22/ab[54][15] ) );
  NOR2_X1 U9124 ( .A1(n2477), .A2(n3066), .ZN(\mult_22/ab[55][16] ) );
  NOR2_X1 U9125 ( .A1(n2634), .A2(n2835), .ZN(\mult_22/ab[16][42] ) );
  NOR2_X1 U9126 ( .A1(n2411), .A2(n3070), .ZN(\mult_22/ab[55][5] ) );
  NOR2_X1 U9127 ( .A1(n2423), .A2(n3059), .ZN(\mult_22/ab[53][7] ) );
  NOR2_X1 U9128 ( .A1(n2634), .A2(n2829), .ZN(\mult_22/ab[15][42] ) );
  NOR2_X1 U9129 ( .A1(n2465), .A2(n3048), .ZN(\mult_22/ab[52][14] ) );
  NOR2_X1 U9130 ( .A1(n2447), .A2(n3042), .ZN(\mult_22/ab[51][11] ) );
  NOR2_X1 U9131 ( .A1(n2483), .A2(n3072), .ZN(\mult_22/ab[56][17] ) );
  NOR2_X1 U9132 ( .A1(n2471), .A2(n3054), .ZN(\mult_22/ab[53][15] ) );
  NOR2_X1 U9133 ( .A1(n2459), .A2(n3042), .ZN(\mult_22/ab[51][13] ) );
  NOR2_X1 U9134 ( .A1(n2477), .A2(n3060), .ZN(\mult_22/ab[54][16] ) );
  NOR2_X1 U9135 ( .A1(n2483), .A2(n3066), .ZN(\mult_22/ab[55][17] ) );
  NOR2_X1 U9136 ( .A1(n2435), .A2(n3047), .ZN(\mult_22/ab[51][9] ) );
  NOR2_X1 U9137 ( .A1(n2471), .A2(n3048), .ZN(\mult_22/ab[52][15] ) );
  NOR2_X1 U9138 ( .A1(n2447), .A2(n3036), .ZN(\mult_22/ab[50][11] ) );
  NOR2_X1 U9139 ( .A1(n2477), .A2(n3054), .ZN(\mult_22/ab[53][16] ) );
  NOR2_X1 U9140 ( .A1(n2459), .A2(n3036), .ZN(\mult_22/ab[50][13] ) );
  NOR2_X1 U9141 ( .A1(n2483), .A2(n3060), .ZN(\mult_22/ab[54][17] ) );
  NOR2_X1 U9142 ( .A1(n2616), .A2(n2840), .ZN(\mult_22/ab[17][39] ) );
  NOR2_X1 U9143 ( .A1(n2471), .A2(n3042), .ZN(\mult_22/ab[51][15] ) );
  NOR2_X1 U9144 ( .A1(n2634), .A2(n2841), .ZN(\mult_22/ab[17][42] ) );
  NOR2_X1 U9145 ( .A1(n2423), .A2(n3053), .ZN(\mult_22/ab[52][7] ) );
  NOR2_X1 U9146 ( .A1(n2477), .A2(n3048), .ZN(\mult_22/ab[52][16] ) );
  NOR2_X1 U9147 ( .A1(n2411), .A2(n3064), .ZN(\mult_22/ab[54][5] ) );
  NOR2_X1 U9148 ( .A1(n2483), .A2(n3054), .ZN(\mult_22/ab[53][17] ) );
  NOR2_X1 U9149 ( .A1(n2489), .A2(n3066), .ZN(\mult_22/ab[55][18] ) );
  NOR2_X1 U9150 ( .A1(n2471), .A2(n3036), .ZN(\mult_22/ab[50][15] ) );
  NOR2_X1 U9151 ( .A1(n2459), .A2(n3030), .ZN(\mult_22/ab[49][13] ) );
  NOR2_X1 U9152 ( .A1(n2435), .A2(n3041), .ZN(\mult_22/ab[50][9] ) );
  NOR2_X1 U9153 ( .A1(n2447), .A2(n3030), .ZN(\mult_22/ab[49][11] ) );
  NOR2_X1 U9154 ( .A1(n2477), .A2(n3042), .ZN(\mult_22/ab[51][16] ) );
  NOR2_X1 U9155 ( .A1(n2489), .A2(n3060), .ZN(\mult_22/ab[54][18] ) );
  NOR2_X1 U9156 ( .A1(n2636), .A2(n2823), .ZN(\mult_22/ab[14][43] ) );
  NOR2_X1 U9157 ( .A1(n2483), .A2(n3048), .ZN(\mult_22/ab[52][17] ) );
  NOR2_X1 U9158 ( .A1(n2636), .A2(n2829), .ZN(\mult_22/ab[15][43] ) );
  NOR2_X1 U9159 ( .A1(n2471), .A2(n3030), .ZN(\mult_22/ab[49][15] ) );
  NOR2_X1 U9160 ( .A1(n2477), .A2(n3036), .ZN(\mult_22/ab[50][16] ) );
  NOR2_X1 U9161 ( .A1(n2634), .A2(n2846), .ZN(\mult_22/ab[18][42] ) );
  NOR2_X1 U9162 ( .A1(n2489), .A2(n3054), .ZN(\mult_22/ab[53][18] ) );
  NOR2_X1 U9163 ( .A1(n2459), .A2(n3024), .ZN(\mult_22/ab[48][13] ) );
  NOR2_X1 U9164 ( .A1(n2483), .A2(n3042), .ZN(\mult_22/ab[51][17] ) );
  NOR2_X1 U9165 ( .A1(n2636), .A2(n2817), .ZN(\mult_22/ab[13][43] ) );
  NOR2_X1 U9166 ( .A1(n2423), .A2(n3047), .ZN(\mult_22/ab[51][7] ) );
  NOR2_X1 U9167 ( .A1(n2477), .A2(n3030), .ZN(\mult_22/ab[49][16] ) );
  NOR2_X1 U9168 ( .A1(n2447), .A2(n3024), .ZN(\mult_22/ab[48][11] ) );
  NOR2_X1 U9169 ( .A1(n2489), .A2(n3048), .ZN(\mult_22/ab[52][18] ) );
  NOR2_X1 U9170 ( .A1(n2471), .A2(n3024), .ZN(\mult_22/ab[48][15] ) );
  NOR2_X1 U9171 ( .A1(n2611), .A2(n2846), .ZN(\mult_22/ab[18][38] ) );
  NOR2_X1 U9172 ( .A1(n2483), .A2(n3036), .ZN(\mult_22/ab[50][17] ) );
  NOR2_X1 U9173 ( .A1(n2435), .A2(n3035), .ZN(\mult_22/ab[49][9] ) );
  NOR2_X1 U9174 ( .A1(n2495), .A2(n3060), .ZN(\mult_22/ab[54][19] ) );
  NOR2_X1 U9175 ( .A1(n2411), .A2(n3058), .ZN(\mult_22/ab[53][5] ) );
  NOR2_X1 U9176 ( .A1(n2460), .A2(n3018), .ZN(\mult_22/ab[47][13] ) );
  NOR2_X1 U9177 ( .A1(n2489), .A2(n3042), .ZN(\mult_22/ab[51][18] ) );
  NOR2_X1 U9178 ( .A1(n2495), .A2(n3054), .ZN(\mult_22/ab[53][19] ) );
  NOR2_X1 U9179 ( .A1(n2483), .A2(n3030), .ZN(\mult_22/ab[49][17] ) );
  NOR2_X1 U9180 ( .A1(n2636), .A2(n2835), .ZN(\mult_22/ab[16][43] ) );
  NOR2_X1 U9181 ( .A1(n2471), .A2(n3018), .ZN(\mult_22/ab[47][15] ) );
  NOR2_X1 U9182 ( .A1(n2616), .A2(n2834), .ZN(\mult_22/ab[16][39] ) );
  NOR2_X1 U9183 ( .A1(n2495), .A2(n3048), .ZN(\mult_22/ab[52][19] ) );
  NOR2_X1 U9184 ( .A1(n2489), .A2(n3036), .ZN(\mult_22/ab[50][18] ) );
  NOR2_X1 U9185 ( .A1(n2447), .A2(n3018), .ZN(\mult_22/ab[47][11] ) );
  NOR2_X1 U9186 ( .A1(n2483), .A2(n3024), .ZN(\mult_22/ab[48][17] ) );
  NOR2_X1 U9187 ( .A1(n2636), .A2(n2811), .ZN(\mult_22/ab[12][43] ) );
  NOR2_X1 U9188 ( .A1(n2495), .A2(n3042), .ZN(\mult_22/ab[51][19] ) );
  NOR2_X1 U9189 ( .A1(n2489), .A2(n3030), .ZN(\mult_22/ab[49][18] ) );
  NOR2_X1 U9190 ( .A1(n2472), .A2(n3012), .ZN(\mult_22/ab[46][15] ) );
  NOR2_X1 U9191 ( .A1(n2460), .A2(n3012), .ZN(\mult_22/ab[46][13] ) );
  NOR2_X1 U9192 ( .A1(n2423), .A2(n3041), .ZN(\mult_22/ab[50][7] ) );
  NOR2_X1 U9193 ( .A1(n2435), .A2(n3029), .ZN(\mult_22/ab[48][9] ) );
  NOR2_X1 U9194 ( .A1(n2483), .A2(n3018), .ZN(\mult_22/ab[47][17] ) );
  NOR2_X1 U9195 ( .A1(n2495), .A2(n3036), .ZN(\mult_22/ab[50][19] ) );
  NOR2_X1 U9196 ( .A1(n2501), .A2(n3055), .ZN(\mult_22/ab[53][20] ) );
  NOR2_X1 U9197 ( .A1(n2489), .A2(n3024), .ZN(\mult_22/ab[48][18] ) );
  NOR2_X1 U9198 ( .A1(n2646), .A2(n2823), .ZN(\mult_22/ab[14][44] ) );
  NOR2_X1 U9199 ( .A1(n2501), .A2(n3049), .ZN(\mult_22/ab[52][20] ) );
  NOR2_X1 U9200 ( .A1(n2484), .A2(n3012), .ZN(\mult_22/ab[46][17] ) );
  NOR2_X1 U9201 ( .A1(n2495), .A2(n3030), .ZN(\mult_22/ab[49][19] ) );
  NOR2_X1 U9202 ( .A1(n2411), .A2(n3052), .ZN(\mult_22/ab[52][5] ) );
  NOR2_X1 U9203 ( .A1(n2448), .A2(n3012), .ZN(\mult_22/ab[46][11] ) );
  NOR2_X1 U9204 ( .A1(n2472), .A2(n3006), .ZN(\mult_22/ab[45][15] ) );
  NOR2_X1 U9205 ( .A1(n2489), .A2(n3018), .ZN(\mult_22/ab[47][18] ) );
  NOR2_X1 U9206 ( .A1(n2636), .A2(n2841), .ZN(\mult_22/ab[17][43] ) );
  NOR2_X1 U9207 ( .A1(n2501), .A2(n3043), .ZN(\mult_22/ab[51][20] ) );
  NOR2_X1 U9208 ( .A1(n2460), .A2(n3006), .ZN(\mult_22/ab[45][13] ) );
  NOR2_X1 U9209 ( .A1(n2495), .A2(n3024), .ZN(\mult_22/ab[48][19] ) );
  NOR2_X1 U9210 ( .A1(n2501), .A2(n3037), .ZN(\mult_22/ab[50][20] ) );
  NOR2_X1 U9211 ( .A1(n2484), .A2(n3006), .ZN(\mult_22/ab[45][17] ) );
  NOR2_X1 U9212 ( .A1(n2636), .A2(n2805), .ZN(\mult_22/ab[11][43] ) );
  NOR2_X1 U9213 ( .A1(n2435), .A2(n3023), .ZN(\mult_22/ab[47][9] ) );
  NOR2_X1 U9214 ( .A1(n2495), .A2(n3018), .ZN(\mult_22/ab[47][19] ) );
  NOR2_X1 U9215 ( .A1(n2423), .A2(n3035), .ZN(\mult_22/ab[49][7] ) );
  NOR2_X1 U9216 ( .A1(n2611), .A2(n2840), .ZN(\mult_22/ab[17][38] ) );
  NOR2_X1 U9217 ( .A1(n2501), .A2(n3031), .ZN(\mult_22/ab[49][20] ) );
  NOR2_X1 U9218 ( .A1(n2472), .A2(n3000), .ZN(\mult_22/ab[44][15] ) );
  NOR2_X1 U9219 ( .A1(n2646), .A2(n2829), .ZN(\mult_22/ab[15][44] ) );
  NOR2_X1 U9220 ( .A1(n2507), .A2(n3049), .ZN(\mult_22/ab[52][21] ) );
  NOR2_X1 U9221 ( .A1(n2616), .A2(n2828), .ZN(\mult_22/ab[15][39] ) );
  NOR2_X1 U9222 ( .A1(n2484), .A2(n3000), .ZN(\mult_22/ab[44][17] ) );
  NOR2_X1 U9223 ( .A1(n2496), .A2(n3012), .ZN(\mult_22/ab[46][19] ) );
  NOR2_X1 U9224 ( .A1(n2448), .A2(n3006), .ZN(\mult_22/ab[45][11] ) );
  NOR2_X1 U9225 ( .A1(n2501), .A2(n3025), .ZN(\mult_22/ab[48][20] ) );
  NOR2_X1 U9226 ( .A1(n2460), .A2(n3000), .ZN(\mult_22/ab[44][13] ) );
  NOR2_X1 U9227 ( .A1(n2507), .A2(n3043), .ZN(\mult_22/ab[51][21] ) );
  NOR2_X1 U9228 ( .A1(n2507), .A2(n3037), .ZN(\mult_22/ab[50][21] ) );
  NOR2_X1 U9229 ( .A1(n2501), .A2(n3019), .ZN(\mult_22/ab[47][20] ) );
  NOR2_X1 U9230 ( .A1(n2496), .A2(n3006), .ZN(\mult_22/ab[45][19] ) );
  NOR2_X1 U9231 ( .A1(n2411), .A2(n3046), .ZN(\mult_22/ab[51][5] ) );
  NOR2_X1 U9232 ( .A1(n2472), .A2(n2994), .ZN(\mult_22/ab[43][15] ) );
  NOR2_X1 U9233 ( .A1(n2507), .A2(n3031), .ZN(\mult_22/ab[49][21] ) );
  NOR2_X1 U9234 ( .A1(n2484), .A2(n2994), .ZN(\mult_22/ab[43][17] ) );
  NOR2_X1 U9235 ( .A1(n2502), .A2(n3013), .ZN(\mult_22/ab[46][20] ) );
  NOR2_X1 U9236 ( .A1(n2507), .A2(n3025), .ZN(\mult_22/ab[48][21] ) );
  NOR2_X1 U9237 ( .A1(n2429), .A2(n3023), .ZN(\mult_22/ab[47][8] ) );
  NOR2_X1 U9238 ( .A1(n2648), .A2(n2805), .ZN(\mult_22/ab[11][45] ) );
  NOR2_X1 U9239 ( .A1(n2496), .A2(n3000), .ZN(\mult_22/ab[44][19] ) );
  NOR2_X1 U9240 ( .A1(n2443), .A2(n3006), .ZN(\mult_22/ab[45][10] ) );
  NOR2_X1 U9241 ( .A1(n2460), .A2(n2994), .ZN(\mult_22/ab[43][13] ) );
  NOR2_X1 U9242 ( .A1(n2502), .A2(n3007), .ZN(\mult_22/ab[45][20] ) );
  NOR2_X1 U9243 ( .A1(n2636), .A2(n2799), .ZN(\mult_22/ab[10][43] ) );
  NOR2_X1 U9244 ( .A1(n2507), .A2(n3019), .ZN(\mult_22/ab[47][21] ) );
  NOR2_X1 U9245 ( .A1(n2513), .A2(n3043), .ZN(\mult_22/ab[51][22] ) );
  NOR2_X1 U9246 ( .A1(n2648), .A2(n2799), .ZN(\mult_22/ab[10][45] ) );
  NOR2_X1 U9247 ( .A1(n2472), .A2(n2988), .ZN(\mult_22/ab[42][15] ) );
  NOR2_X1 U9248 ( .A1(n2484), .A2(n2988), .ZN(\mult_22/ab[42][17] ) );
  NOR2_X1 U9249 ( .A1(n2513), .A2(n3037), .ZN(\mult_22/ab[50][22] ) );
  NOR2_X1 U9250 ( .A1(n2496), .A2(n2994), .ZN(\mult_22/ab[43][19] ) );
  NOR2_X1 U9251 ( .A1(n2646), .A2(n2835), .ZN(\mult_22/ab[16][44] ) );
  NOR2_X1 U9252 ( .A1(n2508), .A2(n3013), .ZN(\mult_22/ab[46][21] ) );
  NOR2_X1 U9253 ( .A1(n2417), .A2(n3035), .ZN(\mult_22/ab[49][6] ) );
  NOR2_X1 U9254 ( .A1(n2502), .A2(n3001), .ZN(\mult_22/ab[44][20] ) );
  NOR2_X1 U9255 ( .A1(n2454), .A2(n2994), .ZN(\mult_22/ab[43][12] ) );
  NOR2_X1 U9256 ( .A1(n2513), .A2(n3031), .ZN(\mult_22/ab[49][22] ) );
  NOR2_X1 U9257 ( .A1(n2659), .A2(n2799), .ZN(\mult_22/ab[10][46] ) );
  NOR2_X1 U9258 ( .A1(n2508), .A2(n3007), .ZN(\mult_22/ab[45][21] ) );
  NOR2_X1 U9259 ( .A1(n2513), .A2(n3025), .ZN(\mult_22/ab[48][22] ) );
  NOR2_X1 U9260 ( .A1(n2611), .A2(n2834), .ZN(\mult_22/ab[16][38] ) );
  NOR2_X1 U9261 ( .A1(n2648), .A2(n2823), .ZN(\mult_22/ab[14][45] ) );
  NOR2_X1 U9262 ( .A1(n2496), .A2(n2988), .ZN(\mult_22/ab[42][19] ) );
  NOR2_X1 U9263 ( .A1(n2616), .A2(n2822), .ZN(\mult_22/ab[14][39] ) );
  NOR2_X1 U9264 ( .A1(n2484), .A2(n2982), .ZN(\mult_22/ab[41][17] ) );
  NOR2_X1 U9265 ( .A1(n2513), .A2(n3019), .ZN(\mult_22/ab[47][22] ) );
  NOR2_X1 U9266 ( .A1(n2508), .A2(n3001), .ZN(\mult_22/ab[44][21] ) );
  NOR2_X1 U9267 ( .A1(n2443), .A2(n3000), .ZN(\mult_22/ab[44][10] ) );
  NOR2_X1 U9268 ( .A1(n2472), .A2(n2982), .ZN(\mult_22/ab[41][15] ) );
  NOR2_X1 U9269 ( .A1(n2430), .A2(n3017), .ZN(\mult_22/ab[46][8] ) );
  NOR2_X1 U9270 ( .A1(n2653), .A2(n2793), .ZN(\mult_22/ab[9][45] ) );
  NOR2_X1 U9271 ( .A1(n2592), .A2(n2882), .ZN(\mult_22/ab[24][35] ) );
  NOR2_X1 U9272 ( .A1(n2514), .A2(n3013), .ZN(\mult_22/ab[46][22] ) );
  NOR2_X1 U9273 ( .A1(n2519), .A2(n3037), .ZN(\mult_22/ab[50][23] ) );
  NOR2_X1 U9274 ( .A1(n2496), .A2(n2982), .ZN(\mult_22/ab[41][19] ) );
  NOR2_X1 U9275 ( .A1(n2508), .A2(n2995), .ZN(\mult_22/ab[43][21] ) );
  NOR2_X1 U9276 ( .A1(n2514), .A2(n3007), .ZN(\mult_22/ab[45][22] ) );
  NOR2_X1 U9277 ( .A1(n2599), .A2(n2858), .ZN(\mult_22/ab[20][36] ) );
  NOR2_X1 U9278 ( .A1(n2519), .A2(n3031), .ZN(\mult_22/ab[49][23] ) );
  NOR2_X1 U9279 ( .A1(n2454), .A2(n2988), .ZN(\mult_22/ab[42][12] ) );
  NOR2_X1 U9280 ( .A1(n2407), .A2(n3045), .ZN(\mult_22/ab[51][4] ) );
  NOR2_X1 U9281 ( .A1(n2519), .A2(n3025), .ZN(\mult_22/ab[48][23] ) );
  NOR2_X1 U9282 ( .A1(n2484), .A2(n2976), .ZN(\mult_22/ab[40][17] ) );
  NOR2_X1 U9283 ( .A1(n2514), .A2(n3001), .ZN(\mult_22/ab[44][22] ) );
  NOR2_X1 U9284 ( .A1(n2641), .A2(n2793), .ZN(\mult_22/ab[9][43] ) );
  NOR2_X1 U9285 ( .A1(n2417), .A2(n3029), .ZN(\mult_22/ab[48][6] ) );
  NOR2_X1 U9286 ( .A1(n2508), .A2(n2989), .ZN(\mult_22/ab[42][21] ) );
  NOR2_X1 U9287 ( .A1(n2519), .A2(n3019), .ZN(\mult_22/ab[47][23] ) );
  NOR2_X1 U9288 ( .A1(n2496), .A2(n2976), .ZN(\mult_22/ab[40][19] ) );
  NOR2_X1 U9289 ( .A1(n2648), .A2(n2829), .ZN(\mult_22/ab[15][45] ) );
  NOR2_X1 U9290 ( .A1(n2472), .A2(n2976), .ZN(\mult_22/ab[40][15] ) );
  NOR2_X1 U9291 ( .A1(n2520), .A2(n3013), .ZN(\mult_22/ab[46][23] ) );
  NOR2_X1 U9292 ( .A1(n2581), .A2(n2870), .ZN(\mult_22/ab[22][33] ) );
  NOR2_X1 U9293 ( .A1(n2514), .A2(n2995), .ZN(\mult_22/ab[43][22] ) );
  NOR2_X1 U9294 ( .A1(n2508), .A2(n2983), .ZN(\mult_22/ab[41][21] ) );
  NOR2_X1 U9295 ( .A1(n2442), .A2(n2994), .ZN(\mult_22/ab[43][10] ) );
  NOR2_X1 U9296 ( .A1(n2557), .A2(n2923), .ZN(\mult_22/ab[31][29] ) );
  NOR2_X1 U9297 ( .A1(n2611), .A2(n2828), .ZN(\mult_22/ab[15][38] ) );
  NOR2_X1 U9298 ( .A1(n2520), .A2(n3007), .ZN(\mult_22/ab[45][23] ) );
  NOR2_X1 U9299 ( .A1(n2605), .A2(n2852), .ZN(\mult_22/ab[19][37] ) );
  NOR2_X1 U9300 ( .A1(n2527), .A2(n3031), .ZN(\mult_22/ab[49][24] ) );
  NOR2_X1 U9301 ( .A1(n2616), .A2(n2816), .ZN(\mult_22/ab[13][39] ) );
  NOR2_X1 U9302 ( .A1(n2484), .A2(n2970), .ZN(\mult_22/ab[39][17] ) );
  NOR2_X1 U9303 ( .A1(n2658), .A2(n2817), .ZN(\mult_22/ab[13][46] ) );
  NOR2_X1 U9304 ( .A1(n2430), .A2(n3011), .ZN(\mult_22/ab[45][8] ) );
  NOR2_X1 U9305 ( .A1(n2587), .A2(n2870), .ZN(\mult_22/ab[22][34] ) );
  NOR2_X1 U9306 ( .A1(n2653), .A2(n2787), .ZN(\mult_22/ab[8][45] ) );
  NOR2_X1 U9307 ( .A1(n2496), .A2(n2970), .ZN(\mult_22/ab[39][19] ) );
  NOR2_X1 U9308 ( .A1(n2599), .A2(n2852), .ZN(\mult_22/ab[19][36] ) );
  NOR2_X1 U9309 ( .A1(n2520), .A2(n3001), .ZN(\mult_22/ab[44][23] ) );
  NOR2_X1 U9310 ( .A1(n2454), .A2(n2982), .ZN(\mult_22/ab[41][12] ) );
  NOR2_X1 U9311 ( .A1(n2527), .A2(n3025), .ZN(\mult_22/ab[48][24] ) );
  NOR2_X1 U9312 ( .A1(n2587), .A2(n2864), .ZN(\mult_22/ab[21][34] ) );
  NOR2_X1 U9313 ( .A1(n2508), .A2(n2977), .ZN(\mult_22/ab[40][21] ) );
  NOR2_X1 U9314 ( .A1(n2563), .A2(n2923), .ZN(\mult_22/ab[31][30] ) );
  NOR2_X1 U9315 ( .A1(n2407), .A2(n3039), .ZN(\mult_22/ab[50][4] ) );
  NOR2_X1 U9316 ( .A1(n2573), .A2(n2894), .ZN(\mult_22/ab[26][32] ) );
  NOR2_X1 U9317 ( .A1(n2581), .A2(n2864), .ZN(\mult_22/ab[21][33] ) );
  NOR2_X1 U9318 ( .A1(n2514), .A2(n2983), .ZN(\mult_22/ab[41][22] ) );
  NOR2_X1 U9319 ( .A1(n2527), .A2(n3019), .ZN(\mult_22/ab[47][24] ) );
  NOR2_X1 U9320 ( .A1(n2520), .A2(n2995), .ZN(\mult_22/ab[43][23] ) );
  NOR2_X1 U9321 ( .A1(n2472), .A2(n2970), .ZN(\mult_22/ab[39][15] ) );
  NOR2_X1 U9322 ( .A1(n2417), .A2(n3023), .ZN(\mult_22/ab[47][6] ) );
  NOR2_X1 U9323 ( .A1(n2666), .A2(n2793), .ZN(\mult_22/ab[9][48] ) );
  NOR2_X1 U9324 ( .A1(n2527), .A2(n3013), .ZN(\mult_22/ab[46][24] ) );
  NOR2_X1 U9325 ( .A1(n2605), .A2(n2846), .ZN(\mult_22/ab[18][37] ) );
  NOR2_X1 U9326 ( .A1(n2520), .A2(n2989), .ZN(\mult_22/ab[42][23] ) );
  NOR2_X1 U9327 ( .A1(n2527), .A2(n3007), .ZN(\mult_22/ab[45][24] ) );
  NOR2_X1 U9328 ( .A1(n2658), .A2(n2823), .ZN(\mult_22/ab[14][46] ) );
  NOR2_X1 U9329 ( .A1(n2593), .A2(n2864), .ZN(\mult_22/ab[21][35] ) );
  NOR2_X1 U9330 ( .A1(n2508), .A2(n2971), .ZN(\mult_22/ab[39][21] ) );
  NOR2_X1 U9331 ( .A1(n2641), .A2(n2787), .ZN(\mult_22/ab[8][43] ) );
  NOR2_X1 U9332 ( .A1(n2563), .A2(n2917), .ZN(\mult_22/ab[30][30] ) );
  NOR2_X1 U9333 ( .A1(n2599), .A2(n2846), .ZN(\mult_22/ab[18][36] ) );
  NOR2_X1 U9334 ( .A1(n2611), .A2(n2822), .ZN(\mult_22/ab[14][38] ) );
  NOR2_X1 U9335 ( .A1(n2527), .A2(n3001), .ZN(\mult_22/ab[44][24] ) );
  NOR2_X1 U9336 ( .A1(n2442), .A2(n2988), .ZN(\mult_22/ab[42][10] ) );
  NOR2_X1 U9337 ( .A1(n2694), .A2(n2775), .ZN(\mult_22/ab[6][52] ) );
  NOR2_X1 U9338 ( .A1(n2520), .A2(n2983), .ZN(\mult_22/ab[41][23] ) );
  NOR2_X1 U9339 ( .A1(n2496), .A2(n2964), .ZN(\mult_22/ab[38][19] ) );
  NOR2_X1 U9340 ( .A1(n2484), .A2(n2964), .ZN(\mult_22/ab[38][17] ) );
  NOR2_X1 U9341 ( .A1(n2617), .A2(n2810), .ZN(\mult_22/ab[12][39] ) );
  NOR2_X1 U9342 ( .A1(n2538), .A2(n2953), .ZN(\mult_22/ab[36][26] ) );
  NOR2_X1 U9343 ( .A1(n2526), .A2(n2971), .ZN(\mult_22/ab[39][24] ) );
  NOR2_X1 U9344 ( .A1(n2538), .A2(n2959), .ZN(\mult_22/ab[37][26] ) );
  NOR2_X1 U9345 ( .A1(n2526), .A2(n2977), .ZN(\mult_22/ab[40][24] ) );
  NOR2_X1 U9346 ( .A1(n2538), .A2(n2965), .ZN(\mult_22/ab[38][26] ) );
  NOR2_X1 U9347 ( .A1(n2526), .A2(n2983), .ZN(\mult_22/ab[41][24] ) );
  NOR2_X1 U9348 ( .A1(n2538), .A2(n2971), .ZN(\mult_22/ab[39][26] ) );
  NOR2_X1 U9349 ( .A1(n2532), .A2(n2953), .ZN(\mult_22/ab[36][25] ) );
  NOR2_X1 U9350 ( .A1(n2532), .A2(n2959), .ZN(\mult_22/ab[37][25] ) );
  NOR2_X1 U9351 ( .A1(n2520), .A2(n2965), .ZN(\mult_22/ab[38][23] ) );
  NOR2_X1 U9352 ( .A1(n2520), .A2(n2971), .ZN(\mult_22/ab[39][23] ) );
  NOR2_X1 U9353 ( .A1(n2520), .A2(n2977), .ZN(\mult_22/ab[40][23] ) );
  NOR2_X1 U9354 ( .A1(n2532), .A2(n2965), .ZN(\mult_22/ab[38][25] ) );
  NOR2_X1 U9355 ( .A1(n2532), .A2(n2971), .ZN(\mult_22/ab[39][25] ) );
  NOR2_X1 U9356 ( .A1(n2532), .A2(n2977), .ZN(\mult_22/ab[40][25] ) );
  NOR2_X1 U9357 ( .A1(n2538), .A2(n2977), .ZN(\mult_22/ab[40][26] ) );
  NOR2_X1 U9358 ( .A1(n2544), .A2(n2953), .ZN(\mult_22/ab[36][27] ) );
  NOR2_X1 U9359 ( .A1(n2544), .A2(n2959), .ZN(\mult_22/ab[37][27] ) );
  NOR2_X1 U9360 ( .A1(n2684), .A2(n2787), .ZN(\mult_22/ab[8][51] ) );
  NOR2_X1 U9361 ( .A1(n2665), .A2(n2811), .ZN(\mult_22/ab[12][47] ) );
  NOR2_X1 U9362 ( .A1(n2544), .A2(n2965), .ZN(\mult_22/ab[38][27] ) );
  NOR2_X1 U9363 ( .A1(n2526), .A2(n2989), .ZN(\mult_22/ab[42][24] ) );
  NOR2_X1 U9364 ( .A1(n2532), .A2(n2983), .ZN(\mult_22/ab[41][25] ) );
  NOR2_X1 U9365 ( .A1(n2573), .A2(n2906), .ZN(\mult_22/ab[28][32] ) );
  NOR2_X1 U9366 ( .A1(n2676), .A2(n2781), .ZN(\mult_22/ab[7][49] ) );
  NOR2_X1 U9367 ( .A1(n2544), .A2(n2971), .ZN(\mult_22/ab[39][27] ) );
  NOR2_X1 U9368 ( .A1(n2587), .A2(n2858), .ZN(\mult_22/ab[20][34] ) );
  NOR2_X1 U9369 ( .A1(n2569), .A2(n2912), .ZN(\mult_22/ab[29][31] ) );
  NOR2_X1 U9370 ( .A1(n2532), .A2(n2989), .ZN(\mult_22/ab[42][25] ) );
  NOR2_X1 U9371 ( .A1(n2671), .A2(n2805), .ZN(\mult_22/ab[11][48] ) );
  NOR2_X1 U9372 ( .A1(n2694), .A2(n2781), .ZN(\mult_22/ab[7][52] ) );
  NOR2_X1 U9373 ( .A1(n2593), .A2(n2858), .ZN(\mult_22/ab[20][35] ) );
  NOR2_X1 U9374 ( .A1(n2544), .A2(n2977), .ZN(\mult_22/ab[40][27] ) );
  NOR2_X1 U9375 ( .A1(n2580), .A2(n2906), .ZN(\mult_22/ab[28][33] ) );
  NOR2_X1 U9376 ( .A1(n2569), .A2(n2918), .ZN(\mult_22/ab[30][31] ) );
  NOR2_X1 U9377 ( .A1(n2573), .A2(n2912), .ZN(\mult_22/ab[29][32] ) );
  NOR2_X1 U9378 ( .A1(n2665), .A2(n2805), .ZN(\mult_22/ab[11][47] ) );
  NOR2_X1 U9379 ( .A1(n2696), .A2(n2763), .ZN(\mult_22/ab[4][53] ) );
  NOR2_X1 U9380 ( .A1(n2526), .A2(n2995), .ZN(\mult_22/ab[43][24] ) );
  NOR2_X1 U9381 ( .A1(n2538), .A2(n2983), .ZN(\mult_22/ab[41][26] ) );
  NOR2_X1 U9382 ( .A1(n2598), .A2(n2888), .ZN(\mult_22/ab[25][36] ) );
  NOR2_X1 U9383 ( .A1(n2551), .A2(n2947), .ZN(\mult_22/ab[35][28] ) );
  NOR2_X1 U9384 ( .A1(n2550), .A2(n2953), .ZN(\mult_22/ab[36][28] ) );
  NOR2_X1 U9385 ( .A1(n2550), .A2(n2959), .ZN(\mult_22/ab[37][28] ) );
  NOR2_X1 U9386 ( .A1(n2430), .A2(n3005), .ZN(\mult_22/ab[44][8] ) );
  NOR2_X1 U9387 ( .A1(n2550), .A2(n2965), .ZN(\mult_22/ab[38][28] ) );
  NOR2_X1 U9388 ( .A1(n2611), .A2(n2804), .ZN(\mult_22/ab[11][38] ) );
  NOR2_X1 U9389 ( .A1(n2599), .A2(n2840), .ZN(\mult_22/ab[17][36] ) );
  NOR2_X1 U9390 ( .A1(n2612), .A2(n2786), .ZN(\mult_22/ab[8][39] ) );
  NOR2_X1 U9391 ( .A1(n2612), .A2(n2792), .ZN(\mult_22/ab[9][39] ) );
  NOR2_X1 U9392 ( .A1(n2617), .A2(n2798), .ZN(\mult_22/ab[10][39] ) );
  NOR2_X1 U9393 ( .A1(n2617), .A2(n2804), .ZN(\mult_22/ab[11][39] ) );
  NOR2_X1 U9394 ( .A1(n2606), .A2(n2804), .ZN(\mult_22/ab[11][37] ) );
  NOR2_X1 U9395 ( .A1(n2605), .A2(n2810), .ZN(\mult_22/ab[12][37] ) );
  NOR2_X1 U9396 ( .A1(n2605), .A2(n2816), .ZN(\mult_22/ab[13][37] ) );
  NOR2_X1 U9397 ( .A1(n2605), .A2(n2822), .ZN(\mult_22/ab[14][37] ) );
  NOR2_X1 U9398 ( .A1(n2593), .A2(n2822), .ZN(\mult_22/ab[14][35] ) );
  NOR2_X1 U9399 ( .A1(n2605), .A2(n2828), .ZN(\mult_22/ab[15][37] ) );
  NOR2_X1 U9400 ( .A1(n2593), .A2(n2828), .ZN(\mult_22/ab[15][35] ) );
  NOR2_X1 U9401 ( .A1(n2593), .A2(n2834), .ZN(\mult_22/ab[16][35] ) );
  NOR2_X1 U9402 ( .A1(n2581), .A2(n2840), .ZN(\mult_22/ab[17][33] ) );
  NOR2_X1 U9403 ( .A1(n2593), .A2(n2840), .ZN(\mult_22/ab[17][35] ) );
  NOR2_X1 U9404 ( .A1(n2581), .A2(n2846), .ZN(\mult_22/ab[18][33] ) );
  NOR2_X1 U9405 ( .A1(n2593), .A2(n2846), .ZN(\mult_22/ab[18][35] ) );
  NOR2_X1 U9406 ( .A1(n2581), .A2(n2852), .ZN(\mult_22/ab[19][33] ) );
  NOR2_X1 U9407 ( .A1(n2581), .A2(n2858), .ZN(\mult_22/ab[20][33] ) );
  NOR2_X1 U9408 ( .A1(n2612), .A2(n2780), .ZN(\mult_22/ab[7][39] ) );
  NOR2_X1 U9409 ( .A1(n2606), .A2(n2798), .ZN(\mult_22/ab[10][37] ) );
  NOR2_X1 U9410 ( .A1(n2593), .A2(n2816), .ZN(\mult_22/ab[13][35] ) );
  NOR2_X1 U9411 ( .A1(n2581), .A2(n2834), .ZN(\mult_22/ab[16][33] ) );
  NOR2_X1 U9412 ( .A1(n2605), .A2(n2834), .ZN(\mult_22/ab[16][37] ) );
  NOR2_X1 U9413 ( .A1(n2593), .A2(n2852), .ZN(\mult_22/ab[19][35] ) );
  NOR2_X1 U9414 ( .A1(n2612), .A2(n2774), .ZN(\mult_22/ab[6][39] ) );
  NOR2_X1 U9415 ( .A1(n2601), .A2(n2792), .ZN(\mult_22/ab[9][37] ) );
  NOR2_X1 U9416 ( .A1(n2593), .A2(n2810), .ZN(\mult_22/ab[12][35] ) );
  NOR2_X1 U9417 ( .A1(n2581), .A2(n2828), .ZN(\mult_22/ab[15][33] ) );
  NOR2_X1 U9418 ( .A1(n2601), .A2(n2786), .ZN(\mult_22/ab[8][37] ) );
  NOR2_X1 U9419 ( .A1(n2594), .A2(n2804), .ZN(\mult_22/ab[11][35] ) );
  NOR2_X1 U9420 ( .A1(n2581), .A2(n2822), .ZN(\mult_22/ab[14][33] ) );
  NOR2_X1 U9421 ( .A1(n2605), .A2(n2840), .ZN(\mult_22/ab[17][37] ) );
  NOR2_X1 U9422 ( .A1(n2594), .A2(n2798), .ZN(\mult_22/ab[10][35] ) );
  NOR2_X1 U9423 ( .A1(n2582), .A2(n2816), .ZN(\mult_22/ab[13][33] ) );
  NOR2_X1 U9424 ( .A1(n2582), .A2(n2810), .ZN(\mult_22/ab[12][33] ) );
  NOR2_X1 U9425 ( .A1(n2677), .A2(n2787), .ZN(\mult_22/ab[8][49] ) );
  NOR2_X1 U9426 ( .A1(n2640), .A2(n2781), .ZN(\mult_22/ab[7][43] ) );
  NOR2_X1 U9427 ( .A1(n2607), .A2(n2774), .ZN(\mult_22/ab[6][38] ) );
  NOR2_X1 U9428 ( .A1(n2607), .A2(n2768), .ZN(\mult_22/ab[5][38] ) );
  NOR2_X1 U9429 ( .A1(n2595), .A2(n2786), .ZN(\mult_22/ab[8][36] ) );
  NOR2_X1 U9430 ( .A1(n2595), .A2(n2780), .ZN(\mult_22/ab[7][36] ) );
  NOR2_X1 U9431 ( .A1(n2588), .A2(n2798), .ZN(\mult_22/ab[10][34] ) );
  NOR2_X1 U9432 ( .A1(n2583), .A2(n2792), .ZN(\mult_22/ab[9][34] ) );
  NOR2_X1 U9433 ( .A1(n2652), .A2(n2781), .ZN(\mult_22/ab[7][45] ) );
  NOR2_X1 U9434 ( .A1(n2652), .A2(n2775), .ZN(\mult_22/ab[6][45] ) );
  NOR2_X1 U9435 ( .A1(n2652), .A2(n2769), .ZN(\mult_22/ab[5][45] ) );
  NOR2_X1 U9436 ( .A1(n2640), .A2(n2775), .ZN(\mult_22/ab[6][43] ) );
  NOR2_X1 U9437 ( .A1(n2580), .A2(n2912), .ZN(\mult_22/ab[29][33] ) );
  NOR2_X1 U9438 ( .A1(n2569), .A2(n2924), .ZN(\mult_22/ab[31][31] ) );
  NOR2_X1 U9439 ( .A1(n2557), .A2(n2935), .ZN(\mult_22/ab[33][29] ) );
  NOR2_X1 U9440 ( .A1(n2569), .A2(n2930), .ZN(\mult_22/ab[32][31] ) );
  NOR2_X1 U9441 ( .A1(n2557), .A2(n2941), .ZN(\mult_22/ab[34][29] ) );
  NOR2_X1 U9442 ( .A1(n2557), .A2(n2947), .ZN(\mult_22/ab[35][29] ) );
  NOR2_X1 U9443 ( .A1(n2592), .A2(n2900), .ZN(\mult_22/ab[27][35] ) );
  NOR2_X1 U9444 ( .A1(n2580), .A2(n2918), .ZN(\mult_22/ab[30][33] ) );
  NOR2_X1 U9445 ( .A1(n2569), .A2(n2935), .ZN(\mult_22/ab[33][31] ) );
  NOR2_X1 U9446 ( .A1(n2640), .A2(n2769), .ZN(\mult_22/ab[5][43] ) );
  NOR2_X1 U9447 ( .A1(n2592), .A2(n2906), .ZN(\mult_22/ab[28][35] ) );
  NOR2_X1 U9448 ( .A1(n2580), .A2(n2924), .ZN(\mult_22/ab[31][33] ) );
  NOR2_X1 U9449 ( .A1(n2604), .A2(n2888), .ZN(\mult_22/ab[25][37] ) );
  NOR2_X1 U9450 ( .A1(n2592), .A2(n2912), .ZN(\mult_22/ab[29][35] ) );
  NOR2_X1 U9451 ( .A1(n2604), .A2(n2894), .ZN(\mult_22/ab[26][37] ) );
  NOR2_X1 U9452 ( .A1(n2604), .A2(n2900), .ZN(\mult_22/ab[27][37] ) );
  NOR2_X1 U9453 ( .A1(n2563), .A2(n2929), .ZN(\mult_22/ab[32][30] ) );
  NOR2_X1 U9454 ( .A1(n2573), .A2(n2918), .ZN(\mult_22/ab[30][32] ) );
  NOR2_X1 U9455 ( .A1(n2563), .A2(n2935), .ZN(\mult_22/ab[33][30] ) );
  NOR2_X1 U9456 ( .A1(n2573), .A2(n2924), .ZN(\mult_22/ab[31][32] ) );
  NOR2_X1 U9457 ( .A1(n2563), .A2(n2941), .ZN(\mult_22/ab[34][30] ) );
  NOR2_X1 U9458 ( .A1(n2586), .A2(n2906), .ZN(\mult_22/ab[28][34] ) );
  NOR2_X1 U9459 ( .A1(n2573), .A2(n2930), .ZN(\mult_22/ab[32][32] ) );
  NOR2_X1 U9460 ( .A1(n2563), .A2(n2947), .ZN(\mult_22/ab[35][30] ) );
  NOR2_X1 U9461 ( .A1(n2586), .A2(n2912), .ZN(\mult_22/ab[29][34] ) );
  NOR2_X1 U9462 ( .A1(n2556), .A2(n2953), .ZN(\mult_22/ab[36][29] ) );
  NOR2_X1 U9463 ( .A1(n2573), .A2(n2936), .ZN(\mult_22/ab[33][32] ) );
  NOR2_X1 U9464 ( .A1(n2586), .A2(n2918), .ZN(\mult_22/ab[30][34] ) );
  NOR2_X1 U9465 ( .A1(n2569), .A2(n2942), .ZN(\mult_22/ab[34][31] ) );
  NOR2_X1 U9466 ( .A1(n2586), .A2(n2924), .ZN(\mult_22/ab[31][34] ) );
  NOR2_X1 U9467 ( .A1(n2580), .A2(n2930), .ZN(\mult_22/ab[32][33] ) );
  NOR2_X1 U9468 ( .A1(n2592), .A2(n2918), .ZN(\mult_22/ab[30][35] ) );
  NOR2_X1 U9469 ( .A1(n2604), .A2(n2906), .ZN(\mult_22/ab[28][37] ) );
  NOR2_X1 U9470 ( .A1(n2581), .A2(n2882), .ZN(\mult_22/ab[24][33] ) );
  NOR2_X1 U9471 ( .A1(n2598), .A2(n2894), .ZN(\mult_22/ab[26][36] ) );
  NOR2_X1 U9472 ( .A1(n2598), .A2(n2900), .ZN(\mult_22/ab[27][36] ) );
  NOR2_X1 U9473 ( .A1(n2598), .A2(n2906), .ZN(\mult_22/ab[28][36] ) );
  NOR2_X1 U9474 ( .A1(n2598), .A2(n2912), .ZN(\mult_22/ab[29][36] ) );
  NOR2_X1 U9475 ( .A1(n2651), .A2(n2763), .ZN(\mult_22/ab[4][45] ) );
  NOR2_X1 U9476 ( .A1(n2550), .A2(n2971), .ZN(\mult_22/ab[39][28] ) );
  NOR2_X1 U9477 ( .A1(n2701), .A2(n2764), .ZN(\mult_22/ab[4][54] ) );
  NOR2_X1 U9478 ( .A1(n2610), .A2(n2888), .ZN(\mult_22/ab[25][38] ) );
  NOR2_X1 U9479 ( .A1(n2610), .A2(n2894), .ZN(\mult_22/ab[26][38] ) );
  NOR2_X1 U9480 ( .A1(n2610), .A2(n2900), .ZN(\mult_22/ab[27][38] ) );
  NOR2_X1 U9481 ( .A1(n2650), .A2(n2757), .ZN(\mult_22/ab[3][45] ) );
  NOR2_X1 U9482 ( .A1(n2587), .A2(n2876), .ZN(\mult_22/ab[23][34] ) );
  NOR2_X1 U9483 ( .A1(n2562), .A2(n2953), .ZN(\mult_22/ab[36][30] ) );
  NOR2_X1 U9484 ( .A1(n2574), .A2(n2942), .ZN(\mult_22/ab[34][32] ) );
  NOR2_X1 U9485 ( .A1(n2586), .A2(n2930), .ZN(\mult_22/ab[32][34] ) );
  NOR2_X1 U9486 ( .A1(n2556), .A2(n2959), .ZN(\mult_22/ab[37][29] ) );
  NOR2_X1 U9487 ( .A1(n2569), .A2(n2948), .ZN(\mult_22/ab[35][31] ) );
  NOR2_X1 U9488 ( .A1(n2580), .A2(n2936), .ZN(\mult_22/ab[33][33] ) );
  NOR2_X1 U9489 ( .A1(n2592), .A2(n2924), .ZN(\mult_22/ab[31][35] ) );
  NOR2_X1 U9490 ( .A1(n2604), .A2(n2912), .ZN(\mult_22/ab[29][37] ) );
  NOR2_X1 U9491 ( .A1(n2598), .A2(n2918), .ZN(\mult_22/ab[30][36] ) );
  NOR2_X1 U9492 ( .A1(n2610), .A2(n2906), .ZN(\mult_22/ab[28][38] ) );
  NOR2_X1 U9493 ( .A1(n2532), .A2(n2995), .ZN(\mult_22/ab[43][25] ) );
  NOR2_X1 U9494 ( .A1(n2544), .A2(n2983), .ZN(\mult_22/ab[41][27] ) );
  NOR2_X1 U9495 ( .A1(n2675), .A2(n2763), .ZN(\mult_22/ab[4][49] ) );
  NOR2_X1 U9496 ( .A1(n2556), .A2(n2965), .ZN(\mult_22/ab[38][29] ) );
  NOR2_X1 U9497 ( .A1(n2569), .A2(n2954), .ZN(\mult_22/ab[36][31] ) );
  NOR2_X1 U9498 ( .A1(n2580), .A2(n2942), .ZN(\mult_22/ab[34][33] ) );
  NOR2_X1 U9499 ( .A1(n2592), .A2(n2930), .ZN(\mult_22/ab[32][35] ) );
  NOR2_X1 U9500 ( .A1(n2604), .A2(n2918), .ZN(\mult_22/ab[30][37] ) );
  NOR2_X1 U9501 ( .A1(n2538), .A2(n2989), .ZN(\mult_22/ab[42][26] ) );
  NOR2_X1 U9502 ( .A1(n2684), .A2(n2793), .ZN(\mult_22/ab[9][51] ) );
  NOR2_X1 U9503 ( .A1(n2672), .A2(n2805), .ZN(\mult_22/ab[11][49] ) );
  NOR2_X1 U9504 ( .A1(n2665), .A2(n2817), .ZN(\mult_22/ab[13][47] ) );
  NOR2_X1 U9505 ( .A1(n2614), .A2(n2756), .ZN(\mult_22/ab[3][39] ) );
  NOR2_X1 U9506 ( .A1(n2601), .A2(n2768), .ZN(\mult_22/ab[5][37] ) );
  NOR2_X1 U9507 ( .A1(n2589), .A2(n2780), .ZN(\mult_22/ab[7][35] ) );
  NOR2_X1 U9508 ( .A1(n2577), .A2(n2792), .ZN(\mult_22/ab[9][33] ) );
  NOR2_X1 U9509 ( .A1(n2729), .A2(n2770), .ZN(\mult_22/ab[5][59] ) );
  NOR2_X1 U9510 ( .A1(n2718), .A2(n2782), .ZN(\mult_22/ab[7][57] ) );
  NOR2_X1 U9511 ( .A1(n2708), .A2(n2794), .ZN(\mult_22/ab[9][55] ) );
  NOR2_X1 U9512 ( .A1(n2695), .A2(n2805), .ZN(\mult_22/ab[11][53] ) );
  NOR2_X1 U9513 ( .A1(n2689), .A2(n2817), .ZN(\mult_22/ab[13][51] ) );
  NOR2_X1 U9514 ( .A1(n2672), .A2(n2829), .ZN(\mult_22/ab[15][49] ) );
  NOR2_X1 U9515 ( .A1(n2664), .A2(n2841), .ZN(\mult_22/ab[17][47] ) );
  NOR2_X1 U9516 ( .A1(n2648), .A2(n2853), .ZN(\mult_22/ab[19][45] ) );
  NOR2_X1 U9517 ( .A1(n2636), .A2(n2865), .ZN(\mult_22/ab[21][43] ) );
  NOR2_X1 U9518 ( .A1(n2625), .A2(n2876), .ZN(\mult_22/ab[23][41] ) );
  NOR2_X1 U9519 ( .A1(n2615), .A2(n2888), .ZN(\mult_22/ab[25][39] ) );
  NOR2_X1 U9520 ( .A1(n2716), .A2(n2788), .ZN(\mult_22/ab[8][57] ) );
  NOR2_X1 U9521 ( .A1(n2695), .A2(n2812), .ZN(\mult_22/ab[12][53] ) );
  NOR2_X1 U9522 ( .A1(n2689), .A2(n2823), .ZN(\mult_22/ab[14][51] ) );
  NOR2_X1 U9523 ( .A1(n2672), .A2(n2835), .ZN(\mult_22/ab[16][49] ) );
  NOR2_X1 U9524 ( .A1(n2664), .A2(n2847), .ZN(\mult_22/ab[18][47] ) );
  NOR2_X1 U9525 ( .A1(n2648), .A2(n2859), .ZN(\mult_22/ab[20][45] ) );
  NOR2_X1 U9526 ( .A1(n2637), .A2(n2871), .ZN(\mult_22/ab[22][43] ) );
  NOR2_X1 U9527 ( .A1(n2625), .A2(n2882), .ZN(\mult_22/ab[24][41] ) );
  NOR2_X1 U9528 ( .A1(n2615), .A2(n2894), .ZN(\mult_22/ab[26][39] ) );
  NOR2_X1 U9529 ( .A1(n2730), .A2(n2776), .ZN(\mult_22/ab[6][59] ) );
  NOR2_X1 U9530 ( .A1(n2545), .A2(n2935), .ZN(\mult_22/ab[33][27] ) );
  NOR2_X1 U9531 ( .A1(n2533), .A2(n2947), .ZN(\mult_22/ab[35][25] ) );
  NOR2_X1 U9532 ( .A1(n2520), .A2(n2959), .ZN(\mult_22/ab[37][23] ) );
  NOR2_X1 U9533 ( .A1(n2694), .A2(n2787), .ZN(\mult_22/ab[8][52] ) );
  NOR2_X1 U9534 ( .A1(n2683), .A2(n2799), .ZN(\mult_22/ab[10][50] ) );
  NOR2_X1 U9535 ( .A1(n2671), .A2(n2811), .ZN(\mult_22/ab[12][48] ) );
  NOR2_X1 U9536 ( .A1(n2734), .A2(n2764), .ZN(\mult_22/ab[4][60] ) );
  NOR2_X1 U9537 ( .A1(n2723), .A2(n2776), .ZN(\mult_22/ab[6][58] ) );
  NOR2_X1 U9538 ( .A1(n2723), .A2(n2782), .ZN(\mult_22/ab[7][58] ) );
  NOR2_X1 U9539 ( .A1(n2705), .A2(n2806), .ZN(\mult_22/ab[11][54] ) );
  NOR2_X1 U9540 ( .A1(n2690), .A2(n2811), .ZN(\mult_22/ab[12][52] ) );
  NOR2_X1 U9541 ( .A1(n2690), .A2(n2817), .ZN(\mult_22/ab[13][52] ) );
  NOR2_X1 U9542 ( .A1(n2682), .A2(n2823), .ZN(\mult_22/ab[14][50] ) );
  NOR2_X1 U9543 ( .A1(n2682), .A2(n2829), .ZN(\mult_22/ab[15][50] ) );
  NOR2_X1 U9544 ( .A1(n2670), .A2(n2835), .ZN(\mult_22/ab[16][48] ) );
  NOR2_X1 U9545 ( .A1(n2670), .A2(n2841), .ZN(\mult_22/ab[17][48] ) );
  NOR2_X1 U9546 ( .A1(n2658), .A2(n2847), .ZN(\mult_22/ab[18][46] ) );
  NOR2_X1 U9547 ( .A1(n2658), .A2(n2853), .ZN(\mult_22/ab[19][46] ) );
  NOR2_X1 U9548 ( .A1(n2646), .A2(n2859), .ZN(\mult_22/ab[20][44] ) );
  NOR2_X1 U9549 ( .A1(n2646), .A2(n2865), .ZN(\mult_22/ab[21][44] ) );
  NOR2_X1 U9550 ( .A1(n2634), .A2(n2870), .ZN(\mult_22/ab[22][42] ) );
  NOR2_X1 U9551 ( .A1(n2634), .A2(n2876), .ZN(\mult_22/ab[23][42] ) );
  NOR2_X1 U9552 ( .A1(n2622), .A2(n2882), .ZN(\mult_22/ab[24][40] ) );
  NOR2_X1 U9553 ( .A1(n2621), .A2(n2888), .ZN(\mult_22/ab[25][40] ) );
  NOR2_X1 U9554 ( .A1(n2562), .A2(n2959), .ZN(\mult_22/ab[37][30] ) );
  NOR2_X1 U9555 ( .A1(n2574), .A2(n2948), .ZN(\mult_22/ab[35][32] ) );
  NOR2_X1 U9556 ( .A1(n2586), .A2(n2936), .ZN(\mult_22/ab[33][34] ) );
  NOR2_X1 U9557 ( .A1(n2581), .A2(n2888), .ZN(\mult_22/ab[25][33] ) );
  NOR2_X1 U9558 ( .A1(n2580), .A2(n2894), .ZN(\mult_22/ab[26][33] ) );
  NOR2_X1 U9559 ( .A1(n2569), .A2(n2905), .ZN(\mult_22/ab[28][31] ) );
  NOR2_X1 U9560 ( .A1(n2598), .A2(n2924), .ZN(\mult_22/ab[31][36] ) );
  NOR2_X1 U9561 ( .A1(n2711), .A2(n2806), .ZN(\mult_22/ab[11][55] ) );
  NOR2_X1 U9562 ( .A1(n2367), .A2(n2818), .ZN(\mult_22/ab[13][53] ) );
  NOR2_X1 U9563 ( .A1(n2688), .A2(n2829), .ZN(\mult_22/ab[15][51] ) );
  NOR2_X1 U9564 ( .A1(n2672), .A2(n2841), .ZN(\mult_22/ab[17][49] ) );
  NOR2_X1 U9565 ( .A1(n2664), .A2(n2853), .ZN(\mult_22/ab[19][47] ) );
  NOR2_X1 U9566 ( .A1(n2648), .A2(n2865), .ZN(\mult_22/ab[21][45] ) );
  NOR2_X1 U9567 ( .A1(n2637), .A2(n2877), .ZN(\mult_22/ab[23][43] ) );
  NOR2_X1 U9568 ( .A1(n2625), .A2(n2888), .ZN(\mult_22/ab[25][41] ) );
  NOR2_X1 U9569 ( .A1(n2615), .A2(n2900), .ZN(\mult_22/ab[27][39] ) );
  NOR2_X1 U9570 ( .A1(n2716), .A2(n2794), .ZN(\mult_22/ab[9][57] ) );
  NOR2_X1 U9571 ( .A1(n2725), .A2(n2782), .ZN(\mult_22/ab[7][59] ) );
  NOR2_X1 U9572 ( .A1(n2741), .A2(n2758), .ZN(\mult_22/ab[3][61] ) );
  NOR2_X1 U9573 ( .A1(n2610), .A2(n2912), .ZN(\mult_22/ab[29][38] ) );
  NOR2_X1 U9574 ( .A1(n2735), .A2(n2770), .ZN(\mult_22/ab[5][60] ) );
  NOR2_X1 U9575 ( .A1(n2705), .A2(n2812), .ZN(\mult_22/ab[12][54] ) );
  NOR2_X1 U9576 ( .A1(n2690), .A2(n2823), .ZN(\mult_22/ab[14][52] ) );
  NOR2_X1 U9577 ( .A1(n2682), .A2(n2835), .ZN(\mult_22/ab[16][50] ) );
  NOR2_X1 U9578 ( .A1(n2670), .A2(n2847), .ZN(\mult_22/ab[18][48] ) );
  NOR2_X1 U9579 ( .A1(n2658), .A2(n2859), .ZN(\mult_22/ab[20][46] ) );
  NOR2_X1 U9580 ( .A1(n2646), .A2(n2871), .ZN(\mult_22/ab[22][44] ) );
  NOR2_X1 U9581 ( .A1(n2634), .A2(n2882), .ZN(\mult_22/ab[24][42] ) );
  NOR2_X1 U9582 ( .A1(n2621), .A2(n2894), .ZN(\mult_22/ab[26][40] ) );
  NOR2_X1 U9583 ( .A1(n2724), .A2(n2788), .ZN(\mult_22/ab[8][58] ) );
  NOR2_X1 U9584 ( .A1(n2723), .A2(n2770), .ZN(\mult_22/ab[5][58] ) );
  NOR2_X1 U9585 ( .A1(n2699), .A2(n2824), .ZN(\mult_22/ab[14][53] ) );
  NOR2_X1 U9586 ( .A1(n2688), .A2(n2835), .ZN(\mult_22/ab[16][51] ) );
  NOR2_X1 U9587 ( .A1(n2672), .A2(n2847), .ZN(\mult_22/ab[18][49] ) );
  NOR2_X1 U9588 ( .A1(n2664), .A2(n2859), .ZN(\mult_22/ab[20][47] ) );
  NOR2_X1 U9589 ( .A1(n2649), .A2(n2871), .ZN(\mult_22/ab[22][45] ) );
  NOR2_X1 U9590 ( .A1(n2637), .A2(n2883), .ZN(\mult_22/ab[24][43] ) );
  NOR2_X1 U9591 ( .A1(n2625), .A2(n2894), .ZN(\mult_22/ab[26][41] ) );
  NOR2_X1 U9592 ( .A1(n2615), .A2(n2906), .ZN(\mult_22/ab[28][39] ) );
  NOR2_X1 U9593 ( .A1(n2711), .A2(n2812), .ZN(\mult_22/ab[12][55] ) );
  NOR2_X1 U9594 ( .A1(n2716), .A2(n2800), .ZN(\mult_22/ab[10][57] ) );
  NOR2_X1 U9595 ( .A1(n2726), .A2(n2788), .ZN(\mult_22/ab[8][59] ) );
  NOR2_X1 U9596 ( .A1(n2735), .A2(n2776), .ZN(\mult_22/ab[6][60] ) );
  NOR2_X1 U9597 ( .A1(n2609), .A2(n2756), .ZN(\mult_22/ab[3][38] ) );
  NOR2_X1 U9598 ( .A1(n2595), .A2(n2768), .ZN(\mult_22/ab[5][36] ) );
  NOR2_X1 U9599 ( .A1(n2583), .A2(n2780), .ZN(\mult_22/ab[7][34] ) );
  NOR2_X1 U9600 ( .A1(n2728), .A2(n2764), .ZN(\mult_22/ab[4][59] ) );
  NOR2_X1 U9601 ( .A1(n2718), .A2(n2776), .ZN(\mult_22/ab[6][57] ) );
  NOR2_X1 U9602 ( .A1(n2689), .A2(n2811), .ZN(\mult_22/ab[12][51] ) );
  NOR2_X1 U9603 ( .A1(n2672), .A2(n2823), .ZN(\mult_22/ab[14][49] ) );
  NOR2_X1 U9604 ( .A1(n2664), .A2(n2835), .ZN(\mult_22/ab[16][47] ) );
  NOR2_X1 U9605 ( .A1(n2648), .A2(n2847), .ZN(\mult_22/ab[18][45] ) );
  NOR2_X1 U9606 ( .A1(n2636), .A2(n2859), .ZN(\mult_22/ab[20][43] ) );
  NOR2_X1 U9607 ( .A1(n2625), .A2(n2870), .ZN(\mult_22/ab[22][41] ) );
  NOR2_X1 U9608 ( .A1(n2616), .A2(n2882), .ZN(\mult_22/ab[24][39] ) );
  NOR2_X1 U9609 ( .A1(n2545), .A2(n2929), .ZN(\mult_22/ab[32][27] ) );
  NOR2_X1 U9610 ( .A1(n2545), .A2(n2923), .ZN(\mult_22/ab[31][27] ) );
  NOR2_X1 U9611 ( .A1(n2533), .A2(n2941), .ZN(\mult_22/ab[34][25] ) );
  NOR2_X1 U9612 ( .A1(n2533), .A2(n2935), .ZN(\mult_22/ab[33][25] ) );
  NOR2_X1 U9613 ( .A1(n2520), .A2(n2953), .ZN(\mult_22/ab[36][23] ) );
  NOR2_X1 U9614 ( .A1(n2521), .A2(n2947), .ZN(\mult_22/ab[35][23] ) );
  NOR2_X1 U9615 ( .A1(n2508), .A2(n2959), .ZN(\mult_22/ab[37][21] ) );
  NOR2_X1 U9616 ( .A1(n2508), .A2(n2965), .ZN(\mult_22/ab[38][21] ) );
  NOR2_X1 U9617 ( .A1(n2717), .A2(n2758), .ZN(\mult_22/ab[3][57] ) );
  NOR2_X1 U9618 ( .A1(n2550), .A2(n2977), .ZN(\mult_22/ab[40][28] ) );
  NOR2_X1 U9619 ( .A1(n2570), .A2(n2858), .ZN(\mult_22/ab[20][31] ) );
  NOR2_X1 U9620 ( .A1(n2570), .A2(n2864), .ZN(\mult_22/ab[21][31] ) );
  NOR2_X1 U9621 ( .A1(n2570), .A2(n2870), .ZN(\mult_22/ab[22][31] ) );
  NOR2_X1 U9622 ( .A1(n2570), .A2(n2876), .ZN(\mult_22/ab[23][31] ) );
  NOR2_X1 U9623 ( .A1(n2570), .A2(n2882), .ZN(\mult_22/ab[24][31] ) );
  NOR2_X1 U9624 ( .A1(n2570), .A2(n2852), .ZN(\mult_22/ab[19][31] ) );
  NOR2_X1 U9625 ( .A1(n2570), .A2(n2846), .ZN(\mult_22/ab[18][31] ) );
  NOR2_X1 U9626 ( .A1(n2570), .A2(n2840), .ZN(\mult_22/ab[17][31] ) );
  NOR2_X1 U9627 ( .A1(n2570), .A2(n2834), .ZN(\mult_22/ab[16][31] ) );
  NOR2_X1 U9628 ( .A1(n2570), .A2(n2828), .ZN(\mult_22/ab[15][31] ) );
  NOR2_X1 U9629 ( .A1(n2570), .A2(n2822), .ZN(\mult_22/ab[14][31] ) );
  NOR2_X1 U9630 ( .A1(n2704), .A2(n2818), .ZN(\mult_22/ab[13][54] ) );
  NOR2_X1 U9631 ( .A1(n2690), .A2(n2829), .ZN(\mult_22/ab[15][52] ) );
  NOR2_X1 U9632 ( .A1(n2682), .A2(n2841), .ZN(\mult_22/ab[17][50] ) );
  NOR2_X1 U9633 ( .A1(n2670), .A2(n2853), .ZN(\mult_22/ab[19][48] ) );
  NOR2_X1 U9634 ( .A1(n2658), .A2(n2865), .ZN(\mult_22/ab[21][46] ) );
  NOR2_X1 U9635 ( .A1(n2646), .A2(n2877), .ZN(\mult_22/ab[23][44] ) );
  NOR2_X1 U9636 ( .A1(n2634), .A2(n2888), .ZN(\mult_22/ab[25][42] ) );
  NOR2_X1 U9637 ( .A1(n2621), .A2(n2900), .ZN(\mult_22/ab[27][40] ) );
  NOR2_X1 U9638 ( .A1(n2724), .A2(n2794), .ZN(\mult_22/ab[9][58] ) );
  NOR2_X1 U9639 ( .A1(n2556), .A2(n2971), .ZN(\mult_22/ab[39][29] ) );
  NOR2_X1 U9640 ( .A1(n2568), .A2(n2960), .ZN(\mult_22/ab[37][31] ) );
  NOR2_X1 U9641 ( .A1(n2580), .A2(n2948), .ZN(\mult_22/ab[35][33] ) );
  NOR2_X1 U9642 ( .A1(n2592), .A2(n2936), .ZN(\mult_22/ab[33][35] ) );
  NOR2_X1 U9643 ( .A1(n2604), .A2(n2924), .ZN(\mult_22/ab[31][37] ) );
  NOR2_X1 U9644 ( .A1(n2738), .A2(n2776), .ZN(\mult_22/ab[6][61] ) );
  NOR2_X1 U9645 ( .A1(n2735), .A2(n2782), .ZN(\mult_22/ab[7][60] ) );
  NOR2_X1 U9646 ( .A1(n2557), .A2(n2905), .ZN(\mult_22/ab[28][29] ) );
  NOR2_X1 U9647 ( .A1(n2557), .A2(n2899), .ZN(\mult_22/ab[27][29] ) );
  NOR2_X1 U9648 ( .A1(n2603), .A2(n2756), .ZN(\mult_22/ab[3][37] ) );
  NOR2_X1 U9649 ( .A1(n2589), .A2(n2768), .ZN(\mult_22/ab[5][35] ) );
  NOR2_X1 U9650 ( .A1(n2577), .A2(n2780), .ZN(\mult_22/ab[7][33] ) );
  NOR2_X1 U9651 ( .A1(n2562), .A2(n2965), .ZN(\mult_22/ab[38][30] ) );
  NOR2_X1 U9652 ( .A1(n2574), .A2(n2954), .ZN(\mult_22/ab[36][32] ) );
  NOR2_X1 U9653 ( .A1(n2586), .A2(n2942), .ZN(\mult_22/ab[34][34] ) );
  NOR2_X1 U9654 ( .A1(n2598), .A2(n2930), .ZN(\mult_22/ab[32][36] ) );
  NOR2_X1 U9655 ( .A1(n2597), .A2(n2756), .ZN(\mult_22/ab[3][36] ) );
  NOR2_X1 U9656 ( .A1(n2583), .A2(n2768), .ZN(\mult_22/ab[5][34] ) );
  NOR2_X1 U9657 ( .A1(n2727), .A2(n2758), .ZN(\mult_22/ab[3][59] ) );
  NOR2_X1 U9658 ( .A1(n2689), .A2(n2805), .ZN(\mult_22/ab[11][51] ) );
  NOR2_X1 U9659 ( .A1(n2672), .A2(n2817), .ZN(\mult_22/ab[13][49] ) );
  NOR2_X1 U9660 ( .A1(n2610), .A2(n2918), .ZN(\mult_22/ab[30][38] ) );
  NOR2_X1 U9661 ( .A1(n2688), .A2(n2841), .ZN(\mult_22/ab[17][51] ) );
  NOR2_X1 U9662 ( .A1(n2672), .A2(n2853), .ZN(\mult_22/ab[19][49] ) );
  NOR2_X1 U9663 ( .A1(n2664), .A2(n2865), .ZN(\mult_22/ab[21][47] ) );
  NOR2_X1 U9664 ( .A1(n2649), .A2(n2877), .ZN(\mult_22/ab[23][45] ) );
  NOR2_X1 U9665 ( .A1(n2637), .A2(n2889), .ZN(\mult_22/ab[25][43] ) );
  NOR2_X1 U9666 ( .A1(n2625), .A2(n2900), .ZN(\mult_22/ab[27][41] ) );
  NOR2_X1 U9667 ( .A1(n2615), .A2(n2912), .ZN(\mult_22/ab[29][39] ) );
  NOR2_X1 U9668 ( .A1(n2696), .A2(n2830), .ZN(\mult_22/ab[15][53] ) );
  NOR2_X1 U9669 ( .A1(n2711), .A2(n2818), .ZN(\mult_22/ab[13][55] ) );
  NOR2_X1 U9670 ( .A1(n2716), .A2(n2806), .ZN(\mult_22/ab[11][57] ) );
  NOR2_X1 U9671 ( .A1(n2727), .A2(n2794), .ZN(\mult_22/ab[9][59] ) );
  NOR2_X1 U9672 ( .A1(n2722), .A2(n2764), .ZN(\mult_22/ab[4][58] ) );
  NOR2_X1 U9673 ( .A1(n2690), .A2(n2799), .ZN(\mult_22/ab[10][52] ) );
  NOR2_X1 U9674 ( .A1(n2682), .A2(n2811), .ZN(\mult_22/ab[12][50] ) );
  NOR2_X1 U9675 ( .A1(n2670), .A2(n2823), .ZN(\mult_22/ab[14][48] ) );
  NOR2_X1 U9676 ( .A1(n2646), .A2(n2847), .ZN(\mult_22/ab[18][44] ) );
  NOR2_X1 U9677 ( .A1(n2634), .A2(n2859), .ZN(\mult_22/ab[20][42] ) );
  NOR2_X1 U9678 ( .A1(n2622), .A2(n2870), .ZN(\mult_22/ab[22][40] ) );
  NOR2_X1 U9679 ( .A1(n2571), .A2(n2804), .ZN(\mult_22/ab[11][31] ) );
  NOR2_X1 U9680 ( .A1(n2454), .A2(n2976), .ZN(\mult_22/ab[40][12] ) );
  NOR2_X1 U9681 ( .A1(n2690), .A2(n2835), .ZN(\mult_22/ab[16][52] ) );
  NOR2_X1 U9682 ( .A1(n2682), .A2(n2847), .ZN(\mult_22/ab[18][50] ) );
  NOR2_X1 U9683 ( .A1(n2670), .A2(n2859), .ZN(\mult_22/ab[20][48] ) );
  NOR2_X1 U9684 ( .A1(n2658), .A2(n2871), .ZN(\mult_22/ab[22][46] ) );
  NOR2_X1 U9685 ( .A1(n2646), .A2(n2883), .ZN(\mult_22/ab[24][44] ) );
  NOR2_X1 U9686 ( .A1(n2633), .A2(n2895), .ZN(\mult_22/ab[26][42] ) );
  NOR2_X1 U9687 ( .A1(n2621), .A2(n2906), .ZN(\mult_22/ab[28][40] ) );
  NOR2_X1 U9688 ( .A1(n2704), .A2(n2824), .ZN(\mult_22/ab[14][54] ) );
  NOR2_X1 U9689 ( .A1(n2719), .A2(n2800), .ZN(\mult_22/ab[10][58] ) );
  NOR2_X1 U9690 ( .A1(n2616), .A2(n2870), .ZN(\mult_22/ab[22][39] ) );
  NOR2_X1 U9691 ( .A1(n2538), .A2(n2995), .ZN(\mult_22/ab[43][26] ) );
  NOR2_X1 U9692 ( .A1(n2740), .A2(n2782), .ZN(\mult_22/ab[7][61] ) );
  NOR2_X1 U9693 ( .A1(n2591), .A2(n2756), .ZN(\mult_22/ab[3][35] ) );
  NOR2_X1 U9694 ( .A1(n2577), .A2(n2768), .ZN(\mult_22/ab[5][33] ) );
  NOR2_X1 U9695 ( .A1(n2532), .A2(n3001), .ZN(\mult_22/ab[44][25] ) );
  NOR2_X1 U9696 ( .A1(n2544), .A2(n2989), .ZN(\mult_22/ab[42][27] ) );
  NOR2_X1 U9697 ( .A1(n2736), .A2(n2788), .ZN(\mult_22/ab[8][60] ) );
  NOR2_X1 U9698 ( .A1(n2672), .A2(n2811), .ZN(\mult_22/ab[12][49] ) );
  NOR2_X1 U9699 ( .A1(n2648), .A2(n2835), .ZN(\mult_22/ab[16][45] ) );
  NOR2_X1 U9700 ( .A1(n2636), .A2(n2847), .ZN(\mult_22/ab[18][43] ) );
  NOR2_X1 U9701 ( .A1(n2624), .A2(n2858), .ZN(\mult_22/ab[20][41] ) );
  NOR2_X1 U9702 ( .A1(n2684), .A2(n2799), .ZN(\mult_22/ab[10][51] ) );
  NOR2_X1 U9703 ( .A1(n2646), .A2(n2841), .ZN(\mult_22/ab[17][44] ) );
  NOR2_X1 U9704 ( .A1(n2634), .A2(n2853), .ZN(\mult_22/ab[19][42] ) );
  NOR2_X1 U9705 ( .A1(n2622), .A2(n2864), .ZN(\mult_22/ab[21][40] ) );
  NOR2_X1 U9706 ( .A1(n2683), .A2(n2805), .ZN(\mult_22/ab[11][50] ) );
  NOR2_X1 U9707 ( .A1(n2670), .A2(n2817), .ZN(\mult_22/ab[13][48] ) );
  NOR2_X1 U9708 ( .A1(n2658), .A2(n2829), .ZN(\mult_22/ab[15][46] ) );
  NOR2_X1 U9709 ( .A1(n2721), .A2(n2758), .ZN(\mult_22/ab[3][58] ) );
  NOR2_X1 U9710 ( .A1(n2531), .A2(n3025), .ZN(\mult_22/ab[48][25] ) );
  NOR2_X1 U9711 ( .A1(n2585), .A2(n2756), .ZN(\mult_22/ab[3][34] ) );
  NOR2_X1 U9712 ( .A1(n2545), .A2(n2917), .ZN(\mult_22/ab[30][27] ) );
  NOR2_X1 U9713 ( .A1(n2533), .A2(n2929), .ZN(\mult_22/ab[32][25] ) );
  NOR2_X1 U9714 ( .A1(n2521), .A2(n2941), .ZN(\mult_22/ab[34][23] ) );
  NOR2_X1 U9715 ( .A1(n2508), .A2(n2953), .ZN(\mult_22/ab[36][21] ) );
  NOR2_X1 U9716 ( .A1(n2545), .A2(n2911), .ZN(\mult_22/ab[29][27] ) );
  NOR2_X1 U9717 ( .A1(n2533), .A2(n2923), .ZN(\mult_22/ab[31][25] ) );
  NOR2_X1 U9718 ( .A1(n2521), .A2(n2935), .ZN(\mult_22/ab[33][23] ) );
  NOR2_X1 U9719 ( .A1(n2509), .A2(n2947), .ZN(\mult_22/ab[35][21] ) );
  NOR2_X1 U9720 ( .A1(n2496), .A2(n2958), .ZN(\mult_22/ab[37][19] ) );
  NOR2_X1 U9721 ( .A1(n2558), .A2(n2875), .ZN(\mult_22/ab[23][29] ) );
  NOR2_X1 U9722 ( .A1(n2558), .A2(n2881), .ZN(\mult_22/ab[24][29] ) );
  NOR2_X1 U9723 ( .A1(n2557), .A2(n2887), .ZN(\mult_22/ab[25][29] ) );
  NOR2_X1 U9724 ( .A1(n2557), .A2(n2893), .ZN(\mult_22/ab[26][29] ) );
  NOR2_X1 U9725 ( .A1(n2558), .A2(n2869), .ZN(\mult_22/ab[22][29] ) );
  NOR2_X1 U9726 ( .A1(n2558), .A2(n2863), .ZN(\mult_22/ab[21][29] ) );
  NOR2_X1 U9727 ( .A1(n2558), .A2(n2857), .ZN(\mult_22/ab[20][29] ) );
  NOR2_X1 U9728 ( .A1(n2558), .A2(n2851), .ZN(\mult_22/ab[19][29] ) );
  NOR2_X1 U9729 ( .A1(n2717), .A2(n2764), .ZN(\mult_22/ab[4][57] ) );
  NOR2_X1 U9730 ( .A1(n2558), .A2(n2845), .ZN(\mult_22/ab[18][29] ) );
  NOR2_X1 U9731 ( .A1(n2558), .A2(n2839), .ZN(\mult_22/ab[17][29] ) );
  NOR2_X1 U9732 ( .A1(n2558), .A2(n2833), .ZN(\mult_22/ab[16][29] ) );
  NOR2_X1 U9733 ( .A1(n2407), .A2(n3033), .ZN(\mult_22/ab[49][4] ) );
  NOR2_X1 U9734 ( .A1(n2558), .A2(n2827), .ZN(\mult_22/ab[15][29] ) );
  NOR2_X1 U9735 ( .A1(n2558), .A2(n2821), .ZN(\mult_22/ab[14][29] ) );
  NOR2_X1 U9736 ( .A1(n2550), .A2(n2983), .ZN(\mult_22/ab[41][28] ) );
  NOR2_X1 U9737 ( .A1(n2566), .A2(n2792), .ZN(\mult_22/ab[9][31] ) );
  NOR2_X1 U9738 ( .A1(n2579), .A2(n2756), .ZN(\mult_22/ab[3][33] ) );
  NOR2_X1 U9739 ( .A1(n2562), .A2(n2971), .ZN(\mult_22/ab[39][30] ) );
  NOR2_X1 U9740 ( .A1(n2574), .A2(n2960), .ZN(\mult_22/ab[37][32] ) );
  NOR2_X1 U9741 ( .A1(n2556), .A2(n2977), .ZN(\mult_22/ab[40][29] ) );
  NOR2_X1 U9742 ( .A1(n2586), .A2(n2948), .ZN(\mult_22/ab[35][34] ) );
  NOR2_X1 U9743 ( .A1(n2568), .A2(n2966), .ZN(\mult_22/ab[38][31] ) );
  NOR2_X1 U9744 ( .A1(n2580), .A2(n2954), .ZN(\mult_22/ab[36][33] ) );
  NOR2_X1 U9745 ( .A1(n2592), .A2(n2942), .ZN(\mult_22/ab[34][35] ) );
  NOR2_X1 U9746 ( .A1(n2604), .A2(n2930), .ZN(\mult_22/ab[32][37] ) );
  NOR2_X1 U9747 ( .A1(n2598), .A2(n2936), .ZN(\mult_22/ab[33][36] ) );
  NOR2_X1 U9748 ( .A1(n2532), .A2(n3007), .ZN(\mult_22/ab[45][25] ) );
  NOR2_X1 U9749 ( .A1(n2558), .A2(n2815), .ZN(\mult_22/ab[13][29] ) );
  NOR2_X1 U9750 ( .A1(n2544), .A2(n2995), .ZN(\mult_22/ab[43][27] ) );
  NOR2_X1 U9751 ( .A1(n2610), .A2(n2924), .ZN(\mult_22/ab[31][38] ) );
  NOR2_X1 U9752 ( .A1(n2538), .A2(n3001), .ZN(\mult_22/ab[44][26] ) );
  NOR2_X1 U9753 ( .A1(n2566), .A2(n2780), .ZN(\mult_22/ab[7][31] ) );
  NOR2_X1 U9754 ( .A1(n2672), .A2(n2859), .ZN(\mult_22/ab[20][49] ) );
  NOR2_X1 U9755 ( .A1(n2664), .A2(n2871), .ZN(\mult_22/ab[22][47] ) );
  NOR2_X1 U9756 ( .A1(n2649), .A2(n2883), .ZN(\mult_22/ab[24][45] ) );
  NOR2_X1 U9757 ( .A1(n2637), .A2(n2895), .ZN(\mult_22/ab[26][43] ) );
  NOR2_X1 U9758 ( .A1(n2625), .A2(n2906), .ZN(\mult_22/ab[28][41] ) );
  NOR2_X1 U9759 ( .A1(n2615), .A2(n2918), .ZN(\mult_22/ab[30][39] ) );
  NOR2_X1 U9760 ( .A1(n2688), .A2(n2847), .ZN(\mult_22/ab[18][51] ) );
  NOR2_X1 U9761 ( .A1(n2697), .A2(n2836), .ZN(\mult_22/ab[16][53] ) );
  NOR2_X1 U9762 ( .A1(n2710), .A2(n2824), .ZN(\mult_22/ab[14][55] ) );
  NOR2_X1 U9763 ( .A1(n2716), .A2(n2812), .ZN(\mult_22/ab[12][57] ) );
  NOR2_X1 U9764 ( .A1(n2728), .A2(n2800), .ZN(\mult_22/ab[10][59] ) );
  NOR2_X1 U9765 ( .A1(n2531), .A2(n3019), .ZN(\mult_22/ab[47][25] ) );
  NOR2_X1 U9766 ( .A1(n2682), .A2(n2853), .ZN(\mult_22/ab[19][50] ) );
  NOR2_X1 U9767 ( .A1(n2670), .A2(n2865), .ZN(\mult_22/ab[21][48] ) );
  NOR2_X1 U9768 ( .A1(n2658), .A2(n2877), .ZN(\mult_22/ab[23][46] ) );
  NOR2_X1 U9769 ( .A1(n2646), .A2(n2889), .ZN(\mult_22/ab[25][44] ) );
  NOR2_X1 U9770 ( .A1(n2633), .A2(n2901), .ZN(\mult_22/ab[27][42] ) );
  NOR2_X1 U9771 ( .A1(n2621), .A2(n2912), .ZN(\mult_22/ab[29][40] ) );
  NOR2_X1 U9772 ( .A1(n2690), .A2(n2841), .ZN(\mult_22/ab[17][52] ) );
  NOR2_X1 U9773 ( .A1(n2704), .A2(n2830), .ZN(\mult_22/ab[15][54] ) );
  NOR2_X1 U9774 ( .A1(n2719), .A2(n2806), .ZN(\mult_22/ab[11][58] ) );
  NOR2_X1 U9775 ( .A1(n2418), .A2(n3017), .ZN(\mult_22/ab[46][6] ) );
  NOR2_X1 U9776 ( .A1(n2559), .A2(n2809), .ZN(\mult_22/ab[12][29] ) );
  NOR2_X1 U9777 ( .A1(n2538), .A2(n3007), .ZN(\mult_22/ab[45][26] ) );
  NOR2_X1 U9778 ( .A1(n2545), .A2(n2887), .ZN(\mult_22/ab[25][27] ) );
  NOR2_X1 U9779 ( .A1(n2545), .A2(n2893), .ZN(\mult_22/ab[26][27] ) );
  NOR2_X1 U9780 ( .A1(n2533), .A2(n2905), .ZN(\mult_22/ab[28][25] ) );
  NOR2_X1 U9781 ( .A1(n2533), .A2(n2911), .ZN(\mult_22/ab[29][25] ) );
  NOR2_X1 U9782 ( .A1(n2521), .A2(n2923), .ZN(\mult_22/ab[31][23] ) );
  NOR2_X1 U9783 ( .A1(n2521), .A2(n2929), .ZN(\mult_22/ab[32][23] ) );
  NOR2_X1 U9784 ( .A1(n2509), .A2(n2941), .ZN(\mult_22/ab[34][21] ) );
  NOR2_X1 U9785 ( .A1(n2546), .A2(n2881), .ZN(\mult_22/ab[24][27] ) );
  NOR2_X1 U9786 ( .A1(n2533), .A2(n2899), .ZN(\mult_22/ab[27][25] ) );
  NOR2_X1 U9787 ( .A1(n2545), .A2(n2899), .ZN(\mult_22/ab[27][27] ) );
  NOR2_X1 U9788 ( .A1(n2521), .A2(n2917), .ZN(\mult_22/ab[30][23] ) );
  NOR2_X1 U9789 ( .A1(n2533), .A2(n2917), .ZN(\mult_22/ab[30][25] ) );
  NOR2_X1 U9790 ( .A1(n2509), .A2(n2935), .ZN(\mult_22/ab[33][21] ) );
  NOR2_X1 U9791 ( .A1(n2496), .A2(n2952), .ZN(\mult_22/ab[36][19] ) );
  NOR2_X1 U9792 ( .A1(n2546), .A2(n2875), .ZN(\mult_22/ab[23][27] ) );
  NOR2_X1 U9793 ( .A1(n2533), .A2(n2893), .ZN(\mult_22/ab[26][25] ) );
  NOR2_X1 U9794 ( .A1(n2545), .A2(n2905), .ZN(\mult_22/ab[28][27] ) );
  NOR2_X1 U9795 ( .A1(n2521), .A2(n2911), .ZN(\mult_22/ab[29][23] ) );
  NOR2_X1 U9796 ( .A1(n2509), .A2(n2929), .ZN(\mult_22/ab[32][21] ) );
  NOR2_X1 U9797 ( .A1(n2497), .A2(n2946), .ZN(\mult_22/ab[35][19] ) );
  NOR2_X1 U9798 ( .A1(n2546), .A2(n2869), .ZN(\mult_22/ab[22][27] ) );
  NOR2_X1 U9799 ( .A1(n2533), .A2(n2887), .ZN(\mult_22/ab[25][25] ) );
  NOR2_X1 U9800 ( .A1(n2521), .A2(n2905), .ZN(\mult_22/ab[28][23] ) );
  NOR2_X1 U9801 ( .A1(n2509), .A2(n2923), .ZN(\mult_22/ab[31][21] ) );
  NOR2_X1 U9802 ( .A1(n2497), .A2(n2940), .ZN(\mult_22/ab[34][19] ) );
  NOR2_X1 U9803 ( .A1(n2484), .A2(n2958), .ZN(\mult_22/ab[37][17] ) );
  NOR2_X1 U9804 ( .A1(n2546), .A2(n2863), .ZN(\mult_22/ab[21][27] ) );
  NOR2_X1 U9805 ( .A1(n2534), .A2(n2881), .ZN(\mult_22/ab[24][25] ) );
  NOR2_X1 U9806 ( .A1(n2521), .A2(n2899), .ZN(\mult_22/ab[27][23] ) );
  NOR2_X1 U9807 ( .A1(n2509), .A2(n2917), .ZN(\mult_22/ab[30][21] ) );
  NOR2_X1 U9808 ( .A1(n2497), .A2(n2934), .ZN(\mult_22/ab[33][19] ) );
  NOR2_X1 U9809 ( .A1(n2484), .A2(n2952), .ZN(\mult_22/ab[36][17] ) );
  NOR2_X1 U9810 ( .A1(n2546), .A2(n2857), .ZN(\mult_22/ab[20][27] ) );
  NOR2_X1 U9811 ( .A1(n2534), .A2(n2875), .ZN(\mult_22/ab[23][25] ) );
  NOR2_X1 U9812 ( .A1(n2521), .A2(n2893), .ZN(\mult_22/ab[26][23] ) );
  NOR2_X1 U9813 ( .A1(n2509), .A2(n2911), .ZN(\mult_22/ab[29][21] ) );
  NOR2_X1 U9814 ( .A1(n2497), .A2(n2928), .ZN(\mult_22/ab[32][19] ) );
  NOR2_X1 U9815 ( .A1(n2485), .A2(n2946), .ZN(\mult_22/ab[35][17] ) );
  NOR2_X1 U9816 ( .A1(n2546), .A2(n2851), .ZN(\mult_22/ab[19][27] ) );
  NOR2_X1 U9817 ( .A1(n2534), .A2(n2869), .ZN(\mult_22/ab[22][25] ) );
  NOR2_X1 U9818 ( .A1(n2521), .A2(n2887), .ZN(\mult_22/ab[25][23] ) );
  NOR2_X1 U9819 ( .A1(n2509), .A2(n2905), .ZN(\mult_22/ab[28][21] ) );
  NOR2_X1 U9820 ( .A1(n2497), .A2(n2922), .ZN(\mult_22/ab[31][19] ) );
  NOR2_X1 U9821 ( .A1(n2485), .A2(n2940), .ZN(\mult_22/ab[34][17] ) );
  NOR2_X1 U9822 ( .A1(n2546), .A2(n2845), .ZN(\mult_22/ab[18][27] ) );
  NOR2_X1 U9823 ( .A1(n2534), .A2(n2863), .ZN(\mult_22/ab[21][25] ) );
  NOR2_X1 U9824 ( .A1(n2522), .A2(n2881), .ZN(\mult_22/ab[24][23] ) );
  NOR2_X1 U9825 ( .A1(n2509), .A2(n2899), .ZN(\mult_22/ab[27][21] ) );
  NOR2_X1 U9826 ( .A1(n2497), .A2(n2916), .ZN(\mult_22/ab[30][19] ) );
  NOR2_X1 U9827 ( .A1(n2485), .A2(n2934), .ZN(\mult_22/ab[33][17] ) );
  NOR2_X1 U9828 ( .A1(n2534), .A2(n2857), .ZN(\mult_22/ab[20][25] ) );
  NOR2_X1 U9829 ( .A1(n2522), .A2(n2875), .ZN(\mult_22/ab[23][23] ) );
  NOR2_X1 U9830 ( .A1(n2509), .A2(n2893), .ZN(\mult_22/ab[26][21] ) );
  NOR2_X1 U9831 ( .A1(n2497), .A2(n2910), .ZN(\mult_22/ab[29][19] ) );
  NOR2_X1 U9832 ( .A1(n2485), .A2(n2928), .ZN(\mult_22/ab[32][17] ) );
  NOR2_X1 U9833 ( .A1(n2472), .A2(n2964), .ZN(\mult_22/ab[38][15] ) );
  NOR2_X1 U9834 ( .A1(n2522), .A2(n2869), .ZN(\mult_22/ab[22][23] ) );
  NOR2_X1 U9835 ( .A1(n2509), .A2(n2887), .ZN(\mult_22/ab[25][21] ) );
  NOR2_X1 U9836 ( .A1(n2497), .A2(n2904), .ZN(\mult_22/ab[28][19] ) );
  NOR2_X1 U9837 ( .A1(n2485), .A2(n2922), .ZN(\mult_22/ab[31][17] ) );
  NOR2_X1 U9838 ( .A1(n2472), .A2(n2958), .ZN(\mult_22/ab[37][15] ) );
  NOR2_X1 U9839 ( .A1(n2510), .A2(n2881), .ZN(\mult_22/ab[24][21] ) );
  NOR2_X1 U9840 ( .A1(n2497), .A2(n2898), .ZN(\mult_22/ab[27][19] ) );
  NOR2_X1 U9841 ( .A1(n2485), .A2(n2916), .ZN(\mult_22/ab[30][17] ) );
  NOR2_X1 U9842 ( .A1(n2472), .A2(n2952), .ZN(\mult_22/ab[36][15] ) );
  NOR2_X1 U9843 ( .A1(n2497), .A2(n2892), .ZN(\mult_22/ab[26][19] ) );
  NOR2_X1 U9844 ( .A1(n2485), .A2(n2910), .ZN(\mult_22/ab[29][17] ) );
  NOR2_X1 U9845 ( .A1(n2473), .A2(n2946), .ZN(\mult_22/ab[35][15] ) );
  NOR2_X1 U9846 ( .A1(n2485), .A2(n2904), .ZN(\mult_22/ab[28][17] ) );
  NOR2_X1 U9847 ( .A1(n2473), .A2(n2940), .ZN(\mult_22/ab[34][15] ) );
  NOR2_X1 U9848 ( .A1(n2473), .A2(n2934), .ZN(\mult_22/ab[33][15] ) );
  NOR2_X1 U9849 ( .A1(n2473), .A2(n2928), .ZN(\mult_22/ab[32][15] ) );
  NOR2_X1 U9850 ( .A1(n2473), .A2(n2922), .ZN(\mult_22/ab[31][15] ) );
  NOR2_X1 U9851 ( .A1(n2473), .A2(n2916), .ZN(\mult_22/ab[30][15] ) );
  NOR2_X1 U9852 ( .A1(n2736), .A2(n2794), .ZN(\mult_22/ab[9][60] ) );
  NOR2_X1 U9853 ( .A1(n2454), .A2(n2970), .ZN(\mult_22/ab[39][12] ) );
  NOR2_X1 U9854 ( .A1(n2454), .A2(n2964), .ZN(\mult_22/ab[38][12] ) );
  NOR2_X1 U9855 ( .A1(n2442), .A2(n2982), .ZN(\mult_22/ab[41][10] ) );
  NOR2_X1 U9856 ( .A1(n2454), .A2(n2958), .ZN(\mult_22/ab[37][12] ) );
  NOR2_X1 U9857 ( .A1(n2442), .A2(n2976), .ZN(\mult_22/ab[40][10] ) );
  NOR2_X1 U9858 ( .A1(n2430), .A2(n2999), .ZN(\mult_22/ab[43][8] ) );
  NOR2_X1 U9859 ( .A1(n2454), .A2(n2952), .ZN(\mult_22/ab[36][12] ) );
  NOR2_X1 U9860 ( .A1(n2442), .A2(n2970), .ZN(\mult_22/ab[39][10] ) );
  NOR2_X1 U9861 ( .A1(n2430), .A2(n2993), .ZN(\mult_22/ab[42][8] ) );
  NOR2_X1 U9862 ( .A1(n2418), .A2(n3011), .ZN(\mult_22/ab[45][6] ) );
  NOR2_X1 U9863 ( .A1(n2407), .A2(n3027), .ZN(\mult_22/ab[48][4] ) );
  NOR2_X1 U9864 ( .A1(n2455), .A2(n2946), .ZN(\mult_22/ab[35][12] ) );
  NOR2_X1 U9865 ( .A1(n2442), .A2(n2964), .ZN(\mult_22/ab[38][10] ) );
  NOR2_X1 U9866 ( .A1(n2430), .A2(n2987), .ZN(\mult_22/ab[41][8] ) );
  NOR2_X1 U9867 ( .A1(n2418), .A2(n3005), .ZN(\mult_22/ab[44][6] ) );
  NOR2_X1 U9868 ( .A1(n2407), .A2(n3021), .ZN(\mult_22/ab[47][4] ) );
  NOR2_X1 U9869 ( .A1(n2455), .A2(n2940), .ZN(\mult_22/ab[34][12] ) );
  NOR2_X1 U9870 ( .A1(n2442), .A2(n2958), .ZN(\mult_22/ab[37][10] ) );
  NOR2_X1 U9871 ( .A1(n2430), .A2(n2981), .ZN(\mult_22/ab[40][8] ) );
  NOR2_X1 U9872 ( .A1(n2418), .A2(n2999), .ZN(\mult_22/ab[43][6] ) );
  NOR2_X1 U9873 ( .A1(n2407), .A2(n3015), .ZN(\mult_22/ab[46][4] ) );
  NOR2_X1 U9874 ( .A1(n2455), .A2(n2934), .ZN(\mult_22/ab[33][12] ) );
  NOR2_X1 U9875 ( .A1(n2442), .A2(n2952), .ZN(\mult_22/ab[36][10] ) );
  NOR2_X1 U9876 ( .A1(n2430), .A2(n2975), .ZN(\mult_22/ab[39][8] ) );
  NOR2_X1 U9877 ( .A1(n2418), .A2(n2993), .ZN(\mult_22/ab[42][6] ) );
  NOR2_X1 U9878 ( .A1(n2407), .A2(n3009), .ZN(\mult_22/ab[45][4] ) );
  NOR2_X1 U9879 ( .A1(n2442), .A2(n2946), .ZN(\mult_22/ab[35][10] ) );
  NOR2_X1 U9880 ( .A1(n2430), .A2(n2969), .ZN(\mult_22/ab[38][8] ) );
  NOR2_X1 U9881 ( .A1(n2418), .A2(n2987), .ZN(\mult_22/ab[41][6] ) );
  NOR2_X1 U9882 ( .A1(n2407), .A2(n3003), .ZN(\mult_22/ab[44][4] ) );
  NOR2_X1 U9883 ( .A1(n2430), .A2(n2963), .ZN(\mult_22/ab[37][8] ) );
  NOR2_X1 U9884 ( .A1(n2418), .A2(n2981), .ZN(\mult_22/ab[40][6] ) );
  NOR2_X1 U9885 ( .A1(n2406), .A2(n2997), .ZN(\mult_22/ab[43][4] ) );
  NOR2_X1 U9886 ( .A1(n2418), .A2(n2975), .ZN(\mult_22/ab[39][6] ) );
  NOR2_X1 U9887 ( .A1(n2406), .A2(n2991), .ZN(\mult_22/ab[42][4] ) );
  NOR2_X1 U9888 ( .A1(n2406), .A2(n2985), .ZN(\mult_22/ab[41][4] ) );
  NOR2_X1 U9889 ( .A1(n2540), .A2(n2845), .ZN(\mult_22/ab[18][26] ) );
  NOR2_X1 U9890 ( .A1(n2540), .A2(n2839), .ZN(\mult_22/ab[17][26] ) );
  NOR2_X1 U9891 ( .A1(n2524), .A2(n2857), .ZN(\mult_22/ab[20][24] ) );
  NOR2_X1 U9892 ( .A1(n2524), .A2(n2851), .ZN(\mult_22/ab[19][24] ) );
  NOR2_X1 U9893 ( .A1(n2516), .A2(n2869), .ZN(\mult_22/ab[22][22] ) );
  NOR2_X1 U9894 ( .A1(n2516), .A2(n2863), .ZN(\mult_22/ab[21][22] ) );
  NOR2_X1 U9895 ( .A1(n2504), .A2(n2881), .ZN(\mult_22/ab[24][20] ) );
  NOR2_X1 U9896 ( .A1(n2504), .A2(n2875), .ZN(\mult_22/ab[23][20] ) );
  NOR2_X1 U9897 ( .A1(n2491), .A2(n2892), .ZN(\mult_22/ab[26][18] ) );
  NOR2_X1 U9898 ( .A1(n2491), .A2(n2886), .ZN(\mult_22/ab[25][18] ) );
  NOR2_X1 U9899 ( .A1(n2479), .A2(n2904), .ZN(\mult_22/ab[28][16] ) );
  NOR2_X1 U9900 ( .A1(n2479), .A2(n2898), .ZN(\mult_22/ab[27][16] ) );
  NOR2_X1 U9901 ( .A1(n2741), .A2(n2788), .ZN(\mult_22/ab[8][61] ) );
  NOR2_X1 U9902 ( .A1(n2467), .A2(n2916), .ZN(\mult_22/ab[30][14] ) );
  NOR2_X1 U9903 ( .A1(n2467), .A2(n2910), .ZN(\mult_22/ab[29][14] ) );
  NOR2_X1 U9904 ( .A1(n2532), .A2(n3013), .ZN(\mult_22/ab[46][25] ) );
  NOR2_X1 U9905 ( .A1(n2544), .A2(n3001), .ZN(\mult_22/ab[44][27] ) );
  NOR2_X1 U9906 ( .A1(n2550), .A2(n2989), .ZN(\mult_22/ab[42][28] ) );
  NOR2_X1 U9907 ( .A1(n2455), .A2(n2928), .ZN(\mult_22/ab[32][12] ) );
  NOR2_X1 U9908 ( .A1(n2455), .A2(n2922), .ZN(\mult_22/ab[31][12] ) );
  NOR2_X1 U9909 ( .A1(n2442), .A2(n2940), .ZN(\mult_22/ab[34][10] ) );
  NOR2_X1 U9910 ( .A1(n2442), .A2(n2934), .ZN(\mult_22/ab[33][10] ) );
  NOR2_X1 U9911 ( .A1(n2430), .A2(n2957), .ZN(\mult_22/ab[36][8] ) );
  NOR2_X1 U9912 ( .A1(n2431), .A2(n2951), .ZN(\mult_22/ab[35][8] ) );
  NOR2_X1 U9913 ( .A1(n2418), .A2(n2969), .ZN(\mult_22/ab[38][6] ) );
  NOR2_X1 U9914 ( .A1(n2418), .A2(n2963), .ZN(\mult_22/ab[37][6] ) );
  NOR2_X1 U9915 ( .A1(n2406), .A2(n2979), .ZN(\mult_22/ab[40][4] ) );
  NOR2_X1 U9916 ( .A1(n2406), .A2(n2973), .ZN(\mult_22/ab[39][4] ) );
  NOR2_X1 U9917 ( .A1(n2559), .A2(n2803), .ZN(\mult_22/ab[11][29] ) );
  NOR2_X1 U9918 ( .A1(n2556), .A2(n2983), .ZN(\mult_22/ab[41][29] ) );
  NOR2_X1 U9919 ( .A1(n2568), .A2(n2972), .ZN(\mult_22/ab[39][31] ) );
  NOR2_X1 U9920 ( .A1(n2579), .A2(n2960), .ZN(\mult_22/ab[37][33] ) );
  NOR2_X1 U9921 ( .A1(n2592), .A2(n2948), .ZN(\mult_22/ab[35][35] ) );
  NOR2_X1 U9922 ( .A1(n2604), .A2(n2936), .ZN(\mult_22/ab[33][37] ) );
  NOR2_X1 U9923 ( .A1(n2566), .A2(n2768), .ZN(\mult_22/ab[5][31] ) );
  NOR2_X1 U9924 ( .A1(n2559), .A2(n2797), .ZN(\mult_22/ab[10][29] ) );
  NOR2_X1 U9925 ( .A1(n2562), .A2(n2977), .ZN(\mult_22/ab[40][30] ) );
  NOR2_X1 U9926 ( .A1(n2574), .A2(n2966), .ZN(\mult_22/ab[38][32] ) );
  NOR2_X1 U9927 ( .A1(n2585), .A2(n2954), .ZN(\mult_22/ab[36][34] ) );
  NOR2_X1 U9928 ( .A1(n2598), .A2(n2942), .ZN(\mult_22/ab[34][36] ) );
  NOR2_X1 U9929 ( .A1(n2550), .A2(n2995), .ZN(\mult_22/ab[43][28] ) );
  NOR2_X1 U9930 ( .A1(n2546), .A2(n2827), .ZN(\mult_22/ab[15][27] ) );
  NOR2_X1 U9931 ( .A1(n2534), .A2(n2839), .ZN(\mult_22/ab[17][25] ) );
  NOR2_X1 U9932 ( .A1(n2522), .A2(n2851), .ZN(\mult_22/ab[19][23] ) );
  NOR2_X1 U9933 ( .A1(n2510), .A2(n2863), .ZN(\mult_22/ab[21][21] ) );
  NOR2_X1 U9934 ( .A1(n2498), .A2(n2874), .ZN(\mult_22/ab[23][19] ) );
  NOR2_X1 U9935 ( .A1(n2485), .A2(n2886), .ZN(\mult_22/ab[25][17] ) );
  NOR2_X1 U9936 ( .A1(n2473), .A2(n2898), .ZN(\mult_22/ab[27][15] ) );
  NOR2_X1 U9937 ( .A1(n2610), .A2(n2930), .ZN(\mult_22/ab[32][38] ) );
  NOR2_X1 U9938 ( .A1(n2461), .A2(n2910), .ZN(\mult_22/ab[29][13] ) );
  NOR2_X1 U9939 ( .A1(n2449), .A2(n2922), .ZN(\mult_22/ab[31][11] ) );
  NOR2_X1 U9940 ( .A1(n2437), .A2(n2939), .ZN(\mult_22/ab[33][9] ) );
  NOR2_X1 U9941 ( .A1(n2425), .A2(n2951), .ZN(\mult_22/ab[35][7] ) );
  NOR2_X1 U9942 ( .A1(n2412), .A2(n2962), .ZN(\mult_22/ab[37][5] ) );
  NOR2_X1 U9943 ( .A1(n2664), .A2(n2877), .ZN(\mult_22/ab[23][47] ) );
  NOR2_X1 U9944 ( .A1(n2649), .A2(n2889), .ZN(\mult_22/ab[25][45] ) );
  NOR2_X1 U9945 ( .A1(n2637), .A2(n2901), .ZN(\mult_22/ab[27][43] ) );
  NOR2_X1 U9946 ( .A1(n2625), .A2(n2912), .ZN(\mult_22/ab[29][41] ) );
  NOR2_X1 U9947 ( .A1(n2615), .A2(n2924), .ZN(\mult_22/ab[31][39] ) );
  NOR2_X1 U9948 ( .A1(n2672), .A2(n2865), .ZN(\mult_22/ab[21][49] ) );
  NOR2_X1 U9949 ( .A1(n2688), .A2(n2853), .ZN(\mult_22/ab[19][51] ) );
  NOR2_X1 U9950 ( .A1(n2700), .A2(n2842), .ZN(\mult_22/ab[17][53] ) );
  NOR2_X1 U9951 ( .A1(n2710), .A2(n2830), .ZN(\mult_22/ab[15][55] ) );
  NOR2_X1 U9952 ( .A1(n2716), .A2(n2818), .ZN(\mult_22/ab[13][57] ) );
  NOR2_X1 U9953 ( .A1(n2729), .A2(n2806), .ZN(\mult_22/ab[11][59] ) );
  NOR2_X1 U9954 ( .A1(n2562), .A2(n2983), .ZN(\mult_22/ab[41][30] ) );
  NOR2_X1 U9955 ( .A1(n2574), .A2(n2972), .ZN(\mult_22/ab[39][32] ) );
  NOR2_X1 U9956 ( .A1(n2585), .A2(n2960), .ZN(\mult_22/ab[37][34] ) );
  NOR2_X1 U9957 ( .A1(n2598), .A2(n2948), .ZN(\mult_22/ab[35][36] ) );
  NOR2_X1 U9958 ( .A1(n2556), .A2(n2989), .ZN(\mult_22/ab[42][29] ) );
  NOR2_X1 U9959 ( .A1(n2568), .A2(n2978), .ZN(\mult_22/ab[40][31] ) );
  NOR2_X1 U9960 ( .A1(n2579), .A2(n2966), .ZN(\mult_22/ab[38][33] ) );
  NOR2_X1 U9961 ( .A1(n2591), .A2(n2954), .ZN(\mult_22/ab[36][35] ) );
  NOR2_X1 U9962 ( .A1(n2604), .A2(n2942), .ZN(\mult_22/ab[34][37] ) );
  NOR2_X1 U9963 ( .A1(n2538), .A2(n3013), .ZN(\mult_22/ab[46][26] ) );
  NOR2_X1 U9964 ( .A1(n2540), .A2(n2827), .ZN(\mult_22/ab[15][26] ) );
  NOR2_X1 U9965 ( .A1(n2524), .A2(n2839), .ZN(\mult_22/ab[17][24] ) );
  NOR2_X1 U9966 ( .A1(n2516), .A2(n2851), .ZN(\mult_22/ab[19][22] ) );
  NOR2_X1 U9967 ( .A1(n2504), .A2(n2863), .ZN(\mult_22/ab[21][20] ) );
  NOR2_X1 U9968 ( .A1(n2492), .A2(n2874), .ZN(\mult_22/ab[23][18] ) );
  NOR2_X1 U9969 ( .A1(n2479), .A2(n2886), .ZN(\mult_22/ab[25][16] ) );
  NOR2_X1 U9970 ( .A1(n2554), .A2(n2791), .ZN(\mult_22/ab[9][29] ) );
  NOR2_X1 U9971 ( .A1(n2467), .A2(n2898), .ZN(\mult_22/ab[27][14] ) );
  NOR2_X1 U9972 ( .A1(n2544), .A2(n3007), .ZN(\mult_22/ab[45][27] ) );
  NOR2_X1 U9973 ( .A1(n2455), .A2(n2910), .ZN(\mult_22/ab[29][12] ) );
  NOR2_X1 U9974 ( .A1(n2441), .A2(n2922), .ZN(\mult_22/ab[31][10] ) );
  NOR2_X1 U9975 ( .A1(n2431), .A2(n2939), .ZN(\mult_22/ab[33][8] ) );
  NOR2_X1 U9976 ( .A1(n2419), .A2(n2951), .ZN(\mult_22/ab[35][6] ) );
  NOR2_X1 U9977 ( .A1(n2406), .A2(n2961), .ZN(\mult_22/ab[37][4] ) );
  NOR2_X1 U9978 ( .A1(n2670), .A2(n2871), .ZN(\mult_22/ab[22][48] ) );
  NOR2_X1 U9979 ( .A1(n2658), .A2(n2883), .ZN(\mult_22/ab[24][46] ) );
  NOR2_X1 U9980 ( .A1(n2645), .A2(n2895), .ZN(\mult_22/ab[26][44] ) );
  NOR2_X1 U9981 ( .A1(n2633), .A2(n2906), .ZN(\mult_22/ab[28][42] ) );
  NOR2_X1 U9982 ( .A1(n2621), .A2(n2918), .ZN(\mult_22/ab[30][40] ) );
  NOR2_X1 U9983 ( .A1(n2682), .A2(n2859), .ZN(\mult_22/ab[20][50] ) );
  NOR2_X1 U9984 ( .A1(n2690), .A2(n2847), .ZN(\mult_22/ab[18][52] ) );
  NOR2_X1 U9985 ( .A1(n2704), .A2(n2836), .ZN(\mult_22/ab[16][54] ) );
  NOR2_X1 U9986 ( .A1(n2719), .A2(n2812), .ZN(\mult_22/ab[12][58] ) );
  NOR2_X1 U9987 ( .A1(n2610), .A2(n2936), .ZN(\mult_22/ab[33][38] ) );
  NOR2_X1 U9988 ( .A1(n2737), .A2(n2794), .ZN(\mult_22/ab[9][61] ) );
  NOR2_X1 U9989 ( .A1(n2731), .A2(n2800), .ZN(\mult_22/ab[10][60] ) );
  NOR2_X1 U9990 ( .A1(n2554), .A2(n2785), .ZN(\mult_22/ab[8][29] ) );
  NOR2_X1 U9991 ( .A1(n2649), .A2(n2895), .ZN(\mult_22/ab[26][45] ) );
  NOR2_X1 U9992 ( .A1(n2637), .A2(n2907), .ZN(\mult_22/ab[28][43] ) );
  NOR2_X1 U9993 ( .A1(n2625), .A2(n2918), .ZN(\mult_22/ab[30][41] ) );
  NOR2_X1 U9994 ( .A1(n2615), .A2(n2930), .ZN(\mult_22/ab[32][39] ) );
  NOR2_X1 U9995 ( .A1(n2664), .A2(n2883), .ZN(\mult_22/ab[24][47] ) );
  NOR2_X1 U9996 ( .A1(n2673), .A2(n2871), .ZN(\mult_22/ab[22][49] ) );
  NOR2_X1 U9997 ( .A1(n2688), .A2(n2859), .ZN(\mult_22/ab[20][51] ) );
  NOR2_X1 U9998 ( .A1(n2568), .A2(n2756), .ZN(\mult_22/ab[3][31] ) );
  NOR2_X1 U9999 ( .A1(n2695), .A2(n2847), .ZN(\mult_22/ab[18][53] ) );
  NOR2_X1 U10000 ( .A1(n2710), .A2(n2836), .ZN(\mult_22/ab[16][55] ) );
  NOR2_X1 U10001 ( .A1(n2716), .A2(n2824), .ZN(\mult_22/ab[14][57] ) );
  NOR2_X1 U10002 ( .A1(n2730), .A2(n2812), .ZN(\mult_22/ab[12][59] ) );
  NOR2_X1 U10003 ( .A1(n2657), .A2(n2889), .ZN(\mult_22/ab[25][46] ) );
  NOR2_X1 U10004 ( .A1(n2645), .A2(n2901), .ZN(\mult_22/ab[27][44] ) );
  NOR2_X1 U10005 ( .A1(n2633), .A2(n2913), .ZN(\mult_22/ab[29][42] ) );
  NOR2_X1 U10006 ( .A1(n2621), .A2(n2924), .ZN(\mult_22/ab[31][40] ) );
  NOR2_X1 U10007 ( .A1(n2670), .A2(n2877), .ZN(\mult_22/ab[23][48] ) );
  NOR2_X1 U10008 ( .A1(n2682), .A2(n2865), .ZN(\mult_22/ab[21][50] ) );
  NOR2_X1 U10009 ( .A1(n2690), .A2(n2853), .ZN(\mult_22/ab[19][52] ) );
  NOR2_X1 U10010 ( .A1(n2704), .A2(n2842), .ZN(\mult_22/ab[17][54] ) );
  NOR2_X1 U10011 ( .A1(n2719), .A2(n2818), .ZN(\mult_22/ab[13][58] ) );
  NOR2_X1 U10012 ( .A1(n2546), .A2(n2815), .ZN(\mult_22/ab[13][27] ) );
  NOR2_X1 U10013 ( .A1(n2534), .A2(n2827), .ZN(\mult_22/ab[15][25] ) );
  NOR2_X1 U10014 ( .A1(n2522), .A2(n2839), .ZN(\mult_22/ab[17][23] ) );
  NOR2_X1 U10015 ( .A1(n2510), .A2(n2851), .ZN(\mult_22/ab[19][21] ) );
  NOR2_X1 U10016 ( .A1(n2498), .A2(n2862), .ZN(\mult_22/ab[21][19] ) );
  NOR2_X1 U10017 ( .A1(n2486), .A2(n2874), .ZN(\mult_22/ab[23][17] ) );
  NOR2_X1 U10018 ( .A1(n2473), .A2(n2886), .ZN(\mult_22/ab[25][15] ) );
  NOR2_X1 U10019 ( .A1(n2455), .A2(n2904), .ZN(\mult_22/ab[28][12] ) );
  NOR2_X1 U10020 ( .A1(n2441), .A2(n2916), .ZN(\mult_22/ab[30][10] ) );
  NOR2_X1 U10021 ( .A1(n2431), .A2(n2933), .ZN(\mult_22/ab[32][8] ) );
  NOR2_X1 U10022 ( .A1(n2419), .A2(n2945), .ZN(\mult_22/ab[34][6] ) );
  NOR2_X1 U10023 ( .A1(n2406), .A2(n2955), .ZN(\mult_22/ab[36][4] ) );
  NOR2_X1 U10024 ( .A1(n2550), .A2(n3001), .ZN(\mult_22/ab[44][28] ) );
  NOR2_X1 U10025 ( .A1(n2731), .A2(n2806), .ZN(\mult_22/ab[11][60] ) );
  NOR2_X1 U10026 ( .A1(n2540), .A2(n2815), .ZN(\mult_22/ab[13][26] ) );
  NOR2_X1 U10027 ( .A1(n2524), .A2(n2827), .ZN(\mult_22/ab[15][24] ) );
  NOR2_X1 U10028 ( .A1(n2516), .A2(n2839), .ZN(\mult_22/ab[17][22] ) );
  NOR2_X1 U10029 ( .A1(n2504), .A2(n2851), .ZN(\mult_22/ab[19][20] ) );
  NOR2_X1 U10030 ( .A1(n2492), .A2(n2862), .ZN(\mult_22/ab[21][18] ) );
  NOR2_X1 U10031 ( .A1(n2480), .A2(n2874), .ZN(\mult_22/ab[23][16] ) );
  NOR2_X1 U10032 ( .A1(n2467), .A2(n2886), .ZN(\mult_22/ab[25][14] ) );
  NOR2_X1 U10033 ( .A1(n2455), .A2(n2898), .ZN(\mult_22/ab[27][12] ) );
  NOR2_X1 U10034 ( .A1(n2441), .A2(n2910), .ZN(\mult_22/ab[29][10] ) );
  NOR2_X1 U10035 ( .A1(n2431), .A2(n2927), .ZN(\mult_22/ab[31][8] ) );
  NOR2_X1 U10036 ( .A1(n2419), .A2(n2938), .ZN(\mult_22/ab[33][6] ) );
  NOR2_X1 U10037 ( .A1(n2406), .A2(n2949), .ZN(\mult_22/ab[35][4] ) );
  NOR2_X1 U10038 ( .A1(n2554), .A2(n2779), .ZN(\mult_22/ab[7][29] ) );
  NOR2_X1 U10039 ( .A1(n2740), .A2(n2800), .ZN(\mult_22/ab[10][61] ) );
  NOR2_X1 U10040 ( .A1(n2556), .A2(n2995), .ZN(\mult_22/ab[43][29] ) );
  NOR2_X1 U10041 ( .A1(n2568), .A2(n2984), .ZN(\mult_22/ab[41][31] ) );
  NOR2_X1 U10042 ( .A1(n2579), .A2(n2972), .ZN(\mult_22/ab[39][33] ) );
  NOR2_X1 U10043 ( .A1(n2591), .A2(n2960), .ZN(\mult_22/ab[37][35] ) );
  NOR2_X1 U10044 ( .A1(n2604), .A2(n2948), .ZN(\mult_22/ab[35][37] ) );
  NOR2_X1 U10045 ( .A1(n2562), .A2(n2989), .ZN(\mult_22/ab[42][30] ) );
  NOR2_X1 U10046 ( .A1(n2574), .A2(n2978), .ZN(\mult_22/ab[40][32] ) );
  NOR2_X1 U10047 ( .A1(n2585), .A2(n2966), .ZN(\mult_22/ab[38][34] ) );
  NOR2_X1 U10048 ( .A1(n2597), .A2(n2954), .ZN(\mult_22/ab[36][36] ) );
  NOR2_X1 U10049 ( .A1(n2610), .A2(n2942), .ZN(\mult_22/ab[34][38] ) );
  NOR2_X1 U10050 ( .A1(n2547), .A2(n2803), .ZN(\mult_22/ab[11][27] ) );
  NOR2_X1 U10051 ( .A1(n2534), .A2(n2815), .ZN(\mult_22/ab[13][25] ) );
  NOR2_X1 U10052 ( .A1(n2522), .A2(n2827), .ZN(\mult_22/ab[15][23] ) );
  NOR2_X1 U10053 ( .A1(n2510), .A2(n2839), .ZN(\mult_22/ab[17][21] ) );
  NOR2_X1 U10054 ( .A1(n2498), .A2(n2850), .ZN(\mult_22/ab[19][19] ) );
  NOR2_X1 U10055 ( .A1(n2486), .A2(n2862), .ZN(\mult_22/ab[21][17] ) );
  NOR2_X1 U10056 ( .A1(n2474), .A2(n2874), .ZN(\mult_22/ab[23][15] ) );
  NOR2_X1 U10057 ( .A1(n2462), .A2(n2886), .ZN(\mult_22/ab[25][13] ) );
  NOR2_X1 U10058 ( .A1(n2449), .A2(n2898), .ZN(\mult_22/ab[27][11] ) );
  NOR2_X1 U10059 ( .A1(n2437), .A2(n2915), .ZN(\mult_22/ab[29][9] ) );
  NOR2_X1 U10060 ( .A1(n2425), .A2(n2927), .ZN(\mult_22/ab[31][7] ) );
  NOR2_X1 U10061 ( .A1(n2413), .A2(n2938), .ZN(\mult_22/ab[33][5] ) );
  NOR2_X1 U10062 ( .A1(n2554), .A2(n2773), .ZN(\mult_22/ab[6][29] ) );
  NOR2_X1 U10063 ( .A1(n2637), .A2(n2913), .ZN(\mult_22/ab[29][43] ) );
  NOR2_X1 U10064 ( .A1(n2625), .A2(n2924), .ZN(\mult_22/ab[31][41] ) );
  NOR2_X1 U10065 ( .A1(n2615), .A2(n2936), .ZN(\mult_22/ab[33][39] ) );
  NOR2_X1 U10066 ( .A1(n2649), .A2(n2901), .ZN(\mult_22/ab[27][45] ) );
  NOR2_X1 U10067 ( .A1(n2664), .A2(n2889), .ZN(\mult_22/ab[25][47] ) );
  NOR2_X1 U10068 ( .A1(n2673), .A2(n2877), .ZN(\mult_22/ab[23][49] ) );
  NOR2_X1 U10069 ( .A1(n2688), .A2(n2865), .ZN(\mult_22/ab[21][51] ) );
  NOR2_X1 U10070 ( .A1(n2700), .A2(n2854), .ZN(\mult_22/ab[19][53] ) );
  NOR2_X1 U10071 ( .A1(n2710), .A2(n2842), .ZN(\mult_22/ab[17][55] ) );
  NOR2_X1 U10072 ( .A1(n2716), .A2(n2830), .ZN(\mult_22/ab[15][57] ) );
  NOR2_X1 U10073 ( .A1(n2725), .A2(n2818), .ZN(\mult_22/ab[13][59] ) );
  NOR2_X1 U10074 ( .A1(n2541), .A2(n2803), .ZN(\mult_22/ab[11][26] ) );
  NOR2_X1 U10075 ( .A1(n2524), .A2(n2815), .ZN(\mult_22/ab[13][24] ) );
  NOR2_X1 U10076 ( .A1(n2516), .A2(n2827), .ZN(\mult_22/ab[15][22] ) );
  NOR2_X1 U10077 ( .A1(n2504), .A2(n2839), .ZN(\mult_22/ab[17][20] ) );
  NOR2_X1 U10078 ( .A1(n2492), .A2(n2850), .ZN(\mult_22/ab[19][18] ) );
  NOR2_X1 U10079 ( .A1(n2480), .A2(n2862), .ZN(\mult_22/ab[21][16] ) );
  NOR2_X1 U10080 ( .A1(n2468), .A2(n2874), .ZN(\mult_22/ab[23][14] ) );
  NOR2_X1 U10081 ( .A1(n2455), .A2(n2886), .ZN(\mult_22/ab[25][12] ) );
  NOR2_X1 U10082 ( .A1(n2441), .A2(n2898), .ZN(\mult_22/ab[27][10] ) );
  NOR2_X1 U10083 ( .A1(n2431), .A2(n2915), .ZN(\mult_22/ab[29][8] ) );
  NOR2_X1 U10084 ( .A1(n2419), .A2(n2927), .ZN(\mult_22/ab[31][6] ) );
  NOR2_X1 U10085 ( .A1(n2406), .A2(n2937), .ZN(\mult_22/ab[33][4] ) );
  NOR2_X1 U10086 ( .A1(n2645), .A2(n2907), .ZN(\mult_22/ab[28][44] ) );
  NOR2_X1 U10087 ( .A1(n2633), .A2(n2919), .ZN(\mult_22/ab[30][42] ) );
  NOR2_X1 U10088 ( .A1(n2621), .A2(n2930), .ZN(\mult_22/ab[32][40] ) );
  NOR2_X1 U10089 ( .A1(n2657), .A2(n2895), .ZN(\mult_22/ab[26][46] ) );
  NOR2_X1 U10090 ( .A1(n2670), .A2(n2883), .ZN(\mult_22/ab[24][48] ) );
  NOR2_X1 U10091 ( .A1(n2682), .A2(n2871), .ZN(\mult_22/ab[22][50] ) );
  NOR2_X1 U10092 ( .A1(n2690), .A2(n2859), .ZN(\mult_22/ab[20][52] ) );
  NOR2_X1 U10093 ( .A1(n2704), .A2(n2848), .ZN(\mult_22/ab[18][54] ) );
  NOR2_X1 U10094 ( .A1(n2719), .A2(n2824), .ZN(\mult_22/ab[14][58] ) );
  NOR2_X1 U10095 ( .A1(n2731), .A2(n2812), .ZN(\mult_22/ab[12][60] ) );
  NOR2_X1 U10096 ( .A1(n2741), .A2(n2806), .ZN(\mult_22/ab[11][61] ) );
  NOR2_X1 U10097 ( .A1(n2554), .A2(n2767), .ZN(\mult_22/ab[5][29] ) );
  NOR2_X1 U10098 ( .A1(n2542), .A2(n2791), .ZN(\mult_22/ab[9][27] ) );
  NOR2_X1 U10099 ( .A1(n2535), .A2(n2803), .ZN(\mult_22/ab[11][25] ) );
  NOR2_X1 U10100 ( .A1(n2522), .A2(n2815), .ZN(\mult_22/ab[13][23] ) );
  NOR2_X1 U10101 ( .A1(n2510), .A2(n2827), .ZN(\mult_22/ab[15][21] ) );
  NOR2_X1 U10102 ( .A1(n2498), .A2(n2838), .ZN(\mult_22/ab[17][19] ) );
  NOR2_X1 U10103 ( .A1(n2486), .A2(n2850), .ZN(\mult_22/ab[19][17] ) );
  NOR2_X1 U10104 ( .A1(n2474), .A2(n2862), .ZN(\mult_22/ab[21][15] ) );
  NOR2_X1 U10105 ( .A1(n2462), .A2(n2874), .ZN(\mult_22/ab[23][13] ) );
  NOR2_X1 U10106 ( .A1(n2449), .A2(n2886), .ZN(\mult_22/ab[25][11] ) );
  NOR2_X1 U10107 ( .A1(n2437), .A2(n2903), .ZN(\mult_22/ab[27][9] ) );
  NOR2_X1 U10108 ( .A1(n2425), .A2(n2915), .ZN(\mult_22/ab[29][7] ) );
  NOR2_X1 U10109 ( .A1(n2413), .A2(n2926), .ZN(\mult_22/ab[31][5] ) );
  NOR2_X1 U10110 ( .A1(n2537), .A2(n3019), .ZN(\mult_22/ab[47][26] ) );
  NOR2_X1 U10111 ( .A1(n2544), .A2(n3013), .ZN(\mult_22/ab[46][27] ) );
  NOR2_X1 U10112 ( .A1(n2550), .A2(n3007), .ZN(\mult_22/ab[45][28] ) );
  NOR2_X1 U10113 ( .A1(n2562), .A2(n2995), .ZN(\mult_22/ab[43][30] ) );
  NOR2_X1 U10114 ( .A1(n2574), .A2(n2984), .ZN(\mult_22/ab[41][32] ) );
  NOR2_X1 U10115 ( .A1(n2585), .A2(n2972), .ZN(\mult_22/ab[39][34] ) );
  NOR2_X1 U10116 ( .A1(n2597), .A2(n2960), .ZN(\mult_22/ab[37][36] ) );
  NOR2_X1 U10117 ( .A1(n2556), .A2(n3001), .ZN(\mult_22/ab[44][29] ) );
  NOR2_X1 U10118 ( .A1(n2568), .A2(n2990), .ZN(\mult_22/ab[42][31] ) );
  NOR2_X1 U10119 ( .A1(n2579), .A2(n2978), .ZN(\mult_22/ab[40][33] ) );
  NOR2_X1 U10120 ( .A1(n2591), .A2(n2966), .ZN(\mult_22/ab[38][35] ) );
  NOR2_X1 U10121 ( .A1(n2603), .A2(n2954), .ZN(\mult_22/ab[36][37] ) );
  NOR2_X1 U10122 ( .A1(n2610), .A2(n2948), .ZN(\mult_22/ab[35][38] ) );
  NOR2_X1 U10123 ( .A1(n2625), .A2(n2930), .ZN(\mult_22/ab[32][41] ) );
  NOR2_X1 U10124 ( .A1(n2615), .A2(n2942), .ZN(\mult_22/ab[34][39] ) );
  NOR2_X1 U10125 ( .A1(n2637), .A2(n2919), .ZN(\mult_22/ab[30][43] ) );
  NOR2_X1 U10126 ( .A1(n2649), .A2(n2907), .ZN(\mult_22/ab[28][45] ) );
  NOR2_X1 U10127 ( .A1(n2663), .A2(n2895), .ZN(\mult_22/ab[26][47] ) );
  NOR2_X1 U10128 ( .A1(n2673), .A2(n2883), .ZN(\mult_22/ab[24][49] ) );
  NOR2_X1 U10129 ( .A1(n2688), .A2(n2871), .ZN(\mult_22/ab[22][51] ) );
  NOR2_X1 U10130 ( .A1(n2367), .A2(n2860), .ZN(\mult_22/ab[20][53] ) );
  NOR2_X1 U10131 ( .A1(n2633), .A2(n2925), .ZN(\mult_22/ab[31][42] ) );
  NOR2_X1 U10132 ( .A1(n2621), .A2(n2936), .ZN(\mult_22/ab[33][40] ) );
  NOR2_X1 U10133 ( .A1(n2710), .A2(n2848), .ZN(\mult_22/ab[18][55] ) );
  NOR2_X1 U10134 ( .A1(n2645), .A2(n2913), .ZN(\mult_22/ab[29][44] ) );
  NOR2_X1 U10135 ( .A1(n2716), .A2(n2836), .ZN(\mult_22/ab[16][57] ) );
  NOR2_X1 U10136 ( .A1(n2657), .A2(n2901), .ZN(\mult_22/ab[27][46] ) );
  NOR2_X1 U10137 ( .A1(n2726), .A2(n2824), .ZN(\mult_22/ab[14][59] ) );
  NOR2_X1 U10138 ( .A1(n2669), .A2(n2889), .ZN(\mult_22/ab[25][48] ) );
  NOR2_X1 U10139 ( .A1(n2682), .A2(n2877), .ZN(\mult_22/ab[23][50] ) );
  NOR2_X1 U10140 ( .A1(n2690), .A2(n2865), .ZN(\mult_22/ab[21][52] ) );
  NOR2_X1 U10141 ( .A1(n2704), .A2(n2854), .ZN(\mult_22/ab[19][54] ) );
  NOR2_X1 U10142 ( .A1(n2719), .A2(n2830), .ZN(\mult_22/ab[15][58] ) );
  NOR2_X1 U10143 ( .A1(n2685), .A2(n2763), .ZN(\mult_22/ab[4][51] ) );
  NOR2_X1 U10144 ( .A1(n2392), .A2(n3109), .ZN(\mult_22/ab[62][2] ) );
  NOR2_X1 U10145 ( .A1(n2408), .A2(n3099), .ZN(\mult_22/ab[60][4] ) );
  NOR2_X1 U10146 ( .A1(n2398), .A2(n3104), .ZN(\mult_22/ab[61][3] ) );
  NOR2_X1 U10147 ( .A1(n2416), .A2(n3089), .ZN(\mult_22/ab[58][6] ) );
  NOR2_X1 U10148 ( .A1(n2408), .A2(n3093), .ZN(\mult_22/ab[59][4] ) );
  NOR2_X1 U10149 ( .A1(n2398), .A2(n3098), .ZN(\mult_22/ab[60][3] ) );
  NOR2_X1 U10150 ( .A1(n2392), .A2(n3103), .ZN(\mult_22/ab[61][2] ) );
  NOR2_X1 U10151 ( .A1(n2417), .A2(n3083), .ZN(\mult_22/ab[57][6] ) );
  NOR2_X1 U10152 ( .A1(n2386), .A2(n3108), .ZN(\mult_22/ab[62][1] ) );
  NOR2_X1 U10153 ( .A1(n2429), .A2(n3077), .ZN(\mult_22/ab[56][8] ) );
  NOR2_X1 U10154 ( .A1(n2408), .A2(n3087), .ZN(\mult_22/ab[58][4] ) );
  NOR2_X1 U10155 ( .A1(n2429), .A2(n3071), .ZN(\mult_22/ab[55][8] ) );
  NOR2_X1 U10156 ( .A1(n2417), .A2(n3077), .ZN(\mult_22/ab[56][6] ) );
  NOR2_X1 U10157 ( .A1(n2398), .A2(n3092), .ZN(\mult_22/ab[59][3] ) );
  NOR2_X1 U10158 ( .A1(n2392), .A2(n3097), .ZN(\mult_22/ab[60][2] ) );
  NOR2_X1 U10159 ( .A1(n2686), .A2(n2757), .ZN(\mult_22/ab[3][51] ) );
  NOR2_X1 U10160 ( .A1(n2443), .A2(n3060), .ZN(\mult_22/ab[54][10] ) );
  NOR2_X1 U10161 ( .A1(n2429), .A2(n3065), .ZN(\mult_22/ab[54][8] ) );
  NOR2_X1 U10162 ( .A1(n2417), .A2(n3071), .ZN(\mult_22/ab[55][6] ) );
  NOR2_X1 U10163 ( .A1(n2386), .A2(n3102), .ZN(\mult_22/ab[61][1] ) );
  NOR2_X1 U10164 ( .A1(n2624), .A2(n2834), .ZN(\mult_22/ab[16][41] ) );
  NOR2_X1 U10165 ( .A1(n2443), .A2(n3054), .ZN(\mult_22/ab[53][10] ) );
  NOR2_X1 U10166 ( .A1(n2408), .A2(n3081), .ZN(\mult_22/ab[57][4] ) );
  NOR2_X1 U10167 ( .A1(n2616), .A2(n2846), .ZN(\mult_22/ab[18][39] ) );
  NOR2_X1 U10168 ( .A1(n2429), .A2(n3059), .ZN(\mult_22/ab[53][8] ) );
  NOR2_X1 U10169 ( .A1(n2398), .A2(n3086), .ZN(\mult_22/ab[58][3] ) );
  NOR2_X1 U10170 ( .A1(n2443), .A2(n3048), .ZN(\mult_22/ab[52][10] ) );
  NOR2_X1 U10171 ( .A1(n2392), .A2(n3091), .ZN(\mult_22/ab[59][2] ) );
  NOR2_X1 U10172 ( .A1(n2622), .A2(n2834), .ZN(\mult_22/ab[16][40] ) );
  NOR2_X1 U10173 ( .A1(n2417), .A2(n3065), .ZN(\mult_22/ab[54][6] ) );
  NOR2_X1 U10174 ( .A1(n2611), .A2(n2852), .ZN(\mult_22/ab[19][38] ) );
  NOR2_X1 U10175 ( .A1(n2624), .A2(n2828), .ZN(\mult_22/ab[15][41] ) );
  NOR2_X1 U10176 ( .A1(n2453), .A2(n3042), .ZN(\mult_22/ab[51][12] ) );
  NOR2_X1 U10177 ( .A1(n2443), .A2(n3042), .ZN(\mult_22/ab[51][10] ) );
  NOR2_X1 U10178 ( .A1(n2429), .A2(n3053), .ZN(\mult_22/ab[52][8] ) );
  NOR2_X1 U10179 ( .A1(n2408), .A2(n3075), .ZN(\mult_22/ab[56][4] ) );
  NOR2_X1 U10180 ( .A1(n2465), .A2(n3042), .ZN(\mult_22/ab[51][14] ) );
  NOR2_X1 U10181 ( .A1(n2384), .A2(n3108), .ZN(\mult_22/ab[62][0] ) );
  NOR2_X1 U10182 ( .A1(n2386), .A2(n3096), .ZN(\mult_22/ab[60][1] ) );
  NOR2_X1 U10183 ( .A1(n2453), .A2(n3036), .ZN(\mult_22/ab[50][12] ) );
  NOR2_X1 U10184 ( .A1(n2399), .A2(n3080), .ZN(\mult_22/ab[57][3] ) );
  NOR2_X1 U10185 ( .A1(n2634), .A2(n2823), .ZN(\mult_22/ab[14][42] ) );
  NOR2_X1 U10186 ( .A1(n2443), .A2(n3036), .ZN(\mult_22/ab[50][10] ) );
  NOR2_X1 U10187 ( .A1(n2465), .A2(n3036), .ZN(\mult_22/ab[50][14] ) );
  NOR2_X1 U10188 ( .A1(n2417), .A2(n3059), .ZN(\mult_22/ab[53][6] ) );
  NOR2_X1 U10189 ( .A1(n2429), .A2(n3047), .ZN(\mult_22/ab[51][8] ) );
  NOR2_X1 U10190 ( .A1(n2453), .A2(n3030), .ZN(\mult_22/ab[49][12] ) );
  NOR2_X1 U10191 ( .A1(n2392), .A2(n3085), .ZN(\mult_22/ab[58][2] ) );
  NOR2_X1 U10192 ( .A1(n2624), .A2(n2822), .ZN(\mult_22/ab[14][41] ) );
  NOR2_X1 U10193 ( .A1(n2408), .A2(n3069), .ZN(\mult_22/ab[55][4] ) );
  NOR2_X1 U10194 ( .A1(n2622), .A2(n2828), .ZN(\mult_22/ab[15][40] ) );
  NOR2_X1 U10195 ( .A1(n2443), .A2(n3030), .ZN(\mult_22/ab[49][10] ) );
  NOR2_X1 U10196 ( .A1(n2453), .A2(n3024), .ZN(\mult_22/ab[48][12] ) );
  NOR2_X1 U10197 ( .A1(n2465), .A2(n3024), .ZN(\mult_22/ab[48][14] ) );
  NOR2_X1 U10198 ( .A1(n2635), .A2(n2817), .ZN(\mult_22/ab[13][42] ) );
  NOR2_X1 U10199 ( .A1(n2429), .A2(n3041), .ZN(\mult_22/ab[50][8] ) );
  NOR2_X1 U10200 ( .A1(n2417), .A2(n3053), .ZN(\mult_22/ab[52][6] ) );
  NOR2_X1 U10201 ( .A1(n2399), .A2(n3074), .ZN(\mult_22/ab[56][3] ) );
  NOR2_X1 U10202 ( .A1(n2465), .A2(n3018), .ZN(\mult_22/ab[47][14] ) );
  NOR2_X1 U10203 ( .A1(n2477), .A2(n3024), .ZN(\mult_22/ab[48][16] ) );
  NOR2_X1 U10204 ( .A1(n2443), .A2(n3024), .ZN(\mult_22/ab[48][10] ) );
  NOR2_X1 U10205 ( .A1(n2386), .A2(n3090), .ZN(\mult_22/ab[59][1] ) );
  NOR2_X1 U10206 ( .A1(n2453), .A2(n3018), .ZN(\mult_22/ab[47][12] ) );
  NOR2_X1 U10207 ( .A1(n2384), .A2(n3102), .ZN(\mult_22/ab[61][0] ) );
  NOR2_X1 U10208 ( .A1(n2407), .A2(n3063), .ZN(\mult_22/ab[54][4] ) );
  NOR2_X1 U10209 ( .A1(n2477), .A2(n3018), .ZN(\mult_22/ab[47][16] ) );
  NOR2_X1 U10210 ( .A1(n2393), .A2(n3079), .ZN(\mult_22/ab[57][2] ) );
  NOR2_X1 U10211 ( .A1(n2466), .A2(n3012), .ZN(\mult_22/ab[46][14] ) );
  NOR2_X1 U10212 ( .A1(n2624), .A2(n2816), .ZN(\mult_22/ab[13][41] ) );
  NOR2_X1 U10213 ( .A1(n2429), .A2(n3035), .ZN(\mult_22/ab[49][8] ) );
  NOR2_X1 U10214 ( .A1(n2454), .A2(n3012), .ZN(\mult_22/ab[46][12] ) );
  NOR2_X1 U10215 ( .A1(n2417), .A2(n3047), .ZN(\mult_22/ab[51][6] ) );
  NOR2_X1 U10216 ( .A1(n2478), .A2(n3012), .ZN(\mult_22/ab[46][16] ) );
  NOR2_X1 U10217 ( .A1(n2622), .A2(n2822), .ZN(\mult_22/ab[14][40] ) );
  NOR2_X1 U10218 ( .A1(n2635), .A2(n2811), .ZN(\mult_22/ab[12][42] ) );
  NOR2_X1 U10219 ( .A1(n2443), .A2(n3018), .ZN(\mult_22/ab[47][10] ) );
  NOR2_X1 U10220 ( .A1(n2647), .A2(n2811), .ZN(\mult_22/ab[12][44] ) );
  NOR2_X1 U10221 ( .A1(n2399), .A2(n3068), .ZN(\mult_22/ab[55][3] ) );
  NOR2_X1 U10222 ( .A1(n2466), .A2(n3006), .ZN(\mult_22/ab[45][14] ) );
  NOR2_X1 U10223 ( .A1(n2478), .A2(n3006), .ZN(\mult_22/ab[45][16] ) );
  NOR2_X1 U10224 ( .A1(n2490), .A2(n3012), .ZN(\mult_22/ab[46][18] ) );
  NOR2_X1 U10225 ( .A1(n2454), .A2(n3006), .ZN(\mult_22/ab[45][12] ) );
  NOR2_X1 U10226 ( .A1(n2647), .A2(n2805), .ZN(\mult_22/ab[11][44] ) );
  NOR2_X1 U10227 ( .A1(n2429), .A2(n3029), .ZN(\mult_22/ab[48][8] ) );
  NOR2_X1 U10228 ( .A1(n2407), .A2(n3057), .ZN(\mult_22/ab[53][4] ) );
  NOR2_X1 U10229 ( .A1(n2443), .A2(n3012), .ZN(\mult_22/ab[46][10] ) );
  NOR2_X1 U10230 ( .A1(n2466), .A2(n3000), .ZN(\mult_22/ab[44][14] ) );
  NOR2_X1 U10231 ( .A1(n2387), .A2(n3084), .ZN(\mult_22/ab[58][1] ) );
  NOR2_X1 U10232 ( .A1(n2478), .A2(n3000), .ZN(\mult_22/ab[44][16] ) );
  NOR2_X1 U10233 ( .A1(n2490), .A2(n3006), .ZN(\mult_22/ab[45][18] ) );
  NOR2_X1 U10234 ( .A1(n2417), .A2(n3041), .ZN(\mult_22/ab[50][6] ) );
  NOR2_X1 U10235 ( .A1(n2393), .A2(n3073), .ZN(\mult_22/ab[56][2] ) );
  NOR2_X1 U10236 ( .A1(n2624), .A2(n2810), .ZN(\mult_22/ab[12][41] ) );
  NOR2_X1 U10237 ( .A1(n2384), .A2(n3096), .ZN(\mult_22/ab[60][0] ) );
  NOR2_X1 U10238 ( .A1(n2490), .A2(n3000), .ZN(\mult_22/ab[44][18] ) );
  NOR2_X1 U10239 ( .A1(n2635), .A2(n2805), .ZN(\mult_22/ab[11][42] ) );
  NOR2_X1 U10240 ( .A1(n2454), .A2(n3000), .ZN(\mult_22/ab[44][12] ) );
  NOR2_X1 U10241 ( .A1(n2478), .A2(n2994), .ZN(\mult_22/ab[43][16] ) );
  NOR2_X1 U10242 ( .A1(n2399), .A2(n3062), .ZN(\mult_22/ab[54][3] ) );
  NOR2_X1 U10243 ( .A1(n2466), .A2(n2994), .ZN(\mult_22/ab[43][14] ) );
  NOR2_X1 U10244 ( .A1(n2622), .A2(n2816), .ZN(\mult_22/ab[13][40] ) );
  NOR2_X1 U10245 ( .A1(n2647), .A2(n2799), .ZN(\mult_22/ab[10][44] ) );
  NOR2_X1 U10246 ( .A1(n2436), .A2(n3017), .ZN(\mult_22/ab[46][9] ) );
  NOR2_X1 U10247 ( .A1(n2490), .A2(n2994), .ZN(\mult_22/ab[43][18] ) );
  NOR2_X1 U10248 ( .A1(n2423), .A2(n3029), .ZN(\mult_22/ab[48][7] ) );
  NOR2_X1 U10249 ( .A1(n2448), .A2(n3000), .ZN(\mult_22/ab[44][11] ) );
  NOR2_X1 U10250 ( .A1(n2407), .A2(n3051), .ZN(\mult_22/ab[52][4] ) );
  NOR2_X1 U10251 ( .A1(n2478), .A2(n2988), .ZN(\mult_22/ab[42][16] ) );
  NOR2_X1 U10252 ( .A1(n2466), .A2(n2988), .ZN(\mult_22/ab[42][14] ) );
  NOR2_X1 U10253 ( .A1(n2490), .A2(n2988), .ZN(\mult_22/ab[42][18] ) );
  NOR2_X1 U10254 ( .A1(n2387), .A2(n3078), .ZN(\mult_22/ab[57][1] ) );
  NOR2_X1 U10255 ( .A1(n2393), .A2(n3067), .ZN(\mult_22/ab[55][2] ) );
  NOR2_X1 U10256 ( .A1(n2502), .A2(n2995), .ZN(\mult_22/ab[43][20] ) );
  NOR2_X1 U10257 ( .A1(n2460), .A2(n2988), .ZN(\mult_22/ab[42][13] ) );
  NOR2_X1 U10258 ( .A1(n2478), .A2(n2982), .ZN(\mult_22/ab[41][16] ) );
  NOR2_X1 U10259 ( .A1(n2411), .A2(n3040), .ZN(\mult_22/ab[50][5] ) );
  NOR2_X1 U10260 ( .A1(n2642), .A2(n2793), .ZN(\mult_22/ab[9][44] ) );
  NOR2_X1 U10261 ( .A1(n2436), .A2(n3011), .ZN(\mult_22/ab[45][9] ) );
  NOR2_X1 U10262 ( .A1(n2490), .A2(n2982), .ZN(\mult_22/ab[41][18] ) );
  NOR2_X1 U10263 ( .A1(n2399), .A2(n3056), .ZN(\mult_22/ab[53][3] ) );
  NOR2_X1 U10264 ( .A1(n2624), .A2(n2804), .ZN(\mult_22/ab[11][41] ) );
  NOR2_X1 U10265 ( .A1(n2448), .A2(n2994), .ZN(\mult_22/ab[43][11] ) );
  NOR2_X1 U10266 ( .A1(n2635), .A2(n2799), .ZN(\mult_22/ab[10][42] ) );
  NOR2_X1 U10267 ( .A1(n2502), .A2(n2989), .ZN(\mult_22/ab[42][20] ) );
  NOR2_X1 U10268 ( .A1(n2423), .A2(n3023), .ZN(\mult_22/ab[47][7] ) );
  NOR2_X1 U10269 ( .A1(n2466), .A2(n2982), .ZN(\mult_22/ab[41][14] ) );
  NOR2_X1 U10270 ( .A1(n2622), .A2(n2810), .ZN(\mult_22/ab[12][40] ) );
  NOR2_X1 U10271 ( .A1(n2384), .A2(n3090), .ZN(\mult_22/ab[59][0] ) );
  NOR2_X1 U10272 ( .A1(n2654), .A2(n2793), .ZN(\mult_22/ab[9][46] ) );
  NOR2_X1 U10273 ( .A1(n2478), .A2(n2976), .ZN(\mult_22/ab[40][16] ) );
  NOR2_X1 U10274 ( .A1(n2502), .A2(n2983), .ZN(\mult_22/ab[41][20] ) );
  NOR2_X1 U10275 ( .A1(n2490), .A2(n2976), .ZN(\mult_22/ab[40][18] ) );
  NOR2_X1 U10276 ( .A1(n2460), .A2(n2982), .ZN(\mult_22/ab[41][13] ) );
  NOR2_X1 U10277 ( .A1(n2387), .A2(n3072), .ZN(\mult_22/ab[56][1] ) );
  NOR2_X1 U10278 ( .A1(n2393), .A2(n3061), .ZN(\mult_22/ab[54][2] ) );
  NOR2_X1 U10279 ( .A1(n2660), .A2(n2793), .ZN(\mult_22/ab[9][47] ) );
  NOR2_X1 U10280 ( .A1(n2502), .A2(n2977), .ZN(\mult_22/ab[40][20] ) );
  NOR2_X1 U10281 ( .A1(n2605), .A2(n2858), .ZN(\mult_22/ab[20][37] ) );
  NOR2_X1 U10282 ( .A1(n2411), .A2(n3034), .ZN(\mult_22/ab[49][5] ) );
  NOR2_X1 U10283 ( .A1(n2436), .A2(n3005), .ZN(\mult_22/ab[44][9] ) );
  NOR2_X1 U10284 ( .A1(n2466), .A2(n2976), .ZN(\mult_22/ab[40][14] ) );
  NOR2_X1 U10285 ( .A1(n2448), .A2(n2988), .ZN(\mult_22/ab[42][11] ) );
  NOR2_X1 U10286 ( .A1(n2490), .A2(n2970), .ZN(\mult_22/ab[39][18] ) );
  NOR2_X1 U10287 ( .A1(n2399), .A2(n3050), .ZN(\mult_22/ab[52][3] ) );
  NOR2_X1 U10288 ( .A1(n2514), .A2(n2989), .ZN(\mult_22/ab[42][22] ) );
  NOR2_X1 U10289 ( .A1(n2478), .A2(n2970), .ZN(\mult_22/ab[39][16] ) );
  NOR2_X1 U10290 ( .A1(n2424), .A2(n3017), .ZN(\mult_22/ab[46][7] ) );
  NOR2_X1 U10291 ( .A1(n2624), .A2(n2798), .ZN(\mult_22/ab[10][41] ) );
  NOR2_X1 U10292 ( .A1(n2654), .A2(n2787), .ZN(\mult_22/ab[8][46] ) );
  NOR2_X1 U10293 ( .A1(n2551), .A2(n2923), .ZN(\mult_22/ab[31][28] ) );
  NOR2_X1 U10294 ( .A1(n2642), .A2(n2787), .ZN(\mult_22/ab[8][44] ) );
  NOR2_X1 U10295 ( .A1(n2630), .A2(n2793), .ZN(\mult_22/ab[9][42] ) );
  NOR2_X1 U10296 ( .A1(n2586), .A2(n2882), .ZN(\mult_22/ab[24][34] ) );
  NOR2_X1 U10297 ( .A1(n2502), .A2(n2971), .ZN(\mult_22/ab[39][20] ) );
  NOR2_X1 U10298 ( .A1(n2573), .A2(n2870), .ZN(\mult_22/ab[22][32] ) );
  NOR2_X1 U10299 ( .A1(n2623), .A2(n2804), .ZN(\mult_22/ab[11][40] ) );
  NOR2_X1 U10300 ( .A1(n2460), .A2(n2976), .ZN(\mult_22/ab[40][13] ) );
  NOR2_X1 U10301 ( .A1(n2605), .A2(n2864), .ZN(\mult_22/ab[21][37] ) );
  NOR2_X1 U10302 ( .A1(n2387), .A2(n3066), .ZN(\mult_22/ab[55][1] ) );
  NOR2_X1 U10303 ( .A1(n2514), .A2(n2977), .ZN(\mult_22/ab[40][22] ) );
  NOR2_X1 U10304 ( .A1(n2490), .A2(n2964), .ZN(\mult_22/ab[38][18] ) );
  NOR2_X1 U10305 ( .A1(n2393), .A2(n3055), .ZN(\mult_22/ab[53][2] ) );
  NOR2_X1 U10306 ( .A1(n2411), .A2(n3028), .ZN(\mult_22/ab[48][5] ) );
  NOR2_X1 U10307 ( .A1(n2660), .A2(n2787), .ZN(\mult_22/ab[8][47] ) );
  NOR2_X1 U10308 ( .A1(n2436), .A2(n2999), .ZN(\mult_22/ab[43][9] ) );
  NOR2_X1 U10309 ( .A1(n2399), .A2(n3044), .ZN(\mult_22/ab[51][3] ) );
  NOR2_X1 U10310 ( .A1(n2526), .A2(n2959), .ZN(\mult_22/ab[37][24] ) );
  NOR2_X1 U10311 ( .A1(n2526), .A2(n2965), .ZN(\mult_22/ab[38][24] ) );
  NOR2_X1 U10312 ( .A1(n2514), .A2(n2971), .ZN(\mult_22/ab[39][22] ) );
  NOR2_X1 U10313 ( .A1(n2668), .A2(n2757), .ZN(\mult_22/ab[3][48] ) );
  NOR2_X1 U10314 ( .A1(n2667), .A2(n2763), .ZN(\mult_22/ab[4][48] ) );
  NOR2_X1 U10315 ( .A1(n2666), .A2(n2769), .ZN(\mult_22/ab[5][48] ) );
  NOR2_X1 U10316 ( .A1(n2666), .A2(n2775), .ZN(\mult_22/ab[6][48] ) );
  NOR2_X1 U10317 ( .A1(n2666), .A2(n2781), .ZN(\mult_22/ab[7][48] ) );
  NOR2_X1 U10318 ( .A1(n2666), .A2(n2787), .ZN(\mult_22/ab[8][48] ) );
  NOR2_X1 U10319 ( .A1(n2466), .A2(n2970), .ZN(\mult_22/ab[39][14] ) );
  NOR2_X1 U10320 ( .A1(n2448), .A2(n2982), .ZN(\mult_22/ab[41][11] ) );
  NOR2_X1 U10321 ( .A1(n2661), .A2(n2763), .ZN(\mult_22/ab[4][47] ) );
  NOR2_X1 U10322 ( .A1(n2660), .A2(n2769), .ZN(\mult_22/ab[5][47] ) );
  NOR2_X1 U10323 ( .A1(n2660), .A2(n2775), .ZN(\mult_22/ab[6][47] ) );
  NOR2_X1 U10324 ( .A1(n2660), .A2(n2781), .ZN(\mult_22/ab[7][47] ) );
  NOR2_X1 U10325 ( .A1(n2662), .A2(n2757), .ZN(\mult_22/ab[3][47] ) );
  NOR2_X1 U10326 ( .A1(n2631), .A2(n2763), .ZN(\mult_22/ab[4][42] ) );
  NOR2_X1 U10327 ( .A1(n2630), .A2(n2769), .ZN(\mult_22/ab[5][42] ) );
  NOR2_X1 U10328 ( .A1(n2630), .A2(n2775), .ZN(\mult_22/ab[6][42] ) );
  NOR2_X1 U10329 ( .A1(n2630), .A2(n2781), .ZN(\mult_22/ab[7][42] ) );
  NOR2_X1 U10330 ( .A1(n2630), .A2(n2787), .ZN(\mult_22/ab[8][42] ) );
  NOR2_X1 U10331 ( .A1(n2632), .A2(n2757), .ZN(\mult_22/ab[3][42] ) );
  NOR2_X1 U10332 ( .A1(n2628), .A2(n2768), .ZN(\mult_22/ab[5][41] ) );
  NOR2_X1 U10333 ( .A1(n2628), .A2(n2774), .ZN(\mult_22/ab[6][41] ) );
  NOR2_X1 U10334 ( .A1(n2628), .A2(n2780), .ZN(\mult_22/ab[7][41] ) );
  NOR2_X1 U10335 ( .A1(n2629), .A2(n2786), .ZN(\mult_22/ab[8][41] ) );
  NOR2_X1 U10336 ( .A1(n2629), .A2(n2792), .ZN(\mult_22/ab[9][41] ) );
  NOR2_X1 U10337 ( .A1(n2627), .A2(n2762), .ZN(\mult_22/ab[4][41] ) );
  NOR2_X1 U10338 ( .A1(n2654), .A2(n2775), .ZN(\mult_22/ab[6][46] ) );
  NOR2_X1 U10339 ( .A1(n2654), .A2(n2781), .ZN(\mult_22/ab[7][46] ) );
  NOR2_X1 U10340 ( .A1(n2654), .A2(n2769), .ZN(\mult_22/ab[5][46] ) );
  NOR2_X1 U10341 ( .A1(n2655), .A2(n2763), .ZN(\mult_22/ab[4][46] ) );
  NOR2_X1 U10342 ( .A1(n2642), .A2(n2781), .ZN(\mult_22/ab[7][44] ) );
  NOR2_X1 U10343 ( .A1(n2642), .A2(n2775), .ZN(\mult_22/ab[6][44] ) );
  NOR2_X1 U10344 ( .A1(n2618), .A2(n2780), .ZN(\mult_22/ab[7][40] ) );
  NOR2_X1 U10345 ( .A1(n2618), .A2(n2786), .ZN(\mult_22/ab[8][40] ) );
  NOR2_X1 U10346 ( .A1(n2618), .A2(n2792), .ZN(\mult_22/ab[9][40] ) );
  NOR2_X1 U10347 ( .A1(n2623), .A2(n2798), .ZN(\mult_22/ab[10][40] ) );
  NOR2_X1 U10348 ( .A1(n2618), .A2(n2774), .ZN(\mult_22/ab[6][40] ) );
  NOR2_X1 U10349 ( .A1(n2618), .A2(n2768), .ZN(\mult_22/ab[5][40] ) );
  NOR2_X1 U10350 ( .A1(n2626), .A2(n2756), .ZN(\mult_22/ab[3][41] ) );
  NOR2_X1 U10351 ( .A1(n2502), .A2(n2965), .ZN(\mult_22/ab[38][20] ) );
  NOR2_X1 U10352 ( .A1(n2611), .A2(n2810), .ZN(\mult_22/ab[12][38] ) );
  NOR2_X1 U10353 ( .A1(n2611), .A2(n2816), .ZN(\mult_22/ab[13][38] ) );
  NOR2_X1 U10354 ( .A1(n2599), .A2(n2816), .ZN(\mult_22/ab[13][36] ) );
  NOR2_X1 U10355 ( .A1(n2599), .A2(n2822), .ZN(\mult_22/ab[14][36] ) );
  NOR2_X1 U10356 ( .A1(n2599), .A2(n2828), .ZN(\mult_22/ab[15][36] ) );
  NOR2_X1 U10357 ( .A1(n2587), .A2(n2834), .ZN(\mult_22/ab[16][34] ) );
  NOR2_X1 U10358 ( .A1(n2599), .A2(n2834), .ZN(\mult_22/ab[16][36] ) );
  NOR2_X1 U10359 ( .A1(n2587), .A2(n2840), .ZN(\mult_22/ab[17][34] ) );
  NOR2_X1 U10360 ( .A1(n2587), .A2(n2846), .ZN(\mult_22/ab[18][34] ) );
  NOR2_X1 U10361 ( .A1(n2587), .A2(n2852), .ZN(\mult_22/ab[19][34] ) );
  NOR2_X1 U10362 ( .A1(n2607), .A2(n2792), .ZN(\mult_22/ab[9][38] ) );
  NOR2_X1 U10363 ( .A1(n2599), .A2(n2810), .ZN(\mult_22/ab[12][36] ) );
  NOR2_X1 U10364 ( .A1(n2587), .A2(n2828), .ZN(\mult_22/ab[15][34] ) );
  NOR2_X1 U10365 ( .A1(n2607), .A2(n2786), .ZN(\mult_22/ab[8][38] ) );
  NOR2_X1 U10366 ( .A1(n2600), .A2(n2804), .ZN(\mult_22/ab[11][36] ) );
  NOR2_X1 U10367 ( .A1(n2587), .A2(n2822), .ZN(\mult_22/ab[14][34] ) );
  NOR2_X1 U10368 ( .A1(n2607), .A2(n2780), .ZN(\mult_22/ab[7][38] ) );
  NOR2_X1 U10369 ( .A1(n2600), .A2(n2798), .ZN(\mult_22/ab[10][36] ) );
  NOR2_X1 U10370 ( .A1(n2587), .A2(n2816), .ZN(\mult_22/ab[13][34] ) );
  NOR2_X1 U10371 ( .A1(n2595), .A2(n2792), .ZN(\mult_22/ab[9][36] ) );
  NOR2_X1 U10372 ( .A1(n2587), .A2(n2810), .ZN(\mult_22/ab[12][34] ) );
  NOR2_X1 U10373 ( .A1(n2588), .A2(n2804), .ZN(\mult_22/ab[11][34] ) );
  NOR2_X1 U10374 ( .A1(n2619), .A2(n2762), .ZN(\mult_22/ab[4][40] ) );
  NOR2_X1 U10375 ( .A1(n2620), .A2(n2756), .ZN(\mult_22/ab[3][40] ) );
  NOR2_X1 U10376 ( .A1(n2678), .A2(n2769), .ZN(\mult_22/ab[5][50] ) );
  NOR2_X1 U10377 ( .A1(n2679), .A2(n2763), .ZN(\mult_22/ab[4][50] ) );
  NOR2_X1 U10378 ( .A1(n2612), .A2(n2768), .ZN(\mult_22/ab[5][39] ) );
  NOR2_X1 U10379 ( .A1(n2613), .A2(n2762), .ZN(\mult_22/ab[4][39] ) );
  NOR2_X1 U10380 ( .A1(n2601), .A2(n2780), .ZN(\mult_22/ab[7][37] ) );
  NOR2_X1 U10381 ( .A1(n2601), .A2(n2774), .ZN(\mult_22/ab[6][37] ) );
  NOR2_X1 U10382 ( .A1(n2589), .A2(n2792), .ZN(\mult_22/ab[9][35] ) );
  NOR2_X1 U10383 ( .A1(n2589), .A2(n2786), .ZN(\mult_22/ab[8][35] ) );
  NOR2_X1 U10384 ( .A1(n2676), .A2(n2775), .ZN(\mult_22/ab[6][49] ) );
  NOR2_X1 U10385 ( .A1(n2676), .A2(n2769), .ZN(\mult_22/ab[5][49] ) );
  NOR2_X1 U10386 ( .A1(n2582), .A2(n2804), .ZN(\mult_22/ab[11][33] ) );
  NOR2_X1 U10387 ( .A1(n2582), .A2(n2798), .ZN(\mult_22/ab[10][33] ) );
  NOR2_X1 U10388 ( .A1(n2656), .A2(n2757), .ZN(\mult_22/ab[3][46] ) );
  NOR2_X1 U10389 ( .A1(n2642), .A2(n2769), .ZN(\mult_22/ab[5][44] ) );
  NOR2_X1 U10390 ( .A1(n2643), .A2(n2763), .ZN(\mult_22/ab[4][44] ) );
  NOR2_X1 U10391 ( .A1(n2638), .A2(n2757), .ZN(\mult_22/ab[3][43] ) );
  NOR2_X1 U10392 ( .A1(n2639), .A2(n2763), .ZN(\mult_22/ab[4][43] ) );
  NOR2_X1 U10393 ( .A1(n2644), .A2(n2757), .ZN(\mult_22/ab[3][44] ) );
  NOR2_X1 U10394 ( .A1(n2680), .A2(n2757), .ZN(\mult_22/ab[3][50] ) );
  NOR2_X1 U10395 ( .A1(n2573), .A2(n2900), .ZN(\mult_22/ab[27][32] ) );
  NOR2_X1 U10396 ( .A1(n2539), .A2(n2941), .ZN(\mult_22/ab[34][26] ) );
  NOR2_X1 U10397 ( .A1(n2526), .A2(n2953), .ZN(\mult_22/ab[36][24] ) );
  NOR2_X1 U10398 ( .A1(n2514), .A2(n2965), .ZN(\mult_22/ab[38][22] ) );
  NOR2_X1 U10399 ( .A1(n2608), .A2(n2762), .ZN(\mult_22/ab[4][38] ) );
  NOR2_X1 U10400 ( .A1(n2595), .A2(n2774), .ZN(\mult_22/ab[6][36] ) );
  NOR2_X1 U10401 ( .A1(n2583), .A2(n2786), .ZN(\mult_22/ab[8][34] ) );
  NOR2_X1 U10402 ( .A1(n2572), .A2(n2852), .ZN(\mult_22/ab[19][32] ) );
  NOR2_X1 U10403 ( .A1(n2572), .A2(n2858), .ZN(\mult_22/ab[20][32] ) );
  NOR2_X1 U10404 ( .A1(n2572), .A2(n2864), .ZN(\mult_22/ab[21][32] ) );
  NOR2_X1 U10405 ( .A1(n2572), .A2(n2846), .ZN(\mult_22/ab[18][32] ) );
  NOR2_X1 U10406 ( .A1(n2572), .A2(n2840), .ZN(\mult_22/ab[17][32] ) );
  NOR2_X1 U10407 ( .A1(n2572), .A2(n2834), .ZN(\mult_22/ab[16][32] ) );
  NOR2_X1 U10408 ( .A1(n2572), .A2(n2828), .ZN(\mult_22/ab[15][32] ) );
  NOR2_X1 U10409 ( .A1(n2572), .A2(n2822), .ZN(\mult_22/ab[14][32] ) );
  NOR2_X1 U10410 ( .A1(n2572), .A2(n2816), .ZN(\mult_22/ab[13][32] ) );
  NOR2_X1 U10411 ( .A1(n2674), .A2(n2757), .ZN(\mult_22/ab[3][49] ) );
  NOR2_X1 U10412 ( .A1(n2572), .A2(n2810), .ZN(\mult_22/ab[12][32] ) );
  NOR2_X1 U10413 ( .A1(n2572), .A2(n2804), .ZN(\mult_22/ab[11][32] ) );
  NOR2_X1 U10414 ( .A1(n2733), .A2(n2758), .ZN(\mult_22/ab[3][60] ) );
  NOR2_X1 U10415 ( .A1(n2690), .A2(n2805), .ZN(\mult_22/ab[11][52] ) );
  NOR2_X1 U10416 ( .A1(n2682), .A2(n2817), .ZN(\mult_22/ab[13][50] ) );
  NOR2_X1 U10417 ( .A1(n2670), .A2(n2829), .ZN(\mult_22/ab[15][48] ) );
  NOR2_X1 U10418 ( .A1(n2658), .A2(n2841), .ZN(\mult_22/ab[17][46] ) );
  NOR2_X1 U10419 ( .A1(n2646), .A2(n2853), .ZN(\mult_22/ab[19][44] ) );
  NOR2_X1 U10420 ( .A1(n2634), .A2(n2864), .ZN(\mult_22/ab[21][42] ) );
  NOR2_X1 U10421 ( .A1(n2622), .A2(n2876), .ZN(\mult_22/ab[23][40] ) );
  NOR2_X1 U10422 ( .A1(n2602), .A2(n2762), .ZN(\mult_22/ab[4][37] ) );
  NOR2_X1 U10423 ( .A1(n2589), .A2(n2774), .ZN(\mult_22/ab[6][35] ) );
  NOR2_X1 U10424 ( .A1(n2577), .A2(n2786), .ZN(\mult_22/ab[8][33] ) );
  NOR2_X1 U10425 ( .A1(n2539), .A2(n2935), .ZN(\mult_22/ab[33][26] ) );
  NOR2_X1 U10426 ( .A1(n2539), .A2(n2929), .ZN(\mult_22/ab[32][26] ) );
  NOR2_X1 U10427 ( .A1(n2526), .A2(n2947), .ZN(\mult_22/ab[35][24] ) );
  NOR2_X1 U10428 ( .A1(n2526), .A2(n2941), .ZN(\mult_22/ab[34][24] ) );
  NOR2_X1 U10429 ( .A1(n2514), .A2(n2959), .ZN(\mult_22/ab[37][22] ) );
  NOR2_X1 U10430 ( .A1(n2514), .A2(n2953), .ZN(\mult_22/ab[36][22] ) );
  NOR2_X1 U10431 ( .A1(n2572), .A2(n2798), .ZN(\mult_22/ab[10][32] ) );
  NOR2_X1 U10432 ( .A1(n2571), .A2(n2816), .ZN(\mult_22/ab[13][31] ) );
  NOR2_X1 U10433 ( .A1(n2571), .A2(n2810), .ZN(\mult_22/ab[12][31] ) );
  NOR2_X1 U10434 ( .A1(n2596), .A2(n2762), .ZN(\mult_22/ab[4][36] ) );
  NOR2_X1 U10435 ( .A1(n2583), .A2(n2774), .ZN(\mult_22/ab[6][34] ) );
  NOR2_X1 U10436 ( .A1(n2590), .A2(n2762), .ZN(\mult_22/ab[4][35] ) );
  NOR2_X1 U10437 ( .A1(n2577), .A2(n2774), .ZN(\mult_22/ab[6][33] ) );
  NOR2_X1 U10438 ( .A1(n2718), .A2(n2770), .ZN(\mult_22/ab[5][57] ) );
  NOR2_X1 U10439 ( .A1(n2664), .A2(n2829), .ZN(\mult_22/ab[15][47] ) );
  NOR2_X1 U10440 ( .A1(n2648), .A2(n2841), .ZN(\mult_22/ab[17][45] ) );
  NOR2_X1 U10441 ( .A1(n2636), .A2(n2853), .ZN(\mult_22/ab[19][43] ) );
  NOR2_X1 U10442 ( .A1(n2624), .A2(n2864), .ZN(\mult_22/ab[21][41] ) );
  NOR2_X1 U10443 ( .A1(n2616), .A2(n2876), .ZN(\mult_22/ab[23][39] ) );
  NOR2_X1 U10444 ( .A1(n2424), .A2(n3011), .ZN(\mult_22/ab[45][7] ) );
  NOR2_X1 U10445 ( .A1(n2551), .A2(n2911), .ZN(\mult_22/ab[29][28] ) );
  NOR2_X1 U10446 ( .A1(n2551), .A2(n2905), .ZN(\mult_22/ab[28][28] ) );
  NOR2_X1 U10447 ( .A1(n2564), .A2(n2869), .ZN(\mult_22/ab[22][30] ) );
  NOR2_X1 U10448 ( .A1(n2564), .A2(n2875), .ZN(\mult_22/ab[23][30] ) );
  NOR2_X1 U10449 ( .A1(n2563), .A2(n2881), .ZN(\mult_22/ab[24][30] ) );
  NOR2_X1 U10450 ( .A1(n2563), .A2(n2887), .ZN(\mult_22/ab[25][30] ) );
  NOR2_X1 U10451 ( .A1(n2564), .A2(n2864), .ZN(\mult_22/ab[21][30] ) );
  NOR2_X1 U10452 ( .A1(n2564), .A2(n2857), .ZN(\mult_22/ab[20][30] ) );
  NOR2_X1 U10453 ( .A1(n2564), .A2(n2851), .ZN(\mult_22/ab[19][30] ) );
  NOR2_X1 U10454 ( .A1(n2564), .A2(n2845), .ZN(\mult_22/ab[18][30] ) );
  NOR2_X1 U10455 ( .A1(n2564), .A2(n2839), .ZN(\mult_22/ab[17][30] ) );
  NOR2_X1 U10456 ( .A1(n2564), .A2(n2833), .ZN(\mult_22/ab[16][30] ) );
  NOR2_X1 U10457 ( .A1(n2564), .A2(n2827), .ZN(\mult_22/ab[15][30] ) );
  NOR2_X1 U10458 ( .A1(n2478), .A2(n2964), .ZN(\mult_22/ab[38][16] ) );
  NOR2_X1 U10459 ( .A1(n2584), .A2(n2762), .ZN(\mult_22/ab[4][34] ) );
  NOR2_X1 U10460 ( .A1(n2576), .A2(n2786), .ZN(\mult_22/ab[8][32] ) );
  NOR2_X1 U10461 ( .A1(n2564), .A2(n2821), .ZN(\mult_22/ab[14][30] ) );
  NOR2_X1 U10462 ( .A1(n2564), .A2(n2815), .ZN(\mult_22/ab[13][30] ) );
  NOR2_X1 U10463 ( .A1(n2576), .A2(n2780), .ZN(\mult_22/ab[7][32] ) );
  NOR2_X1 U10464 ( .A1(n2571), .A2(n2798), .ZN(\mult_22/ab[10][31] ) );
  NOR2_X1 U10465 ( .A1(n2539), .A2(n2923), .ZN(\mult_22/ab[31][26] ) );
  NOR2_X1 U10466 ( .A1(n2539), .A2(n2917), .ZN(\mult_22/ab[30][26] ) );
  NOR2_X1 U10467 ( .A1(n2526), .A2(n2935), .ZN(\mult_22/ab[33][24] ) );
  NOR2_X1 U10468 ( .A1(n2525), .A2(n2929), .ZN(\mult_22/ab[32][24] ) );
  NOR2_X1 U10469 ( .A1(n2515), .A2(n2947), .ZN(\mult_22/ab[35][22] ) );
  NOR2_X1 U10470 ( .A1(n2515), .A2(n2941), .ZN(\mult_22/ab[34][22] ) );
  NOR2_X1 U10471 ( .A1(n2502), .A2(n2959), .ZN(\mult_22/ab[37][20] ) );
  NOR2_X1 U10472 ( .A1(n2502), .A2(n2953), .ZN(\mult_22/ab[36][20] ) );
  NOR2_X1 U10473 ( .A1(n2564), .A2(n2809), .ZN(\mult_22/ab[12][30] ) );
  NOR2_X1 U10474 ( .A1(n2578), .A2(n2762), .ZN(\mult_22/ab[4][33] ) );
  NOR2_X1 U10475 ( .A1(n2576), .A2(n2774), .ZN(\mult_22/ab[6][32] ) );
  NOR2_X1 U10476 ( .A1(n2566), .A2(n2786), .ZN(\mult_22/ab[8][31] ) );
  NOR2_X1 U10477 ( .A1(n2565), .A2(n2803), .ZN(\mult_22/ab[11][30] ) );
  NOR2_X1 U10478 ( .A1(n2576), .A2(n2768), .ZN(\mult_22/ab[5][32] ) );
  NOR2_X1 U10479 ( .A1(n2551), .A2(n2887), .ZN(\mult_22/ab[25][28] ) );
  NOR2_X1 U10480 ( .A1(n2551), .A2(n2893), .ZN(\mult_22/ab[26][28] ) );
  NOR2_X1 U10481 ( .A1(n2551), .A2(n2899), .ZN(\mult_22/ab[27][28] ) );
  NOR2_X1 U10482 ( .A1(n2551), .A2(n2881), .ZN(\mult_22/ab[24][28] ) );
  NOR2_X1 U10483 ( .A1(n2552), .A2(n2875), .ZN(\mult_22/ab[23][28] ) );
  NOR2_X1 U10484 ( .A1(n2552), .A2(n2869), .ZN(\mult_22/ab[22][28] ) );
  NOR2_X1 U10485 ( .A1(n2552), .A2(n2863), .ZN(\mult_22/ab[21][28] ) );
  NOR2_X1 U10486 ( .A1(n2552), .A2(n2857), .ZN(\mult_22/ab[20][28] ) );
  NOR2_X1 U10487 ( .A1(n2552), .A2(n2851), .ZN(\mult_22/ab[19][28] ) );
  NOR2_X1 U10488 ( .A1(n2552), .A2(n2845), .ZN(\mult_22/ab[18][28] ) );
  NOR2_X1 U10489 ( .A1(n2552), .A2(n2839), .ZN(\mult_22/ab[17][28] ) );
  NOR2_X1 U10490 ( .A1(n2552), .A2(n2833), .ZN(\mult_22/ab[16][28] ) );
  NOR2_X1 U10491 ( .A1(n2552), .A2(n2827), .ZN(\mult_22/ab[15][28] ) );
  NOR2_X1 U10492 ( .A1(n2575), .A2(n2762), .ZN(\mult_22/ab[4][32] ) );
  NOR2_X1 U10493 ( .A1(n2565), .A2(n2797), .ZN(\mult_22/ab[10][30] ) );
  NOR2_X1 U10494 ( .A1(n2560), .A2(n2791), .ZN(\mult_22/ab[9][30] ) );
  NOR2_X1 U10495 ( .A1(n2552), .A2(n2821), .ZN(\mult_22/ab[14][28] ) );
  NOR2_X1 U10496 ( .A1(n2539), .A2(n2905), .ZN(\mult_22/ab[28][26] ) );
  NOR2_X1 U10497 ( .A1(n2539), .A2(n2911), .ZN(\mult_22/ab[29][26] ) );
  NOR2_X1 U10498 ( .A1(n2525), .A2(n2923), .ZN(\mult_22/ab[31][24] ) );
  NOR2_X1 U10499 ( .A1(n2539), .A2(n2899), .ZN(\mult_22/ab[27][26] ) );
  NOR2_X1 U10500 ( .A1(n2525), .A2(n2917), .ZN(\mult_22/ab[30][24] ) );
  NOR2_X1 U10501 ( .A1(n2515), .A2(n2935), .ZN(\mult_22/ab[33][22] ) );
  NOR2_X1 U10502 ( .A1(n2539), .A2(n2893), .ZN(\mult_22/ab[26][26] ) );
  NOR2_X1 U10503 ( .A1(n2525), .A2(n2911), .ZN(\mult_22/ab[29][24] ) );
  NOR2_X1 U10504 ( .A1(n2515), .A2(n2929), .ZN(\mult_22/ab[32][22] ) );
  NOR2_X1 U10505 ( .A1(n2503), .A2(n2947), .ZN(\mult_22/ab[35][20] ) );
  NOR2_X1 U10506 ( .A1(n2539), .A2(n2887), .ZN(\mult_22/ab[25][26] ) );
  NOR2_X1 U10507 ( .A1(n2525), .A2(n2905), .ZN(\mult_22/ab[28][24] ) );
  NOR2_X1 U10508 ( .A1(n2515), .A2(n2923), .ZN(\mult_22/ab[31][22] ) );
  NOR2_X1 U10509 ( .A1(n2503), .A2(n2941), .ZN(\mult_22/ab[34][20] ) );
  NOR2_X1 U10510 ( .A1(n2490), .A2(n2958), .ZN(\mult_22/ab[37][18] ) );
  NOR2_X1 U10511 ( .A1(n2540), .A2(n2881), .ZN(\mult_22/ab[24][26] ) );
  NOR2_X1 U10512 ( .A1(n2525), .A2(n2899), .ZN(\mult_22/ab[27][24] ) );
  NOR2_X1 U10513 ( .A1(n2515), .A2(n2917), .ZN(\mult_22/ab[30][22] ) );
  NOR2_X1 U10514 ( .A1(n2503), .A2(n2935), .ZN(\mult_22/ab[33][20] ) );
  NOR2_X1 U10515 ( .A1(n2490), .A2(n2952), .ZN(\mult_22/ab[36][18] ) );
  NOR2_X1 U10516 ( .A1(n2540), .A2(n2875), .ZN(\mult_22/ab[23][26] ) );
  NOR2_X1 U10517 ( .A1(n2525), .A2(n2893), .ZN(\mult_22/ab[26][24] ) );
  NOR2_X1 U10518 ( .A1(n2515), .A2(n2911), .ZN(\mult_22/ab[29][22] ) );
  NOR2_X1 U10519 ( .A1(n2503), .A2(n2929), .ZN(\mult_22/ab[32][20] ) );
  NOR2_X1 U10520 ( .A1(n2491), .A2(n2946), .ZN(\mult_22/ab[35][18] ) );
  NOR2_X1 U10521 ( .A1(n2540), .A2(n2869), .ZN(\mult_22/ab[22][26] ) );
  NOR2_X1 U10522 ( .A1(n2525), .A2(n2887), .ZN(\mult_22/ab[25][24] ) );
  NOR2_X1 U10523 ( .A1(n2515), .A2(n2905), .ZN(\mult_22/ab[28][22] ) );
  NOR2_X1 U10524 ( .A1(n2503), .A2(n2923), .ZN(\mult_22/ab[31][20] ) );
  NOR2_X1 U10525 ( .A1(n2491), .A2(n2940), .ZN(\mult_22/ab[34][18] ) );
  NOR2_X1 U10526 ( .A1(n2540), .A2(n2863), .ZN(\mult_22/ab[21][26] ) );
  NOR2_X1 U10527 ( .A1(n2525), .A2(n2881), .ZN(\mult_22/ab[24][24] ) );
  NOR2_X1 U10528 ( .A1(n2515), .A2(n2899), .ZN(\mult_22/ab[27][22] ) );
  NOR2_X1 U10529 ( .A1(n2503), .A2(n2917), .ZN(\mult_22/ab[30][20] ) );
  NOR2_X1 U10530 ( .A1(n2491), .A2(n2934), .ZN(\mult_22/ab[33][18] ) );
  NOR2_X1 U10531 ( .A1(n2540), .A2(n2857), .ZN(\mult_22/ab[20][26] ) );
  NOR2_X1 U10532 ( .A1(n2525), .A2(n2875), .ZN(\mult_22/ab[23][24] ) );
  NOR2_X1 U10533 ( .A1(n2515), .A2(n2893), .ZN(\mult_22/ab[26][22] ) );
  NOR2_X1 U10534 ( .A1(n2503), .A2(n2911), .ZN(\mult_22/ab[29][20] ) );
  NOR2_X1 U10535 ( .A1(n2491), .A2(n2928), .ZN(\mult_22/ab[32][18] ) );
  NOR2_X1 U10536 ( .A1(n2540), .A2(n2851), .ZN(\mult_22/ab[19][26] ) );
  NOR2_X1 U10537 ( .A1(n2525), .A2(n2869), .ZN(\mult_22/ab[22][24] ) );
  NOR2_X1 U10538 ( .A1(n2515), .A2(n2887), .ZN(\mult_22/ab[25][22] ) );
  NOR2_X1 U10539 ( .A1(n2503), .A2(n2905), .ZN(\mult_22/ab[28][20] ) );
  NOR2_X1 U10540 ( .A1(n2491), .A2(n2922), .ZN(\mult_22/ab[31][18] ) );
  NOR2_X1 U10541 ( .A1(n2478), .A2(n2958), .ZN(\mult_22/ab[37][16] ) );
  NOR2_X1 U10542 ( .A1(n2524), .A2(n2863), .ZN(\mult_22/ab[21][24] ) );
  NOR2_X1 U10543 ( .A1(n2516), .A2(n2881), .ZN(\mult_22/ab[24][22] ) );
  NOR2_X1 U10544 ( .A1(n2503), .A2(n2899), .ZN(\mult_22/ab[27][20] ) );
  NOR2_X1 U10545 ( .A1(n2491), .A2(n2916), .ZN(\mult_22/ab[30][18] ) );
  NOR2_X1 U10546 ( .A1(n2478), .A2(n2952), .ZN(\mult_22/ab[36][16] ) );
  NOR2_X1 U10547 ( .A1(n2516), .A2(n2875), .ZN(\mult_22/ab[23][22] ) );
  NOR2_X1 U10548 ( .A1(n2503), .A2(n2893), .ZN(\mult_22/ab[26][20] ) );
  NOR2_X1 U10549 ( .A1(n2491), .A2(n2910), .ZN(\mult_22/ab[29][18] ) );
  NOR2_X1 U10550 ( .A1(n2479), .A2(n2946), .ZN(\mult_22/ab[35][16] ) );
  NOR2_X1 U10551 ( .A1(n2503), .A2(n2887), .ZN(\mult_22/ab[25][20] ) );
  NOR2_X1 U10552 ( .A1(n2491), .A2(n2904), .ZN(\mult_22/ab[28][18] ) );
  NOR2_X1 U10553 ( .A1(n2479), .A2(n2940), .ZN(\mult_22/ab[34][16] ) );
  NOR2_X1 U10554 ( .A1(n2491), .A2(n2898), .ZN(\mult_22/ab[27][18] ) );
  NOR2_X1 U10555 ( .A1(n2479), .A2(n2934), .ZN(\mult_22/ab[33][16] ) );
  NOR2_X1 U10556 ( .A1(n2479), .A2(n2928), .ZN(\mult_22/ab[32][16] ) );
  NOR2_X1 U10557 ( .A1(n2479), .A2(n2922), .ZN(\mult_22/ab[31][16] ) );
  NOR2_X1 U10558 ( .A1(n2479), .A2(n2916), .ZN(\mult_22/ab[30][16] ) );
  NOR2_X1 U10559 ( .A1(n2479), .A2(n2910), .ZN(\mult_22/ab[29][16] ) );
  NOR2_X1 U10560 ( .A1(n2466), .A2(n2964), .ZN(\mult_22/ab[38][14] ) );
  NOR2_X1 U10561 ( .A1(n2466), .A2(n2958), .ZN(\mult_22/ab[37][14] ) );
  NOR2_X1 U10562 ( .A1(n2466), .A2(n2952), .ZN(\mult_22/ab[36][14] ) );
  NOR2_X1 U10563 ( .A1(n2467), .A2(n2946), .ZN(\mult_22/ab[35][14] ) );
  NOR2_X1 U10564 ( .A1(n2467), .A2(n2940), .ZN(\mult_22/ab[34][14] ) );
  NOR2_X1 U10565 ( .A1(n2467), .A2(n2934), .ZN(\mult_22/ab[33][14] ) );
  NOR2_X1 U10566 ( .A1(n2460), .A2(n2970), .ZN(\mult_22/ab[39][13] ) );
  NOR2_X1 U10567 ( .A1(n2467), .A2(n2928), .ZN(\mult_22/ab[32][14] ) );
  NOR2_X1 U10568 ( .A1(n2546), .A2(n2839), .ZN(\mult_22/ab[17][27] ) );
  NOR2_X1 U10569 ( .A1(n2460), .A2(n2964), .ZN(\mult_22/ab[38][13] ) );
  NOR2_X1 U10570 ( .A1(n2467), .A2(n2922), .ZN(\mult_22/ab[31][14] ) );
  NOR2_X1 U10571 ( .A1(n2546), .A2(n2833), .ZN(\mult_22/ab[16][27] ) );
  NOR2_X1 U10572 ( .A1(n2534), .A2(n2851), .ZN(\mult_22/ab[19][25] ) );
  NOR2_X1 U10573 ( .A1(n2460), .A2(n2958), .ZN(\mult_22/ab[37][13] ) );
  NOR2_X1 U10574 ( .A1(n2448), .A2(n2976), .ZN(\mult_22/ab[40][11] ) );
  NOR2_X1 U10575 ( .A1(n2534), .A2(n2845), .ZN(\mult_22/ab[18][25] ) );
  NOR2_X1 U10576 ( .A1(n2522), .A2(n2863), .ZN(\mult_22/ab[21][23] ) );
  NOR2_X1 U10577 ( .A1(n2461), .A2(n2952), .ZN(\mult_22/ab[36][13] ) );
  NOR2_X1 U10578 ( .A1(n2448), .A2(n2970), .ZN(\mult_22/ab[39][11] ) );
  NOR2_X1 U10579 ( .A1(n2436), .A2(n2993), .ZN(\mult_22/ab[42][9] ) );
  NOR2_X1 U10580 ( .A1(n2522), .A2(n2857), .ZN(\mult_22/ab[20][23] ) );
  NOR2_X1 U10581 ( .A1(n2510), .A2(n2875), .ZN(\mult_22/ab[23][21] ) );
  NOR2_X1 U10582 ( .A1(n2461), .A2(n2946), .ZN(\mult_22/ab[35][13] ) );
  NOR2_X1 U10583 ( .A1(n2448), .A2(n2964), .ZN(\mult_22/ab[38][11] ) );
  NOR2_X1 U10584 ( .A1(n2436), .A2(n2987), .ZN(\mult_22/ab[41][9] ) );
  NOR2_X1 U10585 ( .A1(n2424), .A2(n3005), .ZN(\mult_22/ab[44][7] ) );
  NOR2_X1 U10586 ( .A1(n2412), .A2(n3022), .ZN(\mult_22/ab[47][5] ) );
  NOR2_X1 U10587 ( .A1(n2510), .A2(n2869), .ZN(\mult_22/ab[22][21] ) );
  NOR2_X1 U10588 ( .A1(n2497), .A2(n2886), .ZN(\mult_22/ab[25][19] ) );
  NOR2_X1 U10589 ( .A1(n2461), .A2(n2940), .ZN(\mult_22/ab[34][13] ) );
  NOR2_X1 U10590 ( .A1(n2448), .A2(n2958), .ZN(\mult_22/ab[37][11] ) );
  NOR2_X1 U10591 ( .A1(n2436), .A2(n2981), .ZN(\mult_22/ab[40][9] ) );
  NOR2_X1 U10592 ( .A1(n2424), .A2(n2999), .ZN(\mult_22/ab[43][7] ) );
  NOR2_X1 U10593 ( .A1(n2412), .A2(n3016), .ZN(\mult_22/ab[46][5] ) );
  NOR2_X1 U10594 ( .A1(n2566), .A2(n2774), .ZN(\mult_22/ab[6][31] ) );
  NOR2_X1 U10595 ( .A1(n2498), .A2(n2880), .ZN(\mult_22/ab[24][19] ) );
  NOR2_X1 U10596 ( .A1(n2485), .A2(n2898), .ZN(\mult_22/ab[27][17] ) );
  NOR2_X1 U10597 ( .A1(n2461), .A2(n2934), .ZN(\mult_22/ab[33][13] ) );
  NOR2_X1 U10598 ( .A1(n2448), .A2(n2952), .ZN(\mult_22/ab[36][11] ) );
  NOR2_X1 U10599 ( .A1(n2436), .A2(n2975), .ZN(\mult_22/ab[39][9] ) );
  NOR2_X1 U10600 ( .A1(n2424), .A2(n2993), .ZN(\mult_22/ab[42][7] ) );
  NOR2_X1 U10601 ( .A1(n2412), .A2(n3010), .ZN(\mult_22/ab[45][5] ) );
  NOR2_X1 U10602 ( .A1(n2485), .A2(n2892), .ZN(\mult_22/ab[26][17] ) );
  NOR2_X1 U10603 ( .A1(n2473), .A2(n2910), .ZN(\mult_22/ab[29][15] ) );
  NOR2_X1 U10604 ( .A1(n2461), .A2(n2928), .ZN(\mult_22/ab[32][13] ) );
  NOR2_X1 U10605 ( .A1(n2449), .A2(n2946), .ZN(\mult_22/ab[35][11] ) );
  NOR2_X1 U10606 ( .A1(n2436), .A2(n2969), .ZN(\mult_22/ab[38][9] ) );
  NOR2_X1 U10607 ( .A1(n2424), .A2(n2987), .ZN(\mult_22/ab[41][7] ) );
  NOR2_X1 U10608 ( .A1(n2412), .A2(n3004), .ZN(\mult_22/ab[44][5] ) );
  NOR2_X1 U10609 ( .A1(n2473), .A2(n2904), .ZN(\mult_22/ab[28][15] ) );
  NOR2_X1 U10610 ( .A1(n2461), .A2(n2922), .ZN(\mult_22/ab[31][13] ) );
  NOR2_X1 U10611 ( .A1(n2449), .A2(n2940), .ZN(\mult_22/ab[34][11] ) );
  NOR2_X1 U10612 ( .A1(n2436), .A2(n2963), .ZN(\mult_22/ab[37][9] ) );
  NOR2_X1 U10613 ( .A1(n2424), .A2(n2981), .ZN(\mult_22/ab[40][7] ) );
  NOR2_X1 U10614 ( .A1(n2412), .A2(n2998), .ZN(\mult_22/ab[43][5] ) );
  NOR2_X1 U10615 ( .A1(n2461), .A2(n2916), .ZN(\mult_22/ab[30][13] ) );
  NOR2_X1 U10616 ( .A1(n2449), .A2(n2934), .ZN(\mult_22/ab[33][11] ) );
  NOR2_X1 U10617 ( .A1(n2436), .A2(n2957), .ZN(\mult_22/ab[36][9] ) );
  NOR2_X1 U10618 ( .A1(n2424), .A2(n2975), .ZN(\mult_22/ab[39][7] ) );
  NOR2_X1 U10619 ( .A1(n2412), .A2(n2992), .ZN(\mult_22/ab[42][5] ) );
  NOR2_X1 U10620 ( .A1(n2449), .A2(n2928), .ZN(\mult_22/ab[32][11] ) );
  NOR2_X1 U10621 ( .A1(n2437), .A2(n2951), .ZN(\mult_22/ab[35][9] ) );
  NOR2_X1 U10622 ( .A1(n2424), .A2(n2969), .ZN(\mult_22/ab[38][7] ) );
  NOR2_X1 U10623 ( .A1(n2412), .A2(n2986), .ZN(\mult_22/ab[41][5] ) );
  NOR2_X1 U10624 ( .A1(n2437), .A2(n2945), .ZN(\mult_22/ab[34][9] ) );
  NOR2_X1 U10625 ( .A1(n2424), .A2(n2963), .ZN(\mult_22/ab[37][7] ) );
  NOR2_X1 U10626 ( .A1(n2412), .A2(n2980), .ZN(\mult_22/ab[40][5] ) );
  NOR2_X1 U10627 ( .A1(n2424), .A2(n2957), .ZN(\mult_22/ab[36][7] ) );
  NOR2_X1 U10628 ( .A1(n2412), .A2(n2974), .ZN(\mult_22/ab[39][5] ) );
  NOR2_X1 U10629 ( .A1(n2412), .A2(n2968), .ZN(\mult_22/ab[38][5] ) );
  NOR2_X1 U10630 ( .A1(n2560), .A2(n2785), .ZN(\mult_22/ab[8][30] ) );
  NOR2_X1 U10631 ( .A1(n2399), .A2(n3038), .ZN(\mult_22/ab[50][3] ) );
  NOR2_X1 U10632 ( .A1(n2399), .A2(n3032), .ZN(\mult_22/ab[49][3] ) );
  NOR2_X1 U10633 ( .A1(n2399), .A2(n3026), .ZN(\mult_22/ab[48][3] ) );
  NOR2_X1 U10634 ( .A1(n2399), .A2(n3020), .ZN(\mult_22/ab[47][3] ) );
  NOR2_X1 U10635 ( .A1(n2400), .A2(n3014), .ZN(\mult_22/ab[46][3] ) );
  NOR2_X1 U10636 ( .A1(n2400), .A2(n3008), .ZN(\mult_22/ab[45][3] ) );
  NOR2_X1 U10637 ( .A1(n2400), .A2(n3002), .ZN(\mult_22/ab[44][3] ) );
  NOR2_X1 U10638 ( .A1(n2400), .A2(n2996), .ZN(\mult_22/ab[43][3] ) );
  NOR2_X1 U10639 ( .A1(n2400), .A2(n2990), .ZN(\mult_22/ab[42][3] ) );
  NOR2_X1 U10640 ( .A1(n2574), .A2(n2756), .ZN(\mult_22/ab[3][32] ) );
  NOR2_X1 U10641 ( .A1(n2400), .A2(n2984), .ZN(\mult_22/ab[41][3] ) );
  NOR2_X1 U10642 ( .A1(n2400), .A2(n2978), .ZN(\mult_22/ab[40][3] ) );
  NOR2_X1 U10643 ( .A1(n2552), .A2(n2815), .ZN(\mult_22/ab[13][28] ) );
  NOR2_X1 U10644 ( .A1(n2540), .A2(n2833), .ZN(\mult_22/ab[16][26] ) );
  NOR2_X1 U10645 ( .A1(n2524), .A2(n2845), .ZN(\mult_22/ab[18][24] ) );
  NOR2_X1 U10646 ( .A1(n2516), .A2(n2857), .ZN(\mult_22/ab[20][22] ) );
  NOR2_X1 U10647 ( .A1(n2504), .A2(n2869), .ZN(\mult_22/ab[22][20] ) );
  NOR2_X1 U10648 ( .A1(n2492), .A2(n2880), .ZN(\mult_22/ab[24][18] ) );
  NOR2_X1 U10649 ( .A1(n2479), .A2(n2892), .ZN(\mult_22/ab[26][16] ) );
  NOR2_X1 U10650 ( .A1(n2467), .A2(n2904), .ZN(\mult_22/ab[28][14] ) );
  NOR2_X1 U10651 ( .A1(n2455), .A2(n2916), .ZN(\mult_22/ab[30][12] ) );
  NOR2_X1 U10652 ( .A1(n2441), .A2(n2928), .ZN(\mult_22/ab[32][10] ) );
  NOR2_X1 U10653 ( .A1(n2431), .A2(n2945), .ZN(\mult_22/ab[34][8] ) );
  NOR2_X1 U10654 ( .A1(n2418), .A2(n2957), .ZN(\mult_22/ab[36][6] ) );
  NOR2_X1 U10655 ( .A1(n2560), .A2(n2779), .ZN(\mult_22/ab[7][30] ) );
  NOR2_X1 U10656 ( .A1(n2406), .A2(n2967), .ZN(\mult_22/ab[38][4] ) );
  NOR2_X1 U10657 ( .A1(n2560), .A2(n2773), .ZN(\mult_22/ab[6][30] ) );
  NOR2_X1 U10658 ( .A1(n2552), .A2(n2809), .ZN(\mult_22/ab[12][28] ) );
  NOR2_X1 U10659 ( .A1(n2400), .A2(n2972), .ZN(\mult_22/ab[39][3] ) );
  NOR2_X1 U10660 ( .A1(n2567), .A2(n2762), .ZN(\mult_22/ab[4][31] ) );
  NOR2_X1 U10661 ( .A1(n2546), .A2(n2821), .ZN(\mult_22/ab[14][27] ) );
  NOR2_X1 U10662 ( .A1(n2534), .A2(n2833), .ZN(\mult_22/ab[16][25] ) );
  NOR2_X1 U10663 ( .A1(n2522), .A2(n2845), .ZN(\mult_22/ab[18][23] ) );
  NOR2_X1 U10664 ( .A1(n2510), .A2(n2857), .ZN(\mult_22/ab[20][21] ) );
  NOR2_X1 U10665 ( .A1(n2498), .A2(n2868), .ZN(\mult_22/ab[22][19] ) );
  NOR2_X1 U10666 ( .A1(n2486), .A2(n2880), .ZN(\mult_22/ab[24][17] ) );
  NOR2_X1 U10667 ( .A1(n2473), .A2(n2892), .ZN(\mult_22/ab[26][15] ) );
  NOR2_X1 U10668 ( .A1(n2461), .A2(n2904), .ZN(\mult_22/ab[28][13] ) );
  NOR2_X1 U10669 ( .A1(n2449), .A2(n2916), .ZN(\mult_22/ab[30][11] ) );
  NOR2_X1 U10670 ( .A1(n2437), .A2(n2933), .ZN(\mult_22/ab[32][9] ) );
  NOR2_X1 U10671 ( .A1(n2425), .A2(n2945), .ZN(\mult_22/ab[34][7] ) );
  NOR2_X1 U10672 ( .A1(n2413), .A2(n2956), .ZN(\mult_22/ab[36][5] ) );
  NOR2_X1 U10673 ( .A1(n2553), .A2(n2803), .ZN(\mult_22/ab[11][28] ) );
  NOR2_X1 U10674 ( .A1(n2400), .A2(n2966), .ZN(\mult_22/ab[38][3] ) );
  NOR2_X1 U10675 ( .A1(n2553), .A2(n2797), .ZN(\mult_22/ab[10][28] ) );
  NOR2_X1 U10676 ( .A1(n2393), .A2(n3049), .ZN(\mult_22/ab[52][2] ) );
  NOR2_X1 U10677 ( .A1(n2393), .A2(n3043), .ZN(\mult_22/ab[51][2] ) );
  NOR2_X1 U10678 ( .A1(n2393), .A2(n3037), .ZN(\mult_22/ab[50][2] ) );
  NOR2_X1 U10679 ( .A1(n2393), .A2(n3031), .ZN(\mult_22/ab[49][2] ) );
  NOR2_X1 U10680 ( .A1(n2393), .A2(n3025), .ZN(\mult_22/ab[48][2] ) );
  NOR2_X1 U10681 ( .A1(n2393), .A2(n3019), .ZN(\mult_22/ab[47][2] ) );
  NOR2_X1 U10682 ( .A1(n2394), .A2(n3013), .ZN(\mult_22/ab[46][2] ) );
  NOR2_X1 U10683 ( .A1(n2394), .A2(n3007), .ZN(\mult_22/ab[45][2] ) );
  NOR2_X1 U10684 ( .A1(n2394), .A2(n3001), .ZN(\mult_22/ab[44][2] ) );
  NOR2_X1 U10685 ( .A1(n2394), .A2(n2995), .ZN(\mult_22/ab[43][2] ) );
  NOR2_X1 U10686 ( .A1(n2540), .A2(n2821), .ZN(\mult_22/ab[14][26] ) );
  NOR2_X1 U10687 ( .A1(n2524), .A2(n2833), .ZN(\mult_22/ab[16][24] ) );
  NOR2_X1 U10688 ( .A1(n2516), .A2(n2845), .ZN(\mult_22/ab[18][22] ) );
  NOR2_X1 U10689 ( .A1(n2504), .A2(n2857), .ZN(\mult_22/ab[20][20] ) );
  NOR2_X1 U10690 ( .A1(n2492), .A2(n2868), .ZN(\mult_22/ab[22][18] ) );
  NOR2_X1 U10691 ( .A1(n2480), .A2(n2880), .ZN(\mult_22/ab[24][16] ) );
  NOR2_X1 U10692 ( .A1(n2467), .A2(n2892), .ZN(\mult_22/ab[26][14] ) );
  NOR2_X1 U10693 ( .A1(n2461), .A2(n2898), .ZN(\mult_22/ab[27][13] ) );
  NOR2_X1 U10694 ( .A1(n2449), .A2(n2910), .ZN(\mult_22/ab[29][11] ) );
  NOR2_X1 U10695 ( .A1(n2437), .A2(n2927), .ZN(\mult_22/ab[31][9] ) );
  NOR2_X1 U10696 ( .A1(n2425), .A2(n2939), .ZN(\mult_22/ab[33][7] ) );
  NOR2_X1 U10697 ( .A1(n2413), .A2(n2950), .ZN(\mult_22/ab[35][5] ) );
  NOR2_X1 U10698 ( .A1(n2394), .A2(n2989), .ZN(\mult_22/ab[42][2] ) );
  NOR2_X1 U10699 ( .A1(n2394), .A2(n2983), .ZN(\mult_22/ab[41][2] ) );
  NOR2_X1 U10700 ( .A1(n2547), .A2(n2809), .ZN(\mult_22/ab[12][27] ) );
  NOR2_X1 U10701 ( .A1(n2534), .A2(n2821), .ZN(\mult_22/ab[14][25] ) );
  NOR2_X1 U10702 ( .A1(n2522), .A2(n2833), .ZN(\mult_22/ab[16][23] ) );
  NOR2_X1 U10703 ( .A1(n2510), .A2(n2845), .ZN(\mult_22/ab[18][21] ) );
  NOR2_X1 U10704 ( .A1(n2498), .A2(n2856), .ZN(\mult_22/ab[20][19] ) );
  NOR2_X1 U10705 ( .A1(n2486), .A2(n2868), .ZN(\mult_22/ab[22][17] ) );
  NOR2_X1 U10706 ( .A1(n2474), .A2(n2880), .ZN(\mult_22/ab[24][15] ) );
  NOR2_X1 U10707 ( .A1(n2461), .A2(n2892), .ZN(\mult_22/ab[26][13] ) );
  NOR2_X1 U10708 ( .A1(n2449), .A2(n2904), .ZN(\mult_22/ab[28][11] ) );
  NOR2_X1 U10709 ( .A1(n2437), .A2(n2921), .ZN(\mult_22/ab[30][9] ) );
  NOR2_X1 U10710 ( .A1(n2425), .A2(n2933), .ZN(\mult_22/ab[32][7] ) );
  NOR2_X1 U10711 ( .A1(n2413), .A2(n2944), .ZN(\mult_22/ab[34][5] ) );
  NOR2_X1 U10712 ( .A1(n2560), .A2(n2767), .ZN(\mult_22/ab[5][30] ) );
  NOR2_X1 U10713 ( .A1(n2400), .A2(n2960), .ZN(\mult_22/ab[37][3] ) );
  NOR2_X1 U10714 ( .A1(n2561), .A2(n2761), .ZN(\mult_22/ab[4][30] ) );
  NOR2_X1 U10715 ( .A1(n2548), .A2(n2791), .ZN(\mult_22/ab[9][28] ) );
  NOR2_X1 U10716 ( .A1(n2400), .A2(n2954), .ZN(\mult_22/ab[36][3] ) );
  NOR2_X1 U10717 ( .A1(n2541), .A2(n2809), .ZN(\mult_22/ab[12][26] ) );
  NOR2_X1 U10718 ( .A1(n2524), .A2(n2821), .ZN(\mult_22/ab[14][24] ) );
  NOR2_X1 U10719 ( .A1(n2516), .A2(n2833), .ZN(\mult_22/ab[16][22] ) );
  NOR2_X1 U10720 ( .A1(n2504), .A2(n2845), .ZN(\mult_22/ab[18][20] ) );
  NOR2_X1 U10721 ( .A1(n2492), .A2(n2856), .ZN(\mult_22/ab[20][18] ) );
  NOR2_X1 U10722 ( .A1(n2480), .A2(n2868), .ZN(\mult_22/ab[22][16] ) );
  NOR2_X1 U10723 ( .A1(n2548), .A2(n2785), .ZN(\mult_22/ab[8][28] ) );
  NOR2_X1 U10724 ( .A1(n2468), .A2(n2880), .ZN(\mult_22/ab[24][14] ) );
  NOR2_X1 U10725 ( .A1(n2394), .A2(n2977), .ZN(\mult_22/ab[40][2] ) );
  NOR2_X1 U10726 ( .A1(n2455), .A2(n2892), .ZN(\mult_22/ab[26][12] ) );
  NOR2_X1 U10727 ( .A1(n2441), .A2(n2904), .ZN(\mult_22/ab[28][10] ) );
  NOR2_X1 U10728 ( .A1(n2431), .A2(n2921), .ZN(\mult_22/ab[30][8] ) );
  NOR2_X1 U10729 ( .A1(n2419), .A2(n2933), .ZN(\mult_22/ab[32][6] ) );
  NOR2_X1 U10730 ( .A1(n2406), .A2(n2943), .ZN(\mult_22/ab[34][4] ) );
  NOR2_X1 U10731 ( .A1(n2547), .A2(n2797), .ZN(\mult_22/ab[10][27] ) );
  NOR2_X1 U10732 ( .A1(n2535), .A2(n2809), .ZN(\mult_22/ab[12][25] ) );
  NOR2_X1 U10733 ( .A1(n2522), .A2(n2821), .ZN(\mult_22/ab[14][23] ) );
  NOR2_X1 U10734 ( .A1(n2510), .A2(n2833), .ZN(\mult_22/ab[16][21] ) );
  NOR2_X1 U10735 ( .A1(n2498), .A2(n2844), .ZN(\mult_22/ab[18][19] ) );
  NOR2_X1 U10736 ( .A1(n2486), .A2(n2856), .ZN(\mult_22/ab[20][17] ) );
  NOR2_X1 U10737 ( .A1(n2474), .A2(n2868), .ZN(\mult_22/ab[22][15] ) );
  NOR2_X1 U10738 ( .A1(n2462), .A2(n2880), .ZN(\mult_22/ab[24][13] ) );
  NOR2_X1 U10739 ( .A1(n2449), .A2(n2892), .ZN(\mult_22/ab[26][11] ) );
  NOR2_X1 U10740 ( .A1(n2437), .A2(n2909), .ZN(\mult_22/ab[28][9] ) );
  NOR2_X1 U10741 ( .A1(n2425), .A2(n2921), .ZN(\mult_22/ab[30][7] ) );
  NOR2_X1 U10742 ( .A1(n2413), .A2(n2932), .ZN(\mult_22/ab[32][5] ) );
  NOR2_X1 U10743 ( .A1(n2401), .A2(n2948), .ZN(\mult_22/ab[35][3] ) );
  NOR2_X1 U10744 ( .A1(n2394), .A2(n2971), .ZN(\mult_22/ab[39][2] ) );
  NOR2_X1 U10745 ( .A1(n2541), .A2(n2797), .ZN(\mult_22/ab[10][26] ) );
  NOR2_X1 U10746 ( .A1(n2524), .A2(n2809), .ZN(\mult_22/ab[12][24] ) );
  NOR2_X1 U10747 ( .A1(n2516), .A2(n2821), .ZN(\mult_22/ab[14][22] ) );
  NOR2_X1 U10748 ( .A1(n2504), .A2(n2833), .ZN(\mult_22/ab[16][20] ) );
  NOR2_X1 U10749 ( .A1(n2492), .A2(n2844), .ZN(\mult_22/ab[18][18] ) );
  NOR2_X1 U10750 ( .A1(n2480), .A2(n2856), .ZN(\mult_22/ab[20][16] ) );
  NOR2_X1 U10751 ( .A1(n2562), .A2(n2755), .ZN(\mult_22/ab[3][30] ) );
  NOR2_X1 U10752 ( .A1(n2468), .A2(n2868), .ZN(\mult_22/ab[22][14] ) );
  NOR2_X1 U10753 ( .A1(n2401), .A2(n2942), .ZN(\mult_22/ab[34][3] ) );
  NOR2_X1 U10754 ( .A1(n2456), .A2(n2880), .ZN(\mult_22/ab[24][12] ) );
  NOR2_X1 U10755 ( .A1(n2441), .A2(n2892), .ZN(\mult_22/ab[26][10] ) );
  NOR2_X1 U10756 ( .A1(n2431), .A2(n2909), .ZN(\mult_22/ab[28][8] ) );
  NOR2_X1 U10757 ( .A1(n2419), .A2(n2921), .ZN(\mult_22/ab[30][6] ) );
  NOR2_X1 U10758 ( .A1(n2548), .A2(n2779), .ZN(\mult_22/ab[7][28] ) );
  NOR2_X1 U10759 ( .A1(n2387), .A2(n3060), .ZN(\mult_22/ab[54][1] ) );
  NOR2_X1 U10760 ( .A1(n2387), .A2(n3054), .ZN(\mult_22/ab[53][1] ) );
  NOR2_X1 U10761 ( .A1(n2387), .A2(n3048), .ZN(\mult_22/ab[52][1] ) );
  NOR2_X1 U10762 ( .A1(n2387), .A2(n3042), .ZN(\mult_22/ab[51][1] ) );
  NOR2_X1 U10763 ( .A1(n2387), .A2(n3036), .ZN(\mult_22/ab[50][1] ) );
  NOR2_X1 U10764 ( .A1(n2387), .A2(n3030), .ZN(\mult_22/ab[49][1] ) );
  NOR2_X1 U10765 ( .A1(n2387), .A2(n3024), .ZN(\mult_22/ab[48][1] ) );
  NOR2_X1 U10766 ( .A1(n2388), .A2(n3018), .ZN(\mult_22/ab[47][1] ) );
  NOR2_X1 U10767 ( .A1(n2388), .A2(n3012), .ZN(\mult_22/ab[46][1] ) );
  NOR2_X1 U10768 ( .A1(n2388), .A2(n3006), .ZN(\mult_22/ab[45][1] ) );
  NOR2_X1 U10769 ( .A1(n2388), .A2(n3000), .ZN(\mult_22/ab[44][1] ) );
  NOR2_X1 U10770 ( .A1(n2405), .A2(n2931), .ZN(\mult_22/ab[32][4] ) );
  NOR2_X1 U10771 ( .A1(n2394), .A2(n2965), .ZN(\mult_22/ab[38][2] ) );
  NOR2_X1 U10772 ( .A1(n2388), .A2(n2994), .ZN(\mult_22/ab[43][1] ) );
  NOR2_X1 U10773 ( .A1(n2388), .A2(n2988), .ZN(\mult_22/ab[42][1] ) );
  NOR2_X1 U10774 ( .A1(n2548), .A2(n2773), .ZN(\mult_22/ab[6][28] ) );
  NOR2_X1 U10775 ( .A1(n2394), .A2(n2959), .ZN(\mult_22/ab[37][2] ) );
  NOR2_X1 U10776 ( .A1(n2401), .A2(n2936), .ZN(\mult_22/ab[33][3] ) );
  NOR2_X1 U10777 ( .A1(n2388), .A2(n2982), .ZN(\mult_22/ab[41][1] ) );
  NOR2_X1 U10778 ( .A1(n2394), .A2(n2953), .ZN(\mult_22/ab[36][2] ) );
  NOR2_X1 U10779 ( .A1(n2395), .A2(n2947), .ZN(\mult_22/ab[35][2] ) );
  NOR2_X1 U10780 ( .A1(n2395), .A2(n2941), .ZN(\mult_22/ab[34][2] ) );
  NOR2_X1 U10781 ( .A1(n2384), .A2(n3084), .ZN(\mult_22/ab[58][0] ) );
  NOR2_X1 U10782 ( .A1(n2384), .A2(n3078), .ZN(\mult_22/ab[57][0] ) );
  NOR2_X1 U10783 ( .A1(n2384), .A2(n3072), .ZN(\mult_22/ab[56][0] ) );
  NOR2_X1 U10784 ( .A1(n2586), .A2(n2888), .ZN(\mult_22/ab[25][34] ) );
  NOR2_X1 U10785 ( .A1(n2692), .A2(n2757), .ZN(\mult_22/ab[3][52] ) );
  INV_X1 U10786 ( .A(\mult_22/CARRYB[2][56] ), .ZN(n740) );
  INV_X1 U10787 ( .A(\mult_22/SUMB[2][57] ), .ZN(n741) );
  INV_X1 U10788 ( .A(\mult_22/SUMB[24][36] ), .ZN(n701) );
  NOR2_X1 U10789 ( .A1(n2464), .A2(n3114), .ZN(\mult_22/ab[63][14] ) );
  NOR2_X1 U10790 ( .A1(n2518), .A2(n3115), .ZN(\mult_22/ab[63][23] ) );
  NOR2_X1 U10791 ( .A1(n2476), .A2(n3114), .ZN(\mult_22/ab[63][16] ) );
  NOR2_X1 U10792 ( .A1(n2528), .A2(n3115), .ZN(\mult_22/ab[63][24] ) );
  NOR2_X1 U10793 ( .A1(n2470), .A2(n3114), .ZN(\mult_22/ab[63][15] ) );
  NOR2_X1 U10794 ( .A1(n2536), .A2(n3115), .ZN(\mult_22/ab[63][26] ) );
  NOR2_X1 U10795 ( .A1(n2482), .A2(n3114), .ZN(\mult_22/ab[63][17] ) );
  NOR2_X1 U10796 ( .A1(n2488), .A2(n3114), .ZN(\mult_22/ab[63][18] ) );
  NOR2_X1 U10797 ( .A1(n2530), .A2(n3115), .ZN(\mult_22/ab[63][25] ) );
  NOR2_X1 U10798 ( .A1(n2512), .A2(n3115), .ZN(\mult_22/ab[63][22] ) );
  NOR2_X1 U10799 ( .A1(n2506), .A2(n3115), .ZN(\mult_22/ab[63][21] ) );
  NOR2_X1 U10800 ( .A1(n2458), .A2(n3114), .ZN(\mult_22/ab[63][13] ) );
  NOR2_X1 U10801 ( .A1(n2500), .A2(n3115), .ZN(\mult_22/ab[63][20] ) );
  NOR2_X1 U10802 ( .A1(n2494), .A2(n3114), .ZN(\mult_22/ab[63][19] ) );
  NOR2_X1 U10803 ( .A1(n2452), .A2(n3114), .ZN(\mult_22/ab[63][12] ) );
  NOR2_X1 U10804 ( .A1(n2446), .A2(n3114), .ZN(\mult_22/ab[63][11] ) );
  NOR2_X1 U10805 ( .A1(n2548), .A2(n3115), .ZN(\mult_22/ab[63][28] ) );
  NOR2_X1 U10806 ( .A1(n2542), .A2(n3115), .ZN(\mult_22/ab[63][27] ) );
  NOR2_X1 U10807 ( .A1(n2748), .A2(n2800), .ZN(\mult_22/ab[10][63] ) );
  NOR2_X1 U10808 ( .A1(n2745), .A2(n2806), .ZN(\mult_22/ab[11][62] ) );
  NOR2_X1 U10809 ( .A1(n2745), .A2(n2812), .ZN(\mult_22/ab[12][62] ) );
  NOR2_X1 U10810 ( .A1(n2753), .A2(n2806), .ZN(\mult_22/ab[11][63] ) );
  NOR2_X1 U10811 ( .A1(n2753), .A2(n2812), .ZN(\mult_22/ab[12][63] ) );
  NOR2_X1 U10812 ( .A1(n2186), .A2(n2818), .ZN(\mult_22/ab[13][62] ) );
  NOR2_X1 U10813 ( .A1(n2185), .A2(n2824), .ZN(\mult_22/ab[14][62] ) );
  NOR2_X1 U10814 ( .A1(n2752), .A2(n2818), .ZN(\mult_22/ab[13][63] ) );
  NOR2_X1 U10815 ( .A1(n2744), .A2(n2830), .ZN(\mult_22/ab[15][62] ) );
  NOR2_X1 U10816 ( .A1(n2752), .A2(n2824), .ZN(\mult_22/ab[14][63] ) );
  NOR2_X1 U10817 ( .A1(n2745), .A2(n2836), .ZN(\mult_22/ab[16][62] ) );
  NOR2_X1 U10818 ( .A1(n2752), .A2(n2830), .ZN(\mult_22/ab[15][63] ) );
  NOR2_X1 U10819 ( .A1(n2746), .A2(n2842), .ZN(\mult_22/ab[17][62] ) );
  NOR2_X1 U10820 ( .A1(n2752), .A2(n2836), .ZN(\mult_22/ab[16][63] ) );
  NOR2_X1 U10821 ( .A1(n2752), .A2(n2842), .ZN(\mult_22/ab[17][63] ) );
  NOR2_X1 U10822 ( .A1(n2747), .A2(n2848), .ZN(\mult_22/ab[18][62] ) );
  NOR2_X1 U10823 ( .A1(n2752), .A2(n2860), .ZN(\mult_22/ab[20][63] ) );
  NOR2_X1 U10824 ( .A1(n2744), .A2(n2866), .ZN(\mult_22/ab[21][62] ) );
  NOR2_X1 U10825 ( .A1(n2744), .A2(n2860), .ZN(\mult_22/ab[20][62] ) );
  NOR2_X1 U10826 ( .A1(n2752), .A2(n2854), .ZN(\mult_22/ab[19][63] ) );
  NOR2_X1 U10827 ( .A1(n2743), .A2(n2854), .ZN(\mult_22/ab[19][62] ) );
  NOR2_X1 U10828 ( .A1(n2752), .A2(n2848), .ZN(\mult_22/ab[18][63] ) );
  NOR2_X1 U10829 ( .A1(n2745), .A2(n2896), .ZN(\mult_22/ab[26][62] ) );
  NOR2_X1 U10830 ( .A1(n2751), .A2(n2890), .ZN(\mult_22/ab[25][63] ) );
  NOR2_X1 U10831 ( .A1(n2746), .A2(n2902), .ZN(\mult_22/ab[27][62] ) );
  NOR2_X1 U10832 ( .A1(n2751), .A2(n2896), .ZN(\mult_22/ab[26][63] ) );
  NOR2_X1 U10833 ( .A1(n2751), .A2(n2902), .ZN(\mult_22/ab[27][63] ) );
  NOR2_X1 U10834 ( .A1(n2747), .A2(n2908), .ZN(\mult_22/ab[28][62] ) );
  NOR2_X1 U10835 ( .A1(n2743), .A2(n2914), .ZN(\mult_22/ab[29][62] ) );
  NOR2_X1 U10836 ( .A1(n2751), .A2(n2908), .ZN(\mult_22/ab[28][63] ) );
  NOR2_X1 U10837 ( .A1(n2744), .A2(n2872), .ZN(\mult_22/ab[22][62] ) );
  NOR2_X1 U10838 ( .A1(n2752), .A2(n2866), .ZN(\mult_22/ab[21][63] ) );
  NOR2_X1 U10839 ( .A1(n2752), .A2(n2872), .ZN(\mult_22/ab[22][63] ) );
  NOR2_X1 U10840 ( .A1(n2186), .A2(n2878), .ZN(\mult_22/ab[23][62] ) );
  NOR2_X1 U10841 ( .A1(n2752), .A2(n2878), .ZN(\mult_22/ab[23][63] ) );
  NOR2_X1 U10842 ( .A1(n2185), .A2(n2884), .ZN(\mult_22/ab[24][62] ) );
  NOR2_X1 U10843 ( .A1(n2744), .A2(n2890), .ZN(\mult_22/ab[25][62] ) );
  NOR2_X1 U10844 ( .A1(n2752), .A2(n2884), .ZN(\mult_22/ab[24][63] ) );
  NOR2_X1 U10845 ( .A1(n2458), .A2(n3108), .ZN(\mult_22/ab[62][13] ) );
  NOR2_X1 U10846 ( .A1(n2452), .A2(n3108), .ZN(\mult_22/ab[62][12] ) );
  NOR2_X1 U10847 ( .A1(n2458), .A2(n3102), .ZN(\mult_22/ab[61][13] ) );
  NOR2_X1 U10848 ( .A1(n2464), .A2(n3108), .ZN(\mult_22/ab[62][14] ) );
  NOR2_X1 U10849 ( .A1(n2506), .A2(n3109), .ZN(\mult_22/ab[62][21] ) );
  NOR2_X1 U10850 ( .A1(n2464), .A2(n3102), .ZN(\mult_22/ab[61][14] ) );
  NOR2_X1 U10851 ( .A1(n2500), .A2(n3109), .ZN(\mult_22/ab[62][20] ) );
  NOR2_X1 U10852 ( .A1(n2464), .A2(n3096), .ZN(\mult_22/ab[60][14] ) );
  NOR2_X1 U10853 ( .A1(n2548), .A2(n3109), .ZN(\mult_22/ab[62][28] ) );
  NOR2_X1 U10854 ( .A1(n2470), .A2(n3108), .ZN(\mult_22/ab[62][15] ) );
  NOR2_X1 U10855 ( .A1(n2512), .A2(n3109), .ZN(\mult_22/ab[62][22] ) );
  NOR2_X1 U10856 ( .A1(n2476), .A2(n3108), .ZN(\mult_22/ab[62][16] ) );
  NOR2_X1 U10857 ( .A1(n2470), .A2(n3102), .ZN(\mult_22/ab[61][15] ) );
  NOR2_X1 U10858 ( .A1(n2554), .A2(n3109), .ZN(\mult_22/ab[62][29] ) );
  NOR2_X1 U10859 ( .A1(n2506), .A2(n3103), .ZN(\mult_22/ab[61][21] ) );
  NOR2_X1 U10860 ( .A1(n2542), .A2(n3109), .ZN(\mult_22/ab[62][27] ) );
  NOR2_X1 U10861 ( .A1(n2470), .A2(n3096), .ZN(\mult_22/ab[60][15] ) );
  NOR2_X1 U10862 ( .A1(n2512), .A2(n3103), .ZN(\mult_22/ab[61][22] ) );
  NOR2_X1 U10863 ( .A1(n2482), .A2(n3108), .ZN(\mult_22/ab[62][17] ) );
  NOR2_X1 U10864 ( .A1(n2476), .A2(n3102), .ZN(\mult_22/ab[61][16] ) );
  NOR2_X1 U10865 ( .A1(n2470), .A2(n3090), .ZN(\mult_22/ab[59][15] ) );
  NOR2_X1 U10866 ( .A1(n2494), .A2(n3108), .ZN(\mult_22/ab[62][19] ) );
  NOR2_X1 U10867 ( .A1(n2500), .A2(n3103), .ZN(\mult_22/ab[61][20] ) );
  NOR2_X1 U10868 ( .A1(n2482), .A2(n3102), .ZN(\mult_22/ab[61][17] ) );
  NOR2_X1 U10869 ( .A1(n2476), .A2(n3096), .ZN(\mult_22/ab[60][16] ) );
  NOR2_X1 U10870 ( .A1(n2554), .A2(n3103), .ZN(\mult_22/ab[61][29] ) );
  NOR2_X1 U10871 ( .A1(n2548), .A2(n3103), .ZN(\mult_22/ab[61][28] ) );
  NOR2_X1 U10872 ( .A1(n2512), .A2(n3097), .ZN(\mult_22/ab[60][22] ) );
  NOR2_X1 U10873 ( .A1(n2476), .A2(n3090), .ZN(\mult_22/ab[59][16] ) );
  NOR2_X1 U10874 ( .A1(n2536), .A2(n3109), .ZN(\mult_22/ab[62][26] ) );
  NOR2_X1 U10875 ( .A1(n2506), .A2(n3097), .ZN(\mult_22/ab[60][21] ) );
  NOR2_X1 U10876 ( .A1(n2488), .A2(n3108), .ZN(\mult_22/ab[62][18] ) );
  NOR2_X1 U10877 ( .A1(n2482), .A2(n3096), .ZN(\mult_22/ab[60][17] ) );
  NOR2_X1 U10878 ( .A1(n2476), .A2(n3084), .ZN(\mult_22/ab[58][16] ) );
  NOR2_X1 U10879 ( .A1(n2542), .A2(n3103), .ZN(\mult_22/ab[61][27] ) );
  NOR2_X1 U10880 ( .A1(n2488), .A2(n3102), .ZN(\mult_22/ab[61][18] ) );
  NOR2_X1 U10881 ( .A1(n2560), .A2(n3103), .ZN(\mult_22/ab[61][30] ) );
  NOR2_X1 U10882 ( .A1(n2518), .A2(n3103), .ZN(\mult_22/ab[61][23] ) );
  NOR2_X1 U10883 ( .A1(n2518), .A2(n3097), .ZN(\mult_22/ab[60][23] ) );
  NOR2_X1 U10884 ( .A1(n2494), .A2(n3102), .ZN(\mult_22/ab[61][19] ) );
  NOR2_X1 U10885 ( .A1(n2482), .A2(n3090), .ZN(\mult_22/ab[59][17] ) );
  NOR2_X1 U10886 ( .A1(n2488), .A2(n3096), .ZN(\mult_22/ab[60][18] ) );
  NOR2_X1 U10887 ( .A1(n2512), .A2(n3091), .ZN(\mult_22/ab[59][22] ) );
  NOR2_X1 U10888 ( .A1(n2500), .A2(n3097), .ZN(\mult_22/ab[60][20] ) );
  NOR2_X1 U10889 ( .A1(n2554), .A2(n3097), .ZN(\mult_22/ab[60][29] ) );
  NOR2_X1 U10890 ( .A1(n2482), .A2(n3084), .ZN(\mult_22/ab[58][17] ) );
  NOR2_X1 U10891 ( .A1(n2518), .A2(n3091), .ZN(\mult_22/ab[59][23] ) );
  NOR2_X1 U10892 ( .A1(n2548), .A2(n3097), .ZN(\mult_22/ab[60][28] ) );
  NOR2_X1 U10893 ( .A1(n2488), .A2(n3090), .ZN(\mult_22/ab[59][18] ) );
  NOR2_X1 U10894 ( .A1(n2483), .A2(n3078), .ZN(\mult_22/ab[57][17] ) );
  NOR2_X1 U10895 ( .A1(n2506), .A2(n3091), .ZN(\mult_22/ab[59][21] ) );
  NOR2_X1 U10896 ( .A1(n2518), .A2(n3109), .ZN(\mult_22/ab[62][23] ) );
  NOR2_X1 U10897 ( .A1(n2560), .A2(n3097), .ZN(\mult_22/ab[60][30] ) );
  NOR2_X1 U10898 ( .A1(n2494), .A2(n3096), .ZN(\mult_22/ab[60][19] ) );
  NOR2_X1 U10899 ( .A1(n2488), .A2(n3084), .ZN(\mult_22/ab[58][18] ) );
  NOR2_X1 U10900 ( .A1(n2494), .A2(n3090), .ZN(\mult_22/ab[59][19] ) );
  NOR2_X1 U10901 ( .A1(n2518), .A2(n3085), .ZN(\mult_22/ab[58][23] ) );
  NOR2_X1 U10902 ( .A1(n2500), .A2(n3091), .ZN(\mult_22/ab[59][20] ) );
  NOR2_X1 U10903 ( .A1(n2536), .A2(n3103), .ZN(\mult_22/ab[61][26] ) );
  NOR2_X1 U10904 ( .A1(n2512), .A2(n3085), .ZN(\mult_22/ab[58][22] ) );
  NOR2_X1 U10905 ( .A1(n2489), .A2(n3078), .ZN(\mult_22/ab[57][18] ) );
  NOR2_X1 U10906 ( .A1(n2542), .A2(n3097), .ZN(\mult_22/ab[60][27] ) );
  NOR2_X1 U10907 ( .A1(n2528), .A2(n3091), .ZN(\mult_22/ab[59][24] ) );
  NOR2_X1 U10908 ( .A1(n2554), .A2(n3091), .ZN(\mult_22/ab[59][29] ) );
  NOR2_X1 U10909 ( .A1(n2489), .A2(n3072), .ZN(\mult_22/ab[56][18] ) );
  NOR2_X1 U10910 ( .A1(n2494), .A2(n3084), .ZN(\mult_22/ab[58][19] ) );
  NOR2_X1 U10911 ( .A1(n2560), .A2(n3091), .ZN(\mult_22/ab[59][30] ) );
  NOR2_X1 U10912 ( .A1(n2566), .A2(n3098), .ZN(\mult_22/ab[60][31] ) );
  NOR2_X1 U10913 ( .A1(n2528), .A2(n3085), .ZN(\mult_22/ab[58][24] ) );
  NOR2_X1 U10914 ( .A1(n2528), .A2(n3097), .ZN(\mult_22/ab[60][24] ) );
  NOR2_X1 U10915 ( .A1(n2506), .A2(n3085), .ZN(\mult_22/ab[58][21] ) );
  NOR2_X1 U10916 ( .A1(n2530), .A2(n3109), .ZN(\mult_22/ab[62][25] ) );
  NOR2_X1 U10917 ( .A1(n2548), .A2(n3091), .ZN(\mult_22/ab[59][28] ) );
  NOR2_X1 U10918 ( .A1(n2495), .A2(n3078), .ZN(\mult_22/ab[57][19] ) );
  NOR2_X1 U10919 ( .A1(n2500), .A2(n3085), .ZN(\mult_22/ab[58][20] ) );
  NOR2_X1 U10920 ( .A1(n2519), .A2(n3079), .ZN(\mult_22/ab[57][23] ) );
  NOR2_X1 U10921 ( .A1(n2495), .A2(n3072), .ZN(\mult_22/ab[56][19] ) );
  NOR2_X1 U10922 ( .A1(n2528), .A2(n3079), .ZN(\mult_22/ab[57][24] ) );
  NOR2_X1 U10923 ( .A1(n2513), .A2(n3079), .ZN(\mult_22/ab[57][22] ) );
  NOR2_X1 U10924 ( .A1(n2566), .A2(n3092), .ZN(\mult_22/ab[59][31] ) );
  NOR2_X1 U10925 ( .A1(n2495), .A2(n3066), .ZN(\mult_22/ab[55][19] ) );
  NOR2_X1 U10926 ( .A1(n2501), .A2(n3079), .ZN(\mult_22/ab[57][20] ) );
  NOR2_X1 U10927 ( .A1(n2507), .A2(n3079), .ZN(\mult_22/ab[57][21] ) );
  NOR2_X1 U10928 ( .A1(n2560), .A2(n3085), .ZN(\mult_22/ab[58][30] ) );
  NOR2_X1 U10929 ( .A1(n2554), .A2(n3085), .ZN(\mult_22/ab[58][29] ) );
  NOR2_X1 U10930 ( .A1(n2501), .A2(n3073), .ZN(\mult_22/ab[56][20] ) );
  NOR2_X1 U10931 ( .A1(n2528), .A2(n3073), .ZN(\mult_22/ab[56][24] ) );
  NOR2_X1 U10932 ( .A1(n2519), .A2(n3073), .ZN(\mult_22/ab[56][23] ) );
  NOR2_X1 U10933 ( .A1(n2528), .A2(n3103), .ZN(\mult_22/ab[61][24] ) );
  NOR2_X1 U10934 ( .A1(n2530), .A2(n3085), .ZN(\mult_22/ab[58][25] ) );
  NOR2_X1 U10935 ( .A1(n2531), .A2(n3079), .ZN(\mult_22/ab[57][25] ) );
  NOR2_X1 U10936 ( .A1(n2542), .A2(n3091), .ZN(\mult_22/ab[59][27] ) );
  NOR2_X1 U10937 ( .A1(n2567), .A2(n3086), .ZN(\mult_22/ab[58][31] ) );
  NOR2_X1 U10938 ( .A1(n2501), .A2(n3067), .ZN(\mult_22/ab[55][20] ) );
  NOR2_X1 U10939 ( .A1(n2513), .A2(n3073), .ZN(\mult_22/ab[56][22] ) );
  NOR2_X1 U10940 ( .A1(n2536), .A2(n3097), .ZN(\mult_22/ab[60][26] ) );
  NOR2_X1 U10941 ( .A1(n2507), .A2(n3073), .ZN(\mult_22/ab[56][21] ) );
  NOR2_X1 U10942 ( .A1(n2501), .A2(n3061), .ZN(\mult_22/ab[54][20] ) );
  NOR2_X1 U10943 ( .A1(n2531), .A2(n3073), .ZN(\mult_22/ab[56][25] ) );
  NOR2_X1 U10944 ( .A1(n2530), .A2(n3091), .ZN(\mult_22/ab[59][25] ) );
  NOR2_X1 U10945 ( .A1(n2548), .A2(n3085), .ZN(\mult_22/ab[58][28] ) );
  NOR2_X1 U10946 ( .A1(n2528), .A2(n3067), .ZN(\mult_22/ab[55][24] ) );
  NOR2_X1 U10947 ( .A1(n2576), .A2(n3092), .ZN(\mult_22/ab[59][32] ) );
  NOR2_X1 U10948 ( .A1(n2507), .A2(n3067), .ZN(\mult_22/ab[55][21] ) );
  NOR2_X1 U10949 ( .A1(n2519), .A2(n3067), .ZN(\mult_22/ab[55][23] ) );
  NOR2_X1 U10950 ( .A1(n2561), .A2(n3079), .ZN(\mult_22/ab[57][30] ) );
  NOR2_X1 U10951 ( .A1(n2513), .A2(n3067), .ZN(\mult_22/ab[55][22] ) );
  NOR2_X1 U10952 ( .A1(n2531), .A2(n3067), .ZN(\mult_22/ab[55][25] ) );
  NOR2_X1 U10953 ( .A1(n2567), .A2(n3080), .ZN(\mult_22/ab[57][31] ) );
  NOR2_X1 U10954 ( .A1(n2507), .A2(n3061), .ZN(\mult_22/ab[54][21] ) );
  NOR2_X1 U10955 ( .A1(n2576), .A2(n3086), .ZN(\mult_22/ab[58][32] ) );
  NOR2_X1 U10956 ( .A1(n2555), .A2(n3079), .ZN(\mult_22/ab[57][29] ) );
  NOR2_X1 U10957 ( .A1(n2530), .A2(n3103), .ZN(\mult_22/ab[61][25] ) );
  NOR2_X1 U10958 ( .A1(n2507), .A2(n3055), .ZN(\mult_22/ab[53][21] ) );
  NOR2_X1 U10959 ( .A1(n2530), .A2(n3097), .ZN(\mult_22/ab[60][25] ) );
  NOR2_X1 U10960 ( .A1(n2527), .A2(n3061), .ZN(\mult_22/ab[54][24] ) );
  NOR2_X1 U10961 ( .A1(n2513), .A2(n3061), .ZN(\mult_22/ab[54][22] ) );
  NOR2_X1 U10962 ( .A1(n2531), .A2(n3061), .ZN(\mult_22/ab[54][25] ) );
  NOR2_X1 U10963 ( .A1(n2519), .A2(n3061), .ZN(\mult_22/ab[54][23] ) );
  NOR2_X1 U10964 ( .A1(n2537), .A2(n3073), .ZN(\mult_22/ab[56][26] ) );
  NOR2_X1 U10965 ( .A1(n2576), .A2(n3080), .ZN(\mult_22/ab[57][32] ) );
  NOR2_X1 U10966 ( .A1(n2536), .A2(n3091), .ZN(\mult_22/ab[59][26] ) );
  NOR2_X1 U10967 ( .A1(n2537), .A2(n3079), .ZN(\mult_22/ab[57][26] ) );
  NOR2_X1 U10968 ( .A1(n2537), .A2(n3067), .ZN(\mult_22/ab[55][26] ) );
  NOR2_X1 U10969 ( .A1(n2542), .A2(n3085), .ZN(\mult_22/ab[58][27] ) );
  NOR2_X1 U10970 ( .A1(n2513), .A2(n3055), .ZN(\mult_22/ab[53][22] ) );
  NOR2_X1 U10971 ( .A1(n2567), .A2(n3074), .ZN(\mult_22/ab[56][31] ) );
  NOR2_X1 U10972 ( .A1(n2536), .A2(n3085), .ZN(\mult_22/ab[58][26] ) );
  NOR2_X1 U10973 ( .A1(n2561), .A2(n3073), .ZN(\mult_22/ab[56][30] ) );
  NOR2_X1 U10974 ( .A1(n2549), .A2(n3079), .ZN(\mult_22/ab[57][28] ) );
  NOR2_X1 U10975 ( .A1(n2537), .A2(n3061), .ZN(\mult_22/ab[54][26] ) );
  NOR2_X1 U10976 ( .A1(n2519), .A2(n3055), .ZN(\mult_22/ab[53][23] ) );
  NOR2_X1 U10977 ( .A1(n2527), .A2(n3055), .ZN(\mult_22/ab[53][24] ) );
  NOR2_X1 U10978 ( .A1(n2513), .A2(n3049), .ZN(\mult_22/ab[52][22] ) );
  NOR2_X1 U10979 ( .A1(n2531), .A2(n3055), .ZN(\mult_22/ab[53][25] ) );
  NOR2_X1 U10980 ( .A1(n2576), .A2(n3074), .ZN(\mult_22/ab[56][32] ) );
  NOR2_X1 U10981 ( .A1(n2555), .A2(n3073), .ZN(\mult_22/ab[56][29] ) );
  NOR2_X1 U10982 ( .A1(n2537), .A2(n3055), .ZN(\mult_22/ab[53][26] ) );
  NOR2_X1 U10983 ( .A1(n2519), .A2(n3049), .ZN(\mult_22/ab[52][23] ) );
  NOR2_X1 U10984 ( .A1(n2578), .A2(n3086), .ZN(\mult_22/ab[58][33] ) );
  NOR2_X1 U10985 ( .A1(n2527), .A2(n3049), .ZN(\mult_22/ab[52][24] ) );
  NOR2_X1 U10986 ( .A1(n2543), .A2(n3079), .ZN(\mult_22/ab[57][27] ) );
  NOR2_X1 U10987 ( .A1(n2531), .A2(n3049), .ZN(\mult_22/ab[52][25] ) );
  NOR2_X1 U10988 ( .A1(n2578), .A2(n3080), .ZN(\mult_22/ab[57][33] ) );
  NOR2_X1 U10989 ( .A1(n2567), .A2(n3068), .ZN(\mult_22/ab[55][31] ) );
  NOR2_X1 U10990 ( .A1(n2543), .A2(n3067), .ZN(\mult_22/ab[55][27] ) );
  NOR2_X1 U10991 ( .A1(n2519), .A2(n3043), .ZN(\mult_22/ab[51][23] ) );
  NOR2_X1 U10992 ( .A1(n2543), .A2(n3073), .ZN(\mult_22/ab[56][27] ) );
  NOR2_X1 U10993 ( .A1(n2537), .A2(n3049), .ZN(\mult_22/ab[52][26] ) );
  NOR2_X1 U10994 ( .A1(n2543), .A2(n3061), .ZN(\mult_22/ab[54][27] ) );
  NOR2_X1 U10995 ( .A1(n2575), .A2(n3068), .ZN(\mult_22/ab[55][32] ) );
  NOR2_X1 U10996 ( .A1(n2561), .A2(n3067), .ZN(\mult_22/ab[55][30] ) );
  NOR2_X1 U10997 ( .A1(n2578), .A2(n3074), .ZN(\mult_22/ab[56][33] ) );
  NOR2_X1 U10998 ( .A1(n2549), .A2(n3073), .ZN(\mult_22/ab[56][28] ) );
  NOR2_X1 U10999 ( .A1(n2543), .A2(n3055), .ZN(\mult_22/ab[53][27] ) );
  NOR2_X1 U11000 ( .A1(n2527), .A2(n3043), .ZN(\mult_22/ab[51][24] ) );
  NOR2_X1 U11001 ( .A1(n2531), .A2(n3043), .ZN(\mult_22/ab[51][25] ) );
  NOR2_X1 U11002 ( .A1(n2543), .A2(n3049), .ZN(\mult_22/ab[52][27] ) );
  NOR2_X1 U11003 ( .A1(n2537), .A2(n3043), .ZN(\mult_22/ab[51][26] ) );
  NOR2_X1 U11004 ( .A1(n2578), .A2(n3068), .ZN(\mult_22/ab[55][33] ) );
  NOR2_X1 U11005 ( .A1(n2527), .A2(n3037), .ZN(\mult_22/ab[50][24] ) );
  NOR2_X1 U11006 ( .A1(n2555), .A2(n3067), .ZN(\mult_22/ab[55][29] ) );
  NOR2_X1 U11007 ( .A1(n2549), .A2(n3067), .ZN(\mult_22/ab[55][28] ) );
  NOR2_X1 U11008 ( .A1(n2543), .A2(n3043), .ZN(\mult_22/ab[51][27] ) );
  NOR2_X1 U11009 ( .A1(n2567), .A2(n3062), .ZN(\mult_22/ab[54][31] ) );
  NOR2_X1 U11010 ( .A1(n2575), .A2(n3062), .ZN(\mult_22/ab[54][32] ) );
  NOR2_X1 U11011 ( .A1(n2531), .A2(n3037), .ZN(\mult_22/ab[50][25] ) );
  NOR2_X1 U11012 ( .A1(n2537), .A2(n3037), .ZN(\mult_22/ab[50][26] ) );
  NOR2_X1 U11013 ( .A1(n2549), .A2(n3061), .ZN(\mult_22/ab[54][28] ) );
  NOR2_X1 U11014 ( .A1(n2528), .A2(n3109), .ZN(\mult_22/ab[62][24] ) );
  NOR2_X1 U11015 ( .A1(n2561), .A2(n3061), .ZN(\mult_22/ab[54][30] ) );
  NOR2_X1 U11016 ( .A1(n2549), .A2(n3055), .ZN(\mult_22/ab[53][28] ) );
  NOR2_X1 U11017 ( .A1(n2578), .A2(n3062), .ZN(\mult_22/ab[54][33] ) );
  NOR2_X1 U11018 ( .A1(n2543), .A2(n3037), .ZN(\mult_22/ab[50][27] ) );
  NOR2_X1 U11019 ( .A1(n2531), .A2(n3031), .ZN(\mult_22/ab[49][25] ) );
  NOR2_X1 U11020 ( .A1(n2549), .A2(n3049), .ZN(\mult_22/ab[52][28] ) );
  NOR2_X1 U11021 ( .A1(n2584), .A2(n3080), .ZN(\mult_22/ab[57][34] ) );
  NOR2_X1 U11022 ( .A1(n2584), .A2(n3074), .ZN(\mult_22/ab[56][34] ) );
  NOR2_X1 U11023 ( .A1(n2555), .A2(n3061), .ZN(\mult_22/ab[54][29] ) );
  NOR2_X1 U11024 ( .A1(n2537), .A2(n3031), .ZN(\mult_22/ab[49][26] ) );
  NOR2_X1 U11025 ( .A1(n2549), .A2(n3043), .ZN(\mult_22/ab[51][28] ) );
  NOR2_X1 U11026 ( .A1(n2584), .A2(n3068), .ZN(\mult_22/ab[55][34] ) );
  NOR2_X1 U11027 ( .A1(n2543), .A2(n3031), .ZN(\mult_22/ab[49][27] ) );
  NOR2_X1 U11028 ( .A1(n2575), .A2(n3056), .ZN(\mult_22/ab[53][32] ) );
  NOR2_X1 U11029 ( .A1(n2555), .A2(n2761), .ZN(\mult_22/ab[4][29] ) );
  NOR2_X1 U11030 ( .A1(n2536), .A2(n2791), .ZN(\mult_22/ab[9][26] ) );
  NOR2_X1 U11031 ( .A1(n2524), .A2(n2803), .ZN(\mult_22/ab[11][24] ) );
  NOR2_X1 U11032 ( .A1(n2516), .A2(n2815), .ZN(\mult_22/ab[13][22] ) );
  NOR2_X1 U11033 ( .A1(n2504), .A2(n2827), .ZN(\mult_22/ab[15][20] ) );
  NOR2_X1 U11034 ( .A1(n2492), .A2(n2838), .ZN(\mult_22/ab[17][18] ) );
  NOR2_X1 U11035 ( .A1(n2480), .A2(n2850), .ZN(\mult_22/ab[19][16] ) );
  NOR2_X1 U11036 ( .A1(n2468), .A2(n2862), .ZN(\mult_22/ab[21][14] ) );
  NOR2_X1 U11037 ( .A1(n2456), .A2(n2874), .ZN(\mult_22/ab[23][12] ) );
  NOR2_X1 U11038 ( .A1(n2441), .A2(n2886), .ZN(\mult_22/ab[25][10] ) );
  NOR2_X1 U11039 ( .A1(n2431), .A2(n2903), .ZN(\mult_22/ab[27][8] ) );
  NOR2_X1 U11040 ( .A1(n2419), .A2(n2915), .ZN(\mult_22/ab[29][6] ) );
  NOR2_X1 U11041 ( .A1(n2405), .A2(n2925), .ZN(\mult_22/ab[31][4] ) );
  NOR2_X1 U11042 ( .A1(n2556), .A2(n2755), .ZN(\mult_22/ab[3][29] ) );
  NOR2_X1 U11043 ( .A1(n2542), .A2(n2779), .ZN(\mult_22/ab[7][27] ) );
  NOR2_X1 U11044 ( .A1(n2530), .A2(n2791), .ZN(\mult_22/ab[9][25] ) );
  NOR2_X1 U11045 ( .A1(n2523), .A2(n2803), .ZN(\mult_22/ab[11][23] ) );
  NOR2_X1 U11046 ( .A1(n2510), .A2(n2815), .ZN(\mult_22/ab[13][21] ) );
  NOR2_X1 U11047 ( .A1(n2498), .A2(n2826), .ZN(\mult_22/ab[15][19] ) );
  NOR2_X1 U11048 ( .A1(n2486), .A2(n2838), .ZN(\mult_22/ab[17][17] ) );
  NOR2_X1 U11049 ( .A1(n2474), .A2(n2850), .ZN(\mult_22/ab[19][15] ) );
  NOR2_X1 U11050 ( .A1(n2462), .A2(n2862), .ZN(\mult_22/ab[21][13] ) );
  NOR2_X1 U11051 ( .A1(n2450), .A2(n2874), .ZN(\mult_22/ab[23][11] ) );
  NOR2_X1 U11052 ( .A1(n2437), .A2(n2891), .ZN(\mult_22/ab[25][9] ) );
  NOR2_X1 U11053 ( .A1(n2425), .A2(n2903), .ZN(\mult_22/ab[27][7] ) );
  NOR2_X1 U11054 ( .A1(n2413), .A2(n2914), .ZN(\mult_22/ab[29][5] ) );
  NOR2_X1 U11055 ( .A1(n2549), .A2(n3037), .ZN(\mult_22/ab[50][28] ) );
  NOR2_X1 U11056 ( .A1(n2536), .A2(n2779), .ZN(\mult_22/ab[7][26] ) );
  NOR2_X1 U11057 ( .A1(n2529), .A2(n2791), .ZN(\mult_22/ab[9][24] ) );
  NOR2_X1 U11058 ( .A1(n2517), .A2(n2803), .ZN(\mult_22/ab[11][22] ) );
  NOR2_X1 U11059 ( .A1(n2504), .A2(n2815), .ZN(\mult_22/ab[13][20] ) );
  NOR2_X1 U11060 ( .A1(n2492), .A2(n2826), .ZN(\mult_22/ab[15][18] ) );
  NOR2_X1 U11061 ( .A1(n2480), .A2(n2838), .ZN(\mult_22/ab[17][16] ) );
  NOR2_X1 U11062 ( .A1(n2468), .A2(n2850), .ZN(\mult_22/ab[19][14] ) );
  NOR2_X1 U11063 ( .A1(n2456), .A2(n2862), .ZN(\mult_22/ab[21][12] ) );
  NOR2_X1 U11064 ( .A1(n2441), .A2(n2874), .ZN(\mult_22/ab[23][10] ) );
  NOR2_X1 U11065 ( .A1(n2431), .A2(n2891), .ZN(\mult_22/ab[25][8] ) );
  NOR2_X1 U11066 ( .A1(n2419), .A2(n2903), .ZN(\mult_22/ab[27][6] ) );
  NOR2_X1 U11067 ( .A1(n2405), .A2(n2913), .ZN(\mult_22/ab[29][4] ) );
  NOR2_X1 U11068 ( .A1(n2542), .A2(n2767), .ZN(\mult_22/ab[5][27] ) );
  NOR2_X1 U11069 ( .A1(n2530), .A2(n2779), .ZN(\mult_22/ab[7][25] ) );
  NOR2_X1 U11070 ( .A1(n2518), .A2(n2791), .ZN(\mult_22/ab[9][23] ) );
  NOR2_X1 U11071 ( .A1(n2511), .A2(n2803), .ZN(\mult_22/ab[11][21] ) );
  NOR2_X1 U11072 ( .A1(n2498), .A2(n2814), .ZN(\mult_22/ab[13][19] ) );
  NOR2_X1 U11073 ( .A1(n2486), .A2(n2826), .ZN(\mult_22/ab[15][17] ) );
  NOR2_X1 U11074 ( .A1(n2474), .A2(n2838), .ZN(\mult_22/ab[17][15] ) );
  NOR2_X1 U11075 ( .A1(n2731), .A2(n2818), .ZN(\mult_22/ab[13][60] ) );
  NOR2_X1 U11076 ( .A1(n2462), .A2(n2850), .ZN(\mult_22/ab[19][13] ) );
  NOR2_X1 U11077 ( .A1(n2450), .A2(n2862), .ZN(\mult_22/ab[21][11] ) );
  NOR2_X1 U11078 ( .A1(n2438), .A2(n2879), .ZN(\mult_22/ab[23][9] ) );
  NOR2_X1 U11079 ( .A1(n2425), .A2(n2891), .ZN(\mult_22/ab[25][7] ) );
  NOR2_X1 U11080 ( .A1(n2413), .A2(n2902), .ZN(\mult_22/ab[27][5] ) );
  NOR2_X1 U11081 ( .A1(n2537), .A2(n3025), .ZN(\mult_22/ab[48][26] ) );
  NOR2_X1 U11082 ( .A1(n2737), .A2(n2812), .ZN(\mult_22/ab[12][61] ) );
  NOR2_X1 U11083 ( .A1(n2543), .A2(n3019), .ZN(\mult_22/ab[47][27] ) );
  NOR2_X1 U11084 ( .A1(n2536), .A2(n2767), .ZN(\mult_22/ab[5][26] ) );
  NOR2_X1 U11085 ( .A1(n2537), .A2(n2761), .ZN(\mult_22/ab[4][26] ) );
  NOR2_X1 U11086 ( .A1(n2528), .A2(n2779), .ZN(\mult_22/ab[7][24] ) );
  NOR2_X1 U11087 ( .A1(n2528), .A2(n2773), .ZN(\mult_22/ab[6][24] ) );
  NOR2_X1 U11088 ( .A1(n2512), .A2(n2791), .ZN(\mult_22/ab[9][22] ) );
  NOR2_X1 U11089 ( .A1(n2512), .A2(n2785), .ZN(\mult_22/ab[8][22] ) );
  NOR2_X1 U11090 ( .A1(n2505), .A2(n2803), .ZN(\mult_22/ab[11][20] ) );
  NOR2_X1 U11091 ( .A1(n2505), .A2(n2797), .ZN(\mult_22/ab[10][20] ) );
  NOR2_X1 U11092 ( .A1(n2492), .A2(n2814), .ZN(\mult_22/ab[13][18] ) );
  NOR2_X1 U11093 ( .A1(n2493), .A2(n2808), .ZN(\mult_22/ab[12][18] ) );
  NOR2_X1 U11094 ( .A1(n2480), .A2(n2826), .ZN(\mult_22/ab[15][16] ) );
  NOR2_X1 U11095 ( .A1(n2480), .A2(n2820), .ZN(\mult_22/ab[14][16] ) );
  NOR2_X1 U11096 ( .A1(n2468), .A2(n2838), .ZN(\mult_22/ab[17][14] ) );
  NOR2_X1 U11097 ( .A1(n2468), .A2(n2832), .ZN(\mult_22/ab[16][14] ) );
  NOR2_X1 U11098 ( .A1(n2456), .A2(n2850), .ZN(\mult_22/ab[19][12] ) );
  NOR2_X1 U11099 ( .A1(n2456), .A2(n2844), .ZN(\mult_22/ab[18][12] ) );
  NOR2_X1 U11100 ( .A1(n2440), .A2(n2862), .ZN(\mult_22/ab[21][10] ) );
  NOR2_X1 U11101 ( .A1(n2440), .A2(n2856), .ZN(\mult_22/ab[20][10] ) );
  NOR2_X1 U11102 ( .A1(n2432), .A2(n2879), .ZN(\mult_22/ab[23][8] ) );
  NOR2_X1 U11103 ( .A1(n2432), .A2(n2873), .ZN(\mult_22/ab[22][8] ) );
  NOR2_X1 U11104 ( .A1(n2419), .A2(n2890), .ZN(\mult_22/ab[25][6] ) );
  NOR2_X1 U11105 ( .A1(n2420), .A2(n2884), .ZN(\mult_22/ab[24][6] ) );
  NOR2_X1 U11106 ( .A1(n2405), .A2(n2901), .ZN(\mult_22/ab[27][4] ) );
  NOR2_X1 U11107 ( .A1(n2405), .A2(n2895), .ZN(\mult_22/ab[26][4] ) );
  NOR2_X1 U11108 ( .A1(n2567), .A2(n3056), .ZN(\mult_22/ab[53][31] ) );
  NOR2_X1 U11109 ( .A1(n2550), .A2(n3013), .ZN(\mult_22/ab[46][28] ) );
  NOR2_X1 U11110 ( .A1(n2538), .A2(n2755), .ZN(\mult_22/ab[3][26] ) );
  NOR2_X1 U11111 ( .A1(n2528), .A2(n2767), .ZN(\mult_22/ab[5][24] ) );
  NOR2_X1 U11112 ( .A1(n2512), .A2(n2779), .ZN(\mult_22/ab[7][22] ) );
  NOR2_X1 U11113 ( .A1(n2500), .A2(n2791), .ZN(\mult_22/ab[9][20] ) );
  NOR2_X1 U11114 ( .A1(n2493), .A2(n2802), .ZN(\mult_22/ab[11][18] ) );
  NOR2_X1 U11115 ( .A1(n2480), .A2(n2814), .ZN(\mult_22/ab[13][16] ) );
  NOR2_X1 U11116 ( .A1(n2468), .A2(n2826), .ZN(\mult_22/ab[15][14] ) );
  NOR2_X1 U11117 ( .A1(n2456), .A2(n2838), .ZN(\mult_22/ab[17][12] ) );
  NOR2_X1 U11118 ( .A1(n2440), .A2(n2850), .ZN(\mult_22/ab[19][10] ) );
  NOR2_X1 U11119 ( .A1(n2432), .A2(n2867), .ZN(\mult_22/ab[21][8] ) );
  NOR2_X1 U11120 ( .A1(n2420), .A2(n2878), .ZN(\mult_22/ab[23][6] ) );
  NOR2_X1 U11121 ( .A1(n2405), .A2(n2889), .ZN(\mult_22/ab[25][4] ) );
  NOR2_X1 U11122 ( .A1(n2556), .A2(n3007), .ZN(\mult_22/ab[45][29] ) );
  NOR2_X1 U11123 ( .A1(n2568), .A2(n2996), .ZN(\mult_22/ab[43][31] ) );
  NOR2_X1 U11124 ( .A1(n2579), .A2(n2984), .ZN(\mult_22/ab[41][33] ) );
  NOR2_X1 U11125 ( .A1(n2527), .A2(n2761), .ZN(\mult_22/ab[4][24] ) );
  NOR2_X1 U11126 ( .A1(n2512), .A2(n2773), .ZN(\mult_22/ab[6][22] ) );
  NOR2_X1 U11127 ( .A1(n2591), .A2(n2972), .ZN(\mult_22/ab[39][35] ) );
  NOR2_X1 U11128 ( .A1(n2500), .A2(n2785), .ZN(\mult_22/ab[8][20] ) );
  NOR2_X1 U11129 ( .A1(n2603), .A2(n2960), .ZN(\mult_22/ab[37][37] ) );
  NOR2_X1 U11130 ( .A1(n2493), .A2(n2796), .ZN(\mult_22/ab[10][18] ) );
  NOR2_X1 U11131 ( .A1(n2481), .A2(n2808), .ZN(\mult_22/ab[12][16] ) );
  NOR2_X1 U11132 ( .A1(n2468), .A2(n2820), .ZN(\mult_22/ab[14][14] ) );
  NOR2_X1 U11133 ( .A1(n2456), .A2(n2832), .ZN(\mult_22/ab[16][12] ) );
  NOR2_X1 U11134 ( .A1(n2440), .A2(n2844), .ZN(\mult_22/ab[18][10] ) );
  NOR2_X1 U11135 ( .A1(n2432), .A2(n2861), .ZN(\mult_22/ab[20][8] ) );
  NOR2_X1 U11136 ( .A1(n2420), .A2(n2872), .ZN(\mult_22/ab[22][6] ) );
  NOR2_X1 U11137 ( .A1(n2405), .A2(n2883), .ZN(\mult_22/ab[24][4] ) );
  NOR2_X1 U11138 ( .A1(n2562), .A2(n3001), .ZN(\mult_22/ab[44][30] ) );
  NOR2_X1 U11139 ( .A1(n2574), .A2(n2990), .ZN(\mult_22/ab[42][32] ) );
  NOR2_X1 U11140 ( .A1(n2585), .A2(n2978), .ZN(\mult_22/ab[40][34] ) );
  NOR2_X1 U11141 ( .A1(n2597), .A2(n2966), .ZN(\mult_22/ab[38][36] ) );
  NOR2_X1 U11142 ( .A1(n2609), .A2(n2954), .ZN(\mult_22/ab[36][38] ) );
  NOR2_X1 U11143 ( .A1(n2615), .A2(n2948), .ZN(\mult_22/ab[35][39] ) );
  NOR2_X1 U11144 ( .A1(n2626), .A2(n2936), .ZN(\mult_22/ab[33][41] ) );
  NOR2_X1 U11145 ( .A1(n2637), .A2(n2925), .ZN(\mult_22/ab[31][43] ) );
  NOR2_X1 U11146 ( .A1(n2649), .A2(n2913), .ZN(\mult_22/ab[29][45] ) );
  NOR2_X1 U11147 ( .A1(n2663), .A2(n2901), .ZN(\mult_22/ab[27][47] ) );
  NOR2_X1 U11148 ( .A1(n2673), .A2(n2889), .ZN(\mult_22/ab[25][49] ) );
  NOR2_X1 U11149 ( .A1(n2688), .A2(n2877), .ZN(\mult_22/ab[23][51] ) );
  NOR2_X1 U11150 ( .A1(n2700), .A2(n2865), .ZN(\mult_22/ab[21][53] ) );
  NOR2_X1 U11151 ( .A1(n2710), .A2(n2854), .ZN(\mult_22/ab[19][55] ) );
  NOR2_X1 U11152 ( .A1(n2716), .A2(n2842), .ZN(\mult_22/ab[17][57] ) );
  NOR2_X1 U11153 ( .A1(n2727), .A2(n2830), .ZN(\mult_22/ab[15][59] ) );
  NOR2_X1 U11154 ( .A1(n2543), .A2(n3025), .ZN(\mult_22/ab[48][27] ) );
  NOR2_X1 U11155 ( .A1(n2526), .A2(n2755), .ZN(\mult_22/ab[3][24] ) );
  NOR2_X1 U11156 ( .A1(n2512), .A2(n2767), .ZN(\mult_22/ab[5][22] ) );
  NOR2_X1 U11157 ( .A1(n2500), .A2(n2779), .ZN(\mult_22/ab[7][20] ) );
  NOR2_X1 U11158 ( .A1(n2488), .A2(n2790), .ZN(\mult_22/ab[9][18] ) );
  NOR2_X1 U11159 ( .A1(n2481), .A2(n2802), .ZN(\mult_22/ab[11][16] ) );
  NOR2_X1 U11160 ( .A1(n2468), .A2(n2814), .ZN(\mult_22/ab[13][14] ) );
  NOR2_X1 U11161 ( .A1(n2456), .A2(n2826), .ZN(\mult_22/ab[15][12] ) );
  NOR2_X1 U11162 ( .A1(n2440), .A2(n2838), .ZN(\mult_22/ab[17][10] ) );
  NOR2_X1 U11163 ( .A1(n2432), .A2(n2855), .ZN(\mult_22/ab[19][8] ) );
  NOR2_X1 U11164 ( .A1(n2420), .A2(n2866), .ZN(\mult_22/ab[21][6] ) );
  NOR2_X1 U11165 ( .A1(n2405), .A2(n2877), .ZN(\mult_22/ab[23][4] ) );
  NOR2_X1 U11166 ( .A1(n2621), .A2(n2942), .ZN(\mult_22/ab[34][40] ) );
  NOR2_X1 U11167 ( .A1(n2633), .A2(n2931), .ZN(\mult_22/ab[32][42] ) );
  NOR2_X1 U11168 ( .A1(n2645), .A2(n2919), .ZN(\mult_22/ab[30][44] ) );
  NOR2_X1 U11169 ( .A1(n2657), .A2(n2907), .ZN(\mult_22/ab[28][46] ) );
  NOR2_X1 U11170 ( .A1(n2669), .A2(n2895), .ZN(\mult_22/ab[26][48] ) );
  NOR2_X1 U11171 ( .A1(n2681), .A2(n2883), .ZN(\mult_22/ab[24][50] ) );
  NOR2_X1 U11172 ( .A1(n2691), .A2(n2871), .ZN(\mult_22/ab[22][52] ) );
  NOR2_X1 U11173 ( .A1(n2704), .A2(n2860), .ZN(\mult_22/ab[20][54] ) );
  NOR2_X1 U11174 ( .A1(n2719), .A2(n2836), .ZN(\mult_22/ab[16][58] ) );
  NOR2_X1 U11175 ( .A1(n2731), .A2(n2824), .ZN(\mult_22/ab[14][60] ) );
  NOR2_X1 U11176 ( .A1(n2740), .A2(n2818), .ZN(\mult_22/ab[13][61] ) );
  NOR2_X1 U11177 ( .A1(n2549), .A2(n3019), .ZN(\mult_22/ab[47][28] ) );
  NOR2_X1 U11178 ( .A1(n2562), .A2(n3007), .ZN(\mult_22/ab[45][30] ) );
  NOR2_X1 U11179 ( .A1(n2574), .A2(n2996), .ZN(\mult_22/ab[43][32] ) );
  NOR2_X1 U11180 ( .A1(n2585), .A2(n2984), .ZN(\mult_22/ab[41][34] ) );
  NOR2_X1 U11181 ( .A1(n2597), .A2(n2972), .ZN(\mult_22/ab[39][36] ) );
  NOR2_X1 U11182 ( .A1(n2556), .A2(n3013), .ZN(\mult_22/ab[46][29] ) );
  NOR2_X1 U11183 ( .A1(n2568), .A2(n3002), .ZN(\mult_22/ab[44][31] ) );
  NOR2_X1 U11184 ( .A1(n2579), .A2(n2990), .ZN(\mult_22/ab[42][33] ) );
  NOR2_X1 U11185 ( .A1(n2591), .A2(n2978), .ZN(\mult_22/ab[40][35] ) );
  NOR2_X1 U11186 ( .A1(n2603), .A2(n2966), .ZN(\mult_22/ab[38][37] ) );
  NOR2_X1 U11187 ( .A1(n2513), .A2(n2761), .ZN(\mult_22/ab[4][22] ) );
  NOR2_X1 U11188 ( .A1(n2500), .A2(n2773), .ZN(\mult_22/ab[6][20] ) );
  NOR2_X1 U11189 ( .A1(n2488), .A2(n2784), .ZN(\mult_22/ab[8][18] ) );
  NOR2_X1 U11190 ( .A1(n2481), .A2(n2796), .ZN(\mult_22/ab[10][16] ) );
  NOR2_X1 U11191 ( .A1(n2469), .A2(n2808), .ZN(\mult_22/ab[12][14] ) );
  NOR2_X1 U11192 ( .A1(n2456), .A2(n2820), .ZN(\mult_22/ab[14][12] ) );
  NOR2_X1 U11193 ( .A1(n2440), .A2(n2832), .ZN(\mult_22/ab[16][10] ) );
  NOR2_X1 U11194 ( .A1(n2432), .A2(n2849), .ZN(\mult_22/ab[18][8] ) );
  NOR2_X1 U11195 ( .A1(n2420), .A2(n2861), .ZN(\mult_22/ab[20][6] ) );
  NOR2_X1 U11196 ( .A1(n2405), .A2(n2871), .ZN(\mult_22/ab[22][4] ) );
  NOR2_X1 U11197 ( .A1(n2609), .A2(n2960), .ZN(\mult_22/ab[37][38] ) );
  NOR2_X1 U11198 ( .A1(n2578), .A2(n3056), .ZN(\mult_22/ab[53][33] ) );
  NOR2_X1 U11199 ( .A1(n2614), .A2(n2954), .ZN(\mult_22/ab[36][39] ) );
  NOR2_X1 U11200 ( .A1(n2626), .A2(n2942), .ZN(\mult_22/ab[34][41] ) );
  NOR2_X1 U11201 ( .A1(n2637), .A2(n2931), .ZN(\mult_22/ab[32][43] ) );
  NOR2_X1 U11202 ( .A1(n2649), .A2(n2919), .ZN(\mult_22/ab[30][45] ) );
  NOR2_X1 U11203 ( .A1(n2663), .A2(n2907), .ZN(\mult_22/ab[28][47] ) );
  NOR2_X1 U11204 ( .A1(n2673), .A2(n2895), .ZN(\mult_22/ab[26][49] ) );
  NOR2_X1 U11205 ( .A1(n2688), .A2(n2883), .ZN(\mult_22/ab[24][51] ) );
  NOR2_X1 U11206 ( .A1(n2699), .A2(n2871), .ZN(\mult_22/ab[22][53] ) );
  NOR2_X1 U11207 ( .A1(n2710), .A2(n2860), .ZN(\mult_22/ab[20][55] ) );
  NOR2_X1 U11208 ( .A1(n2716), .A2(n2848), .ZN(\mult_22/ab[18][57] ) );
  NOR2_X1 U11209 ( .A1(n2728), .A2(n2836), .ZN(\mult_22/ab[16][59] ) );
  NOR2_X1 U11210 ( .A1(n2621), .A2(n2948), .ZN(\mult_22/ab[35][40] ) );
  NOR2_X1 U11211 ( .A1(n2633), .A2(n2936), .ZN(\mult_22/ab[33][42] ) );
  NOR2_X1 U11212 ( .A1(n2645), .A2(n2925), .ZN(\mult_22/ab[31][44] ) );
  NOR2_X1 U11213 ( .A1(n2657), .A2(n2913), .ZN(\mult_22/ab[29][46] ) );
  NOR2_X1 U11214 ( .A1(n2669), .A2(n2901), .ZN(\mult_22/ab[27][48] ) );
  NOR2_X1 U11215 ( .A1(n2681), .A2(n2889), .ZN(\mult_22/ab[25][50] ) );
  NOR2_X1 U11216 ( .A1(n2691), .A2(n2877), .ZN(\mult_22/ab[23][52] ) );
  NOR2_X1 U11217 ( .A1(n2704), .A2(n2866), .ZN(\mult_22/ab[21][54] ) );
  NOR2_X1 U11218 ( .A1(n2719), .A2(n2842), .ZN(\mult_22/ab[17][58] ) );
  NOR2_X1 U11219 ( .A1(n2507), .A2(n2761), .ZN(\mult_22/ab[4][21] ) );
  NOR2_X1 U11220 ( .A1(n2494), .A2(n2772), .ZN(\mult_22/ab[6][19] ) );
  NOR2_X1 U11221 ( .A1(n2482), .A2(n2784), .ZN(\mult_22/ab[8][17] ) );
  NOR2_X1 U11222 ( .A1(n2475), .A2(n2796), .ZN(\mult_22/ab[10][15] ) );
  NOR2_X1 U11223 ( .A1(n2508), .A2(n2755), .ZN(\mult_22/ab[3][21] ) );
  NOR2_X1 U11224 ( .A1(n2494), .A2(n2766), .ZN(\mult_22/ab[5][19] ) );
  NOR2_X1 U11225 ( .A1(n2482), .A2(n2778), .ZN(\mult_22/ab[7][17] ) );
  NOR2_X1 U11226 ( .A1(n2470), .A2(n2790), .ZN(\mult_22/ab[9][15] ) );
  NOR2_X1 U11227 ( .A1(n2463), .A2(n2808), .ZN(\mult_22/ab[12][13] ) );
  NOR2_X1 U11228 ( .A1(n2450), .A2(n2820), .ZN(\mult_22/ab[14][11] ) );
  NOR2_X1 U11229 ( .A1(n2438), .A2(n2837), .ZN(\mult_22/ab[16][9] ) );
  NOR2_X1 U11230 ( .A1(n2426), .A2(n2849), .ZN(\mult_22/ab[18][7] ) );
  NOR2_X1 U11231 ( .A1(n2414), .A2(n2860), .ZN(\mult_22/ab[20][5] ) );
  NOR2_X1 U11232 ( .A1(n2463), .A2(n2802), .ZN(\mult_22/ab[11][13] ) );
  NOR2_X1 U11233 ( .A1(n2450), .A2(n2814), .ZN(\mult_22/ab[13][11] ) );
  NOR2_X1 U11234 ( .A1(n2438), .A2(n2831), .ZN(\mult_22/ab[15][9] ) );
  NOR2_X1 U11235 ( .A1(n2426), .A2(n2843), .ZN(\mult_22/ab[17][7] ) );
  NOR2_X1 U11236 ( .A1(n2414), .A2(n2854), .ZN(\mult_22/ab[19][5] ) );
  NOR2_X1 U11237 ( .A1(n2731), .A2(n2830), .ZN(\mult_22/ab[15][60] ) );
  NOR2_X1 U11238 ( .A1(n2741), .A2(n2824), .ZN(\mult_22/ab[14][61] ) );
  NOR2_X1 U11239 ( .A1(n2502), .A2(n2755), .ZN(\mult_22/ab[3][20] ) );
  NOR2_X1 U11240 ( .A1(n2488), .A2(n2766), .ZN(\mult_22/ab[5][18] ) );
  NOR2_X1 U11241 ( .A1(n2476), .A2(n2778), .ZN(\mult_22/ab[7][16] ) );
  NOR2_X1 U11242 ( .A1(n2464), .A2(n2790), .ZN(\mult_22/ab[9][14] ) );
  NOR2_X1 U11243 ( .A1(n2457), .A2(n2802), .ZN(\mult_22/ab[11][12] ) );
  NOR2_X1 U11244 ( .A1(n2440), .A2(n2814), .ZN(\mult_22/ab[13][10] ) );
  NOR2_X1 U11245 ( .A1(n2432), .A2(n2831), .ZN(\mult_22/ab[15][8] ) );
  NOR2_X1 U11246 ( .A1(n2420), .A2(n2843), .ZN(\mult_22/ab[17][6] ) );
  NOR2_X1 U11247 ( .A1(n2404), .A2(n2853), .ZN(\mult_22/ab[19][4] ) );
  NOR2_X1 U11248 ( .A1(n2549), .A2(n3031), .ZN(\mult_22/ab[49][28] ) );
  NOR2_X1 U11249 ( .A1(n2549), .A2(n3025), .ZN(\mult_22/ab[48][28] ) );
  NOR2_X1 U11250 ( .A1(n2496), .A2(n2754), .ZN(\mult_22/ab[3][19] ) );
  NOR2_X1 U11251 ( .A1(n2482), .A2(n2766), .ZN(\mult_22/ab[5][17] ) );
  NOR2_X1 U11252 ( .A1(n2470), .A2(n2778), .ZN(\mult_22/ab[7][15] ) );
  NOR2_X1 U11253 ( .A1(n2458), .A2(n2790), .ZN(\mult_22/ab[9][13] ) );
  NOR2_X1 U11254 ( .A1(n2451), .A2(n2802), .ZN(\mult_22/ab[11][11] ) );
  NOR2_X1 U11255 ( .A1(n2438), .A2(n2819), .ZN(\mult_22/ab[13][9] ) );
  NOR2_X1 U11256 ( .A1(n2426), .A2(n2831), .ZN(\mult_22/ab[15][7] ) );
  NOR2_X1 U11257 ( .A1(n2414), .A2(n2842), .ZN(\mult_22/ab[17][5] ) );
  NOR2_X1 U11258 ( .A1(n2562), .A2(n3013), .ZN(\mult_22/ab[46][30] ) );
  NOR2_X1 U11259 ( .A1(n2574), .A2(n3002), .ZN(\mult_22/ab[44][32] ) );
  NOR2_X1 U11260 ( .A1(n2585), .A2(n2990), .ZN(\mult_22/ab[42][34] ) );
  NOR2_X1 U11261 ( .A1(n2555), .A2(n3019), .ZN(\mult_22/ab[47][29] ) );
  NOR2_X1 U11262 ( .A1(n2568), .A2(n3008), .ZN(\mult_22/ab[45][31] ) );
  NOR2_X1 U11263 ( .A1(n2579), .A2(n2996), .ZN(\mult_22/ab[43][33] ) );
  NOR2_X1 U11264 ( .A1(n2597), .A2(n2978), .ZN(\mult_22/ab[40][36] ) );
  NOR2_X1 U11265 ( .A1(n2609), .A2(n2966), .ZN(\mult_22/ab[38][38] ) );
  NOR2_X1 U11266 ( .A1(n2591), .A2(n2984), .ZN(\mult_22/ab[41][35] ) );
  NOR2_X1 U11267 ( .A1(n2603), .A2(n2972), .ZN(\mult_22/ab[39][37] ) );
  NOR2_X1 U11268 ( .A1(n2490), .A2(n2754), .ZN(\mult_22/ab[3][18] ) );
  NOR2_X1 U11269 ( .A1(n2476), .A2(n2766), .ZN(\mult_22/ab[5][16] ) );
  NOR2_X1 U11270 ( .A1(n2464), .A2(n2778), .ZN(\mult_22/ab[7][14] ) );
  NOR2_X1 U11271 ( .A1(n2452), .A2(n2790), .ZN(\mult_22/ab[9][12] ) );
  NOR2_X1 U11272 ( .A1(n2440), .A2(n2802), .ZN(\mult_22/ab[11][10] ) );
  NOR2_X1 U11273 ( .A1(n2432), .A2(n2819), .ZN(\mult_22/ab[13][8] ) );
  NOR2_X1 U11274 ( .A1(n2420), .A2(n2831), .ZN(\mult_22/ab[15][6] ) );
  NOR2_X1 U11275 ( .A1(n2404), .A2(n2841), .ZN(\mult_22/ab[17][4] ) );
  NOR2_X1 U11276 ( .A1(n2584), .A2(n3062), .ZN(\mult_22/ab[54][34] ) );
  NOR2_X1 U11277 ( .A1(n2614), .A2(n2960), .ZN(\mult_22/ab[37][39] ) );
  NOR2_X1 U11278 ( .A1(n2626), .A2(n2948), .ZN(\mult_22/ab[35][41] ) );
  NOR2_X1 U11279 ( .A1(n2638), .A2(n2937), .ZN(\mult_22/ab[33][43] ) );
  NOR2_X1 U11280 ( .A1(n2649), .A2(n2925), .ZN(\mult_22/ab[31][45] ) );
  NOR2_X1 U11281 ( .A1(n2663), .A2(n2913), .ZN(\mult_22/ab[29][47] ) );
  NOR2_X1 U11282 ( .A1(n2673), .A2(n2901), .ZN(\mult_22/ab[27][49] ) );
  NOR2_X1 U11283 ( .A1(n2688), .A2(n2889), .ZN(\mult_22/ab[25][51] ) );
  NOR2_X1 U11284 ( .A1(n2696), .A2(n2877), .ZN(\mult_22/ab[23][53] ) );
  NOR2_X1 U11285 ( .A1(n2710), .A2(n2866), .ZN(\mult_22/ab[21][55] ) );
  NOR2_X1 U11286 ( .A1(n2716), .A2(n2854), .ZN(\mult_22/ab[19][57] ) );
  NOR2_X1 U11287 ( .A1(n2729), .A2(n2842), .ZN(\mult_22/ab[17][59] ) );
  NOR2_X1 U11288 ( .A1(n2620), .A2(n2954), .ZN(\mult_22/ab[36][40] ) );
  NOR2_X1 U11289 ( .A1(n2633), .A2(n2943), .ZN(\mult_22/ab[34][42] ) );
  NOR2_X1 U11290 ( .A1(n2645), .A2(n2931), .ZN(\mult_22/ab[32][44] ) );
  NOR2_X1 U11291 ( .A1(n2657), .A2(n2919), .ZN(\mult_22/ab[30][46] ) );
  NOR2_X1 U11292 ( .A1(n2669), .A2(n2907), .ZN(\mult_22/ab[28][48] ) );
  NOR2_X1 U11293 ( .A1(n2681), .A2(n2895), .ZN(\mult_22/ab[26][50] ) );
  NOR2_X1 U11294 ( .A1(n2691), .A2(n2883), .ZN(\mult_22/ab[24][52] ) );
  NOR2_X1 U11295 ( .A1(n2704), .A2(n2872), .ZN(\mult_22/ab[22][54] ) );
  NOR2_X1 U11296 ( .A1(n2719), .A2(n2848), .ZN(\mult_22/ab[18][58] ) );
  NOR2_X1 U11297 ( .A1(n2731), .A2(n2836), .ZN(\mult_22/ab[16][60] ) );
  NOR2_X1 U11298 ( .A1(n2555), .A2(n3055), .ZN(\mult_22/ab[53][29] ) );
  NOR2_X1 U11299 ( .A1(n2484), .A2(n2754), .ZN(\mult_22/ab[3][17] ) );
  NOR2_X1 U11300 ( .A1(n2470), .A2(n2766), .ZN(\mult_22/ab[5][15] ) );
  NOR2_X1 U11301 ( .A1(n2458), .A2(n2778), .ZN(\mult_22/ab[7][13] ) );
  NOR2_X1 U11302 ( .A1(n2446), .A2(n2790), .ZN(\mult_22/ab[9][11] ) );
  NOR2_X1 U11303 ( .A1(n2439), .A2(n2807), .ZN(\mult_22/ab[11][9] ) );
  NOR2_X1 U11304 ( .A1(n2426), .A2(n2819), .ZN(\mult_22/ab[13][7] ) );
  NOR2_X1 U11305 ( .A1(n2414), .A2(n2830), .ZN(\mult_22/ab[15][5] ) );
  NOR2_X1 U11306 ( .A1(n2739), .A2(n2830), .ZN(\mult_22/ab[15][61] ) );
  NOR2_X1 U11307 ( .A1(n2561), .A2(n3019), .ZN(\mult_22/ab[47][30] ) );
  NOR2_X1 U11308 ( .A1(n2575), .A2(n3008), .ZN(\mult_22/ab[45][32] ) );
  NOR2_X1 U11309 ( .A1(n2585), .A2(n2996), .ZN(\mult_22/ab[43][34] ) );
  NOR2_X1 U11310 ( .A1(n2478), .A2(n2754), .ZN(\mult_22/ab[3][16] ) );
  NOR2_X1 U11311 ( .A1(n2555), .A2(n3025), .ZN(\mult_22/ab[48][29] ) );
  NOR2_X1 U11312 ( .A1(n2464), .A2(n2766), .ZN(\mult_22/ab[5][14] ) );
  NOR2_X1 U11313 ( .A1(n2568), .A2(n3014), .ZN(\mult_22/ab[46][31] ) );
  NOR2_X1 U11314 ( .A1(n2579), .A2(n3002), .ZN(\mult_22/ab[44][33] ) );
  NOR2_X1 U11315 ( .A1(n2597), .A2(n2984), .ZN(\mult_22/ab[41][36] ) );
  NOR2_X1 U11316 ( .A1(n2609), .A2(n2972), .ZN(\mult_22/ab[39][38] ) );
  NOR2_X1 U11317 ( .A1(n2452), .A2(n2778), .ZN(\mult_22/ab[7][12] ) );
  NOR2_X1 U11318 ( .A1(n2445), .A2(n2790), .ZN(\mult_22/ab[9][10] ) );
  NOR2_X1 U11319 ( .A1(n2591), .A2(n2990), .ZN(\mult_22/ab[42][35] ) );
  NOR2_X1 U11320 ( .A1(n2433), .A2(n2807), .ZN(\mult_22/ab[11][8] ) );
  NOR2_X1 U11321 ( .A1(n2603), .A2(n2978), .ZN(\mult_22/ab[40][37] ) );
  NOR2_X1 U11322 ( .A1(n2420), .A2(n2819), .ZN(\mult_22/ab[13][6] ) );
  NOR2_X1 U11323 ( .A1(n2404), .A2(n2829), .ZN(\mult_22/ab[15][4] ) );
  NOR2_X1 U11324 ( .A1(n2465), .A2(n2760), .ZN(\mult_22/ab[4][14] ) );
  NOR2_X1 U11325 ( .A1(n2452), .A2(n2772), .ZN(\mult_22/ab[6][12] ) );
  NOR2_X1 U11326 ( .A1(n2445), .A2(n2784), .ZN(\mult_22/ab[8][10] ) );
  NOR2_X1 U11327 ( .A1(n2433), .A2(n2801), .ZN(\mult_22/ab[10][8] ) );
  NOR2_X1 U11328 ( .A1(n2421), .A2(n2813), .ZN(\mult_22/ab[12][6] ) );
  NOR2_X1 U11329 ( .A1(n2404), .A2(n2823), .ZN(\mult_22/ab[14][4] ) );
  NOR2_X1 U11330 ( .A1(n2466), .A2(n2754), .ZN(\mult_22/ab[3][14] ) );
  NOR2_X1 U11331 ( .A1(n2452), .A2(n2766), .ZN(\mult_22/ab[5][12] ) );
  NOR2_X1 U11332 ( .A1(n2444), .A2(n2778), .ZN(\mult_22/ab[7][10] ) );
  NOR2_X1 U11333 ( .A1(n2428), .A2(n2795), .ZN(\mult_22/ab[9][8] ) );
  NOR2_X1 U11334 ( .A1(n2421), .A2(n2806), .ZN(\mult_22/ab[11][6] ) );
  NOR2_X1 U11335 ( .A1(n2404), .A2(n2817), .ZN(\mult_22/ab[13][4] ) );
  NOR2_X1 U11336 ( .A1(n2614), .A2(n2966), .ZN(\mult_22/ab[38][39] ) );
  NOR2_X1 U11337 ( .A1(n2626), .A2(n2954), .ZN(\mult_22/ab[36][41] ) );
  NOR2_X1 U11338 ( .A1(n2638), .A2(n2943), .ZN(\mult_22/ab[34][43] ) );
  NOR2_X1 U11339 ( .A1(n2649), .A2(n2931), .ZN(\mult_22/ab[32][45] ) );
  NOR2_X1 U11340 ( .A1(n2663), .A2(n2919), .ZN(\mult_22/ab[30][47] ) );
  NOR2_X1 U11341 ( .A1(n2673), .A2(n2907), .ZN(\mult_22/ab[28][49] ) );
  NOR2_X1 U11342 ( .A1(n2688), .A2(n2895), .ZN(\mult_22/ab[26][51] ) );
  NOR2_X1 U11343 ( .A1(n2697), .A2(n2883), .ZN(\mult_22/ab[24][53] ) );
  NOR2_X1 U11344 ( .A1(n2710), .A2(n2872), .ZN(\mult_22/ab[22][55] ) );
  NOR2_X1 U11345 ( .A1(n2716), .A2(n2860), .ZN(\mult_22/ab[20][57] ) );
  NOR2_X1 U11346 ( .A1(n2730), .A2(n2848), .ZN(\mult_22/ab[18][59] ) );
  NOR2_X1 U11347 ( .A1(n2620), .A2(n2960), .ZN(\mult_22/ab[37][40] ) );
  NOR2_X1 U11348 ( .A1(n2633), .A2(n2949), .ZN(\mult_22/ab[35][42] ) );
  NOR2_X1 U11349 ( .A1(n2645), .A2(n2937), .ZN(\mult_22/ab[33][44] ) );
  NOR2_X1 U11350 ( .A1(n2657), .A2(n2925), .ZN(\mult_22/ab[31][46] ) );
  NOR2_X1 U11351 ( .A1(n2669), .A2(n2913), .ZN(\mult_22/ab[29][48] ) );
  NOR2_X1 U11352 ( .A1(n2681), .A2(n2901), .ZN(\mult_22/ab[27][50] ) );
  NOR2_X1 U11353 ( .A1(n2691), .A2(n2889), .ZN(\mult_22/ab[25][52] ) );
  NOR2_X1 U11354 ( .A1(n2704), .A2(n2878), .ZN(\mult_22/ab[23][54] ) );
  NOR2_X1 U11355 ( .A1(n2712), .A2(n2866), .ZN(\mult_22/ab[21][56] ) );
  NOR2_X1 U11356 ( .A1(n2719), .A2(n2854), .ZN(\mult_22/ab[19][58] ) );
  NOR2_X1 U11357 ( .A1(n2731), .A2(n2842), .ZN(\mult_22/ab[17][60] ) );
  NOR2_X1 U11358 ( .A1(n2738), .A2(n2836), .ZN(\mult_22/ab[16][61] ) );
  NOR2_X1 U11359 ( .A1(n2460), .A2(n2754), .ZN(\mult_22/ab[3][13] ) );
  NOR2_X1 U11360 ( .A1(n2446), .A2(n2766), .ZN(\mult_22/ab[5][11] ) );
  NOR2_X1 U11361 ( .A1(n2434), .A2(n2783), .ZN(\mult_22/ab[7][9] ) );
  NOR2_X1 U11362 ( .A1(n2422), .A2(n2795), .ZN(\mult_22/ab[9][7] ) );
  NOR2_X1 U11363 ( .A1(n2415), .A2(n2806), .ZN(\mult_22/ab[11][5] ) );
  NOR2_X1 U11364 ( .A1(n2454), .A2(n2754), .ZN(\mult_22/ab[3][12] ) );
  NOR2_X1 U11365 ( .A1(n2444), .A2(n2766), .ZN(\mult_22/ab[5][10] ) );
  NOR2_X1 U11366 ( .A1(n2428), .A2(n2783), .ZN(\mult_22/ab[7][8] ) );
  NOR2_X1 U11367 ( .A1(n2416), .A2(n2795), .ZN(\mult_22/ab[9][6] ) );
  NOR2_X1 U11368 ( .A1(n2404), .A2(n2805), .ZN(\mult_22/ab[11][4] ) );
  NOR2_X1 U11369 ( .A1(n2443), .A2(n2760), .ZN(\mult_22/ab[4][10] ) );
  NOR2_X1 U11370 ( .A1(n2428), .A2(n2777), .ZN(\mult_22/ab[6][8] ) );
  NOR2_X1 U11371 ( .A1(n2416), .A2(n2788), .ZN(\mult_22/ab[8][6] ) );
  NOR2_X1 U11372 ( .A1(n2561), .A2(n3055), .ZN(\mult_22/ab[53][30] ) );
  NOR2_X1 U11373 ( .A1(n2404), .A2(n2799), .ZN(\mult_22/ab[10][4] ) );
  NOR2_X1 U11374 ( .A1(n2442), .A2(n2754), .ZN(\mult_22/ab[3][10] ) );
  NOR2_X1 U11375 ( .A1(n2428), .A2(n2771), .ZN(\mult_22/ab[5][8] ) );
  NOR2_X1 U11376 ( .A1(n2416), .A2(n2783), .ZN(\mult_22/ab[7][6] ) );
  NOR2_X1 U11377 ( .A1(n2409), .A2(n2793), .ZN(\mult_22/ab[9][4] ) );
  NOR2_X1 U11378 ( .A1(n2555), .A2(n3031), .ZN(\mult_22/ab[49][29] ) );
  NOR2_X1 U11379 ( .A1(n2568), .A2(n3020), .ZN(\mult_22/ab[47][31] ) );
  NOR2_X1 U11380 ( .A1(n2579), .A2(n3008), .ZN(\mult_22/ab[45][33] ) );
  NOR2_X1 U11381 ( .A1(n2591), .A2(n2996), .ZN(\mult_22/ab[43][35] ) );
  NOR2_X1 U11382 ( .A1(n2603), .A2(n2984), .ZN(\mult_22/ab[41][37] ) );
  NOR2_X1 U11383 ( .A1(n2561), .A2(n3025), .ZN(\mult_22/ab[48][30] ) );
  NOR2_X1 U11384 ( .A1(n2575), .A2(n3014), .ZN(\mult_22/ab[46][32] ) );
  NOR2_X1 U11385 ( .A1(n2585), .A2(n3002), .ZN(\mult_22/ab[44][34] ) );
  NOR2_X1 U11386 ( .A1(n2555), .A2(n3049), .ZN(\mult_22/ab[52][29] ) );
  NOR2_X1 U11387 ( .A1(n2597), .A2(n2990), .ZN(\mult_22/ab[42][36] ) );
  NOR2_X1 U11388 ( .A1(n2609), .A2(n2978), .ZN(\mult_22/ab[40][38] ) );
  NOR2_X1 U11389 ( .A1(n2429), .A2(n2765), .ZN(\mult_22/ab[4][8] ) );
  NOR2_X1 U11390 ( .A1(n2416), .A2(n2777), .ZN(\mult_22/ab[6][6] ) );
  NOR2_X1 U11391 ( .A1(n2409), .A2(n2787), .ZN(\mult_22/ab[8][4] ) );
  NOR2_X1 U11392 ( .A1(n2614), .A2(n2972), .ZN(\mult_22/ab[39][39] ) );
  NOR2_X1 U11393 ( .A1(n2626), .A2(n2960), .ZN(\mult_22/ab[37][41] ) );
  NOR2_X1 U11394 ( .A1(n2638), .A2(n2949), .ZN(\mult_22/ab[35][43] ) );
  NOR2_X1 U11395 ( .A1(n2650), .A2(n2937), .ZN(\mult_22/ab[33][45] ) );
  NOR2_X1 U11396 ( .A1(n2663), .A2(n2925), .ZN(\mult_22/ab[31][47] ) );
  NOR2_X1 U11397 ( .A1(n2673), .A2(n2913), .ZN(\mult_22/ab[29][49] ) );
  NOR2_X1 U11398 ( .A1(n2687), .A2(n2901), .ZN(\mult_22/ab[27][51] ) );
  NOR2_X1 U11399 ( .A1(n2700), .A2(n2889), .ZN(\mult_22/ab[25][53] ) );
  NOR2_X1 U11400 ( .A1(n2710), .A2(n2878), .ZN(\mult_22/ab[23][55] ) );
  NOR2_X1 U11401 ( .A1(n2716), .A2(n2866), .ZN(\mult_22/ab[21][57] ) );
  NOR2_X1 U11402 ( .A1(n2725), .A2(n2854), .ZN(\mult_22/ab[19][59] ) );
  NOR2_X1 U11403 ( .A1(n2620), .A2(n2966), .ZN(\mult_22/ab[38][40] ) );
  NOR2_X1 U11404 ( .A1(n2633), .A2(n2955), .ZN(\mult_22/ab[36][42] ) );
  NOR2_X1 U11405 ( .A1(n2645), .A2(n2943), .ZN(\mult_22/ab[34][44] ) );
  NOR2_X1 U11406 ( .A1(n2657), .A2(n2931), .ZN(\mult_22/ab[32][46] ) );
  NOR2_X1 U11407 ( .A1(n2669), .A2(n2919), .ZN(\mult_22/ab[30][48] ) );
  NOR2_X1 U11408 ( .A1(n2681), .A2(n2907), .ZN(\mult_22/ab[28][50] ) );
  NOR2_X1 U11409 ( .A1(n2691), .A2(n2895), .ZN(\mult_22/ab[26][52] ) );
  NOR2_X1 U11410 ( .A1(n2430), .A2(n2759), .ZN(\mult_22/ab[3][8] ) );
  NOR2_X1 U11411 ( .A1(n2704), .A2(n2884), .ZN(\mult_22/ab[24][54] ) );
  NOR2_X1 U11412 ( .A1(n2416), .A2(n2771), .ZN(\mult_22/ab[5][6] ) );
  NOR2_X1 U11413 ( .A1(n2712), .A2(n2872), .ZN(\mult_22/ab[22][56] ) );
  NOR2_X1 U11414 ( .A1(n2408), .A2(n2781), .ZN(\mult_22/ab[7][4] ) );
  NOR2_X1 U11415 ( .A1(n2719), .A2(n2860), .ZN(\mult_22/ab[20][58] ) );
  NOR2_X1 U11416 ( .A1(n2731), .A2(n2848), .ZN(\mult_22/ab[18][60] ) );
  NOR2_X1 U11417 ( .A1(n2739), .A2(n2842), .ZN(\mult_22/ab[17][61] ) );
  NOR2_X1 U11418 ( .A1(n2424), .A2(n2759), .ZN(\mult_22/ab[3][7] ) );
  NOR2_X1 U11419 ( .A1(n2410), .A2(n2770), .ZN(\mult_22/ab[5][5] ) );
  NOR2_X1 U11420 ( .A1(n2555), .A2(n3043), .ZN(\mult_22/ab[51][29] ) );
  NOR2_X1 U11421 ( .A1(n2561), .A2(n3031), .ZN(\mult_22/ab[49][30] ) );
  NOR2_X1 U11422 ( .A1(n2575), .A2(n3020), .ZN(\mult_22/ab[47][32] ) );
  NOR2_X1 U11423 ( .A1(n2585), .A2(n3008), .ZN(\mult_22/ab[45][34] ) );
  NOR2_X1 U11424 ( .A1(n2597), .A2(n2996), .ZN(\mult_22/ab[43][36] ) );
  NOR2_X1 U11425 ( .A1(n2555), .A2(n3037), .ZN(\mult_22/ab[50][29] ) );
  NOR2_X1 U11426 ( .A1(n2567), .A2(n3026), .ZN(\mult_22/ab[48][31] ) );
  NOR2_X1 U11427 ( .A1(n2579), .A2(n3014), .ZN(\mult_22/ab[46][33] ) );
  NOR2_X1 U11428 ( .A1(n2591), .A2(n3002), .ZN(\mult_22/ab[44][35] ) );
  NOR2_X1 U11429 ( .A1(n2603), .A2(n2990), .ZN(\mult_22/ab[42][37] ) );
  NOR2_X1 U11430 ( .A1(n2411), .A2(n2764), .ZN(\mult_22/ab[4][5] ) );
  NOR2_X1 U11431 ( .A1(n2412), .A2(n2758), .ZN(\mult_22/ab[3][5] ) );
  NOR2_X1 U11432 ( .A1(n2609), .A2(n2984), .ZN(\mult_22/ab[41][38] ) );
  NOR2_X1 U11433 ( .A1(n2614), .A2(n2978), .ZN(\mult_22/ab[40][39] ) );
  NOR2_X1 U11434 ( .A1(n2626), .A2(n2966), .ZN(\mult_22/ab[38][41] ) );
  NOR2_X1 U11435 ( .A1(n2638), .A2(n2955), .ZN(\mult_22/ab[36][43] ) );
  NOR2_X1 U11436 ( .A1(n2650), .A2(n2943), .ZN(\mult_22/ab[34][45] ) );
  NOR2_X1 U11437 ( .A1(n2663), .A2(n2931), .ZN(\mult_22/ab[32][47] ) );
  NOR2_X1 U11438 ( .A1(n2673), .A2(n2919), .ZN(\mult_22/ab[30][49] ) );
  NOR2_X1 U11439 ( .A1(n2687), .A2(n2907), .ZN(\mult_22/ab[28][51] ) );
  NOR2_X1 U11440 ( .A1(n2695), .A2(n2896), .ZN(\mult_22/ab[26][53] ) );
  NOR2_X1 U11441 ( .A1(n2710), .A2(n2884), .ZN(\mult_22/ab[24][55] ) );
  NOR2_X1 U11442 ( .A1(n2716), .A2(n2872), .ZN(\mult_22/ab[22][57] ) );
  NOR2_X1 U11443 ( .A1(n2726), .A2(n2860), .ZN(\mult_22/ab[20][59] ) );
  NOR2_X1 U11444 ( .A1(n2620), .A2(n2972), .ZN(\mult_22/ab[39][40] ) );
  NOR2_X1 U11445 ( .A1(n2632), .A2(n2961), .ZN(\mult_22/ab[37][42] ) );
  NOR2_X1 U11446 ( .A1(n2645), .A2(n2949), .ZN(\mult_22/ab[35][44] ) );
  NOR2_X1 U11447 ( .A1(n2657), .A2(n2937), .ZN(\mult_22/ab[33][46] ) );
  NOR2_X1 U11448 ( .A1(n2669), .A2(n2925), .ZN(\mult_22/ab[31][48] ) );
  NOR2_X1 U11449 ( .A1(n2681), .A2(n2913), .ZN(\mult_22/ab[29][50] ) );
  NOR2_X1 U11450 ( .A1(n2691), .A2(n2901), .ZN(\mult_22/ab[27][52] ) );
  NOR2_X1 U11451 ( .A1(n2712), .A2(n2878), .ZN(\mult_22/ab[23][56] ) );
  NOR2_X1 U11452 ( .A1(n2719), .A2(n2866), .ZN(\mult_22/ab[21][58] ) );
  NOR2_X1 U11453 ( .A1(n2731), .A2(n2854), .ZN(\mult_22/ab[19][60] ) );
  NOR2_X1 U11454 ( .A1(n2737), .A2(n2848), .ZN(\mult_22/ab[18][61] ) );
  NOR2_X1 U11455 ( .A1(n2406), .A2(n2757), .ZN(\mult_22/ab[3][4] ) );
  NOR2_X1 U11456 ( .A1(n2567), .A2(n3032), .ZN(\mult_22/ab[49][31] ) );
  NOR2_X1 U11457 ( .A1(n2579), .A2(n3020), .ZN(\mult_22/ab[47][33] ) );
  NOR2_X1 U11458 ( .A1(n2591), .A2(n3008), .ZN(\mult_22/ab[45][35] ) );
  NOR2_X1 U11459 ( .A1(n2603), .A2(n2996), .ZN(\mult_22/ab[43][37] ) );
  NOR2_X1 U11460 ( .A1(n2561), .A2(n3037), .ZN(\mult_22/ab[50][30] ) );
  NOR2_X1 U11461 ( .A1(n2575), .A2(n3026), .ZN(\mult_22/ab[48][32] ) );
  NOR2_X1 U11462 ( .A1(n2585), .A2(n3014), .ZN(\mult_22/ab[46][34] ) );
  NOR2_X1 U11463 ( .A1(n2597), .A2(n3002), .ZN(\mult_22/ab[44][36] ) );
  NOR2_X1 U11464 ( .A1(n2609), .A2(n2990), .ZN(\mult_22/ab[42][38] ) );
  NOR2_X1 U11465 ( .A1(n2614), .A2(n2984), .ZN(\mult_22/ab[41][39] ) );
  NOR2_X1 U11466 ( .A1(n2626), .A2(n2972), .ZN(\mult_22/ab[39][41] ) );
  NOR2_X1 U11467 ( .A1(n2638), .A2(n2961), .ZN(\mult_22/ab[37][43] ) );
  NOR2_X1 U11468 ( .A1(n2650), .A2(n2949), .ZN(\mult_22/ab[35][45] ) );
  NOR2_X1 U11469 ( .A1(n2663), .A2(n2937), .ZN(\mult_22/ab[33][47] ) );
  NOR2_X1 U11470 ( .A1(n2673), .A2(n2925), .ZN(\mult_22/ab[31][49] ) );
  NOR2_X1 U11471 ( .A1(n2687), .A2(n2913), .ZN(\mult_22/ab[29][51] ) );
  NOR2_X1 U11472 ( .A1(n2367), .A2(n2902), .ZN(\mult_22/ab[27][53] ) );
  NOR2_X1 U11473 ( .A1(n2710), .A2(n2890), .ZN(\mult_22/ab[25][55] ) );
  NOR2_X1 U11474 ( .A1(n2716), .A2(n2878), .ZN(\mult_22/ab[23][57] ) );
  NOR2_X1 U11475 ( .A1(n2727), .A2(n2866), .ZN(\mult_22/ab[21][59] ) );
  NOR2_X1 U11476 ( .A1(n2620), .A2(n2978), .ZN(\mult_22/ab[40][40] ) );
  NOR2_X1 U11477 ( .A1(n2632), .A2(n2967), .ZN(\mult_22/ab[38][42] ) );
  NOR2_X1 U11478 ( .A1(n2645), .A2(n2955), .ZN(\mult_22/ab[36][44] ) );
  NOR2_X1 U11479 ( .A1(n2657), .A2(n2943), .ZN(\mult_22/ab[34][46] ) );
  NOR2_X1 U11480 ( .A1(n2669), .A2(n2931), .ZN(\mult_22/ab[32][48] ) );
  NOR2_X1 U11481 ( .A1(n2681), .A2(n2919), .ZN(\mult_22/ab[30][50] ) );
  NOR2_X1 U11482 ( .A1(n2691), .A2(n2907), .ZN(\mult_22/ab[28][52] ) );
  NOR2_X1 U11483 ( .A1(n2712), .A2(n2884), .ZN(\mult_22/ab[24][56] ) );
  NOR2_X1 U11484 ( .A1(n2720), .A2(n2872), .ZN(\mult_22/ab[22][58] ) );
  NOR2_X1 U11485 ( .A1(n2731), .A2(n2860), .ZN(\mult_22/ab[20][60] ) );
  NOR2_X1 U11486 ( .A1(n2738), .A2(n2854), .ZN(\mult_22/ab[19][61] ) );
  NOR2_X1 U11487 ( .A1(n2584), .A2(n3056), .ZN(\mult_22/ab[53][34] ) );
  NOR2_X1 U11488 ( .A1(n2567), .A2(n3038), .ZN(\mult_22/ab[50][31] ) );
  NOR2_X1 U11489 ( .A1(n2578), .A2(n3026), .ZN(\mult_22/ab[48][33] ) );
  NOR2_X1 U11490 ( .A1(n2591), .A2(n3014), .ZN(\mult_22/ab[46][35] ) );
  NOR2_X1 U11491 ( .A1(n2603), .A2(n3002), .ZN(\mult_22/ab[44][37] ) );
  NOR2_X1 U11492 ( .A1(n2561), .A2(n3043), .ZN(\mult_22/ab[51][30] ) );
  NOR2_X1 U11493 ( .A1(n2575), .A2(n3032), .ZN(\mult_22/ab[49][32] ) );
  NOR2_X1 U11494 ( .A1(n2584), .A2(n3020), .ZN(\mult_22/ab[47][34] ) );
  NOR2_X1 U11495 ( .A1(n2567), .A2(n3044), .ZN(\mult_22/ab[51][31] ) );
  NOR2_X1 U11496 ( .A1(n2578), .A2(n3032), .ZN(\mult_22/ab[49][33] ) );
  NOR2_X1 U11497 ( .A1(n2590), .A2(n3020), .ZN(\mult_22/ab[47][35] ) );
  NOR2_X1 U11498 ( .A1(n2603), .A2(n3008), .ZN(\mult_22/ab[45][37] ) );
  NOR2_X1 U11499 ( .A1(n2597), .A2(n3008), .ZN(\mult_22/ab[45][36] ) );
  NOR2_X1 U11500 ( .A1(n2561), .A2(n3049), .ZN(\mult_22/ab[52][30] ) );
  NOR2_X1 U11501 ( .A1(n2575), .A2(n3038), .ZN(\mult_22/ab[50][32] ) );
  NOR2_X1 U11502 ( .A1(n2584), .A2(n3026), .ZN(\mult_22/ab[48][34] ) );
  NOR2_X1 U11503 ( .A1(n2614), .A2(n2990), .ZN(\mult_22/ab[42][39] ) );
  NOR2_X1 U11504 ( .A1(n2626), .A2(n2978), .ZN(\mult_22/ab[40][41] ) );
  NOR2_X1 U11505 ( .A1(n2597), .A2(n3014), .ZN(\mult_22/ab[46][36] ) );
  NOR2_X1 U11506 ( .A1(n2638), .A2(n2967), .ZN(\mult_22/ab[38][43] ) );
  NOR2_X1 U11507 ( .A1(n2650), .A2(n2955), .ZN(\mult_22/ab[36][45] ) );
  NOR2_X1 U11508 ( .A1(n2663), .A2(n2943), .ZN(\mult_22/ab[34][47] ) );
  NOR2_X1 U11509 ( .A1(n2673), .A2(n2931), .ZN(\mult_22/ab[32][49] ) );
  NOR2_X1 U11510 ( .A1(n2687), .A2(n2919), .ZN(\mult_22/ab[30][51] ) );
  NOR2_X1 U11511 ( .A1(n2699), .A2(n2907), .ZN(\mult_22/ab[28][53] ) );
  NOR2_X1 U11512 ( .A1(n2709), .A2(n2896), .ZN(\mult_22/ab[26][55] ) );
  NOR2_X1 U11513 ( .A1(n2716), .A2(n2884), .ZN(\mult_22/ab[24][57] ) );
  NOR2_X1 U11514 ( .A1(n2728), .A2(n2872), .ZN(\mult_22/ab[22][59] ) );
  NOR2_X1 U11515 ( .A1(n2609), .A2(n2996), .ZN(\mult_22/ab[43][38] ) );
  NOR2_X1 U11516 ( .A1(n2609), .A2(n3002), .ZN(\mult_22/ab[44][38] ) );
  NOR2_X1 U11517 ( .A1(n2614), .A2(n2996), .ZN(\mult_22/ab[43][39] ) );
  NOR2_X1 U11518 ( .A1(n2626), .A2(n2984), .ZN(\mult_22/ab[41][41] ) );
  NOR2_X1 U11519 ( .A1(n2638), .A2(n2973), .ZN(\mult_22/ab[39][43] ) );
  NOR2_X1 U11520 ( .A1(n2650), .A2(n2961), .ZN(\mult_22/ab[37][45] ) );
  NOR2_X1 U11521 ( .A1(n2663), .A2(n2949), .ZN(\mult_22/ab[35][47] ) );
  NOR2_X1 U11522 ( .A1(n2674), .A2(n2937), .ZN(\mult_22/ab[33][49] ) );
  NOR2_X1 U11523 ( .A1(n2687), .A2(n2925), .ZN(\mult_22/ab[31][51] ) );
  NOR2_X1 U11524 ( .A1(n2696), .A2(n2914), .ZN(\mult_22/ab[29][53] ) );
  NOR2_X1 U11525 ( .A1(n2709), .A2(n2902), .ZN(\mult_22/ab[27][55] ) );
  NOR2_X1 U11526 ( .A1(n2716), .A2(n2890), .ZN(\mult_22/ab[25][57] ) );
  NOR2_X1 U11527 ( .A1(n2729), .A2(n2878), .ZN(\mult_22/ab[23][59] ) );
  NOR2_X1 U11528 ( .A1(n2620), .A2(n2984), .ZN(\mult_22/ab[41][40] ) );
  NOR2_X1 U11529 ( .A1(n2632), .A2(n2973), .ZN(\mult_22/ab[39][42] ) );
  NOR2_X1 U11530 ( .A1(n2644), .A2(n2961), .ZN(\mult_22/ab[37][44] ) );
  NOR2_X1 U11531 ( .A1(n2657), .A2(n2949), .ZN(\mult_22/ab[35][46] ) );
  NOR2_X1 U11532 ( .A1(n2669), .A2(n2937), .ZN(\mult_22/ab[33][48] ) );
  NOR2_X1 U11533 ( .A1(n2681), .A2(n2925), .ZN(\mult_22/ab[31][50] ) );
  NOR2_X1 U11534 ( .A1(n2691), .A2(n2913), .ZN(\mult_22/ab[29][52] ) );
  NOR2_X1 U11535 ( .A1(n2712), .A2(n2890), .ZN(\mult_22/ab[25][56] ) );
  NOR2_X1 U11536 ( .A1(n2720), .A2(n2878), .ZN(\mult_22/ab[23][58] ) );
  NOR2_X1 U11537 ( .A1(n2575), .A2(n3044), .ZN(\mult_22/ab[51][32] ) );
  NOR2_X1 U11538 ( .A1(n2584), .A2(n3032), .ZN(\mult_22/ab[49][34] ) );
  NOR2_X1 U11539 ( .A1(n2596), .A2(n3020), .ZN(\mult_22/ab[47][36] ) );
  NOR2_X1 U11540 ( .A1(n2740), .A2(n2860), .ZN(\mult_22/ab[20][61] ) );
  NOR2_X1 U11541 ( .A1(n2567), .A2(n3050), .ZN(\mult_22/ab[52][31] ) );
  NOR2_X1 U11542 ( .A1(n2578), .A2(n3038), .ZN(\mult_22/ab[50][33] ) );
  NOR2_X1 U11543 ( .A1(n2590), .A2(n3026), .ZN(\mult_22/ab[48][35] ) );
  NOR2_X1 U11544 ( .A1(n2603), .A2(n3014), .ZN(\mult_22/ab[46][37] ) );
  NOR2_X1 U11545 ( .A1(n2620), .A2(n2990), .ZN(\mult_22/ab[42][40] ) );
  NOR2_X1 U11546 ( .A1(n2632), .A2(n2979), .ZN(\mult_22/ab[40][42] ) );
  NOR2_X1 U11547 ( .A1(n2644), .A2(n2967), .ZN(\mult_22/ab[38][44] ) );
  NOR2_X1 U11548 ( .A1(n2656), .A2(n2955), .ZN(\mult_22/ab[36][46] ) );
  NOR2_X1 U11549 ( .A1(n2669), .A2(n2943), .ZN(\mult_22/ab[34][48] ) );
  NOR2_X1 U11550 ( .A1(n2681), .A2(n2931), .ZN(\mult_22/ab[32][50] ) );
  NOR2_X1 U11551 ( .A1(n2691), .A2(n2919), .ZN(\mult_22/ab[30][52] ) );
  NOR2_X1 U11552 ( .A1(n2712), .A2(n2896), .ZN(\mult_22/ab[26][56] ) );
  NOR2_X1 U11553 ( .A1(n2720), .A2(n2884), .ZN(\mult_22/ab[24][58] ) );
  NOR2_X1 U11554 ( .A1(n2731), .A2(n2866), .ZN(\mult_22/ab[21][60] ) );
  NOR2_X1 U11555 ( .A1(n2609), .A2(n3008), .ZN(\mult_22/ab[45][38] ) );
  NOR2_X1 U11556 ( .A1(n2741), .A2(n2866), .ZN(\mult_22/ab[21][61] ) );
  NOR2_X1 U11557 ( .A1(n2732), .A2(n2872), .ZN(\mult_22/ab[22][60] ) );
  NOR2_X1 U11558 ( .A1(n2614), .A2(n3002), .ZN(\mult_22/ab[44][39] ) );
  NOR2_X1 U11559 ( .A1(n2626), .A2(n2990), .ZN(\mult_22/ab[42][41] ) );
  NOR2_X1 U11560 ( .A1(n2638), .A2(n2979), .ZN(\mult_22/ab[40][43] ) );
  NOR2_X1 U11561 ( .A1(n2650), .A2(n2967), .ZN(\mult_22/ab[38][45] ) );
  NOR2_X1 U11562 ( .A1(n2663), .A2(n2955), .ZN(\mult_22/ab[36][47] ) );
  NOR2_X1 U11563 ( .A1(n2674), .A2(n2943), .ZN(\mult_22/ab[34][49] ) );
  NOR2_X1 U11564 ( .A1(n2687), .A2(n2931), .ZN(\mult_22/ab[32][51] ) );
  NOR2_X1 U11565 ( .A1(n2697), .A2(n2920), .ZN(\mult_22/ab[30][53] ) );
  NOR2_X1 U11566 ( .A1(n2709), .A2(n2908), .ZN(\mult_22/ab[28][55] ) );
  NOR2_X1 U11567 ( .A1(n2716), .A2(n2896), .ZN(\mult_22/ab[26][57] ) );
  NOR2_X1 U11568 ( .A1(n2730), .A2(n2884), .ZN(\mult_22/ab[24][59] ) );
  NOR2_X1 U11569 ( .A1(n2620), .A2(n2996), .ZN(\mult_22/ab[43][40] ) );
  NOR2_X1 U11570 ( .A1(n2632), .A2(n2985), .ZN(\mult_22/ab[41][42] ) );
  NOR2_X1 U11571 ( .A1(n2644), .A2(n2973), .ZN(\mult_22/ab[39][44] ) );
  NOR2_X1 U11572 ( .A1(n2656), .A2(n2961), .ZN(\mult_22/ab[37][46] ) );
  NOR2_X1 U11573 ( .A1(n2669), .A2(n2949), .ZN(\mult_22/ab[35][48] ) );
  NOR2_X1 U11574 ( .A1(n2681), .A2(n2937), .ZN(\mult_22/ab[33][50] ) );
  NOR2_X1 U11575 ( .A1(n2691), .A2(n2925), .ZN(\mult_22/ab[31][52] ) );
  NOR2_X1 U11576 ( .A1(n2712), .A2(n2902), .ZN(\mult_22/ab[27][56] ) );
  NOR2_X1 U11577 ( .A1(n2720), .A2(n2890), .ZN(\mult_22/ab[25][58] ) );
  NOR2_X1 U11578 ( .A1(n2732), .A2(n2878), .ZN(\mult_22/ab[23][60] ) );
  NOR2_X1 U11579 ( .A1(n2737), .A2(n2872), .ZN(\mult_22/ab[22][61] ) );
  NOR2_X1 U11580 ( .A1(n2575), .A2(n3050), .ZN(\mult_22/ab[52][32] ) );
  NOR2_X1 U11581 ( .A1(n2584), .A2(n3038), .ZN(\mult_22/ab[50][34] ) );
  NOR2_X1 U11582 ( .A1(n2578), .A2(n3044), .ZN(\mult_22/ab[51][33] ) );
  NOR2_X1 U11583 ( .A1(n2590), .A2(n3032), .ZN(\mult_22/ab[49][35] ) );
  NOR2_X1 U11584 ( .A1(n2602), .A2(n3020), .ZN(\mult_22/ab[47][37] ) );
  NOR2_X1 U11585 ( .A1(n2596), .A2(n3026), .ZN(\mult_22/ab[48][36] ) );
  NOR2_X1 U11586 ( .A1(n2609), .A2(n3014), .ZN(\mult_22/ab[46][38] ) );
  NOR2_X1 U11587 ( .A1(n2614), .A2(n3008), .ZN(\mult_22/ab[45][39] ) );
  NOR2_X1 U11588 ( .A1(n2626), .A2(n2996), .ZN(\mult_22/ab[43][41] ) );
  NOR2_X1 U11589 ( .A1(n2638), .A2(n2985), .ZN(\mult_22/ab[41][43] ) );
  NOR2_X1 U11590 ( .A1(n2650), .A2(n2973), .ZN(\mult_22/ab[39][45] ) );
  NOR2_X1 U11591 ( .A1(n2662), .A2(n2961), .ZN(\mult_22/ab[37][47] ) );
  NOR2_X1 U11592 ( .A1(n2674), .A2(n2949), .ZN(\mult_22/ab[35][49] ) );
  NOR2_X1 U11593 ( .A1(n2687), .A2(n2937), .ZN(\mult_22/ab[33][51] ) );
  NOR2_X1 U11594 ( .A1(n2695), .A2(n2926), .ZN(\mult_22/ab[31][53] ) );
  NOR2_X1 U11595 ( .A1(n2709), .A2(n2914), .ZN(\mult_22/ab[29][55] ) );
  NOR2_X1 U11596 ( .A1(n2716), .A2(n2902), .ZN(\mult_22/ab[27][57] ) );
  NOR2_X1 U11597 ( .A1(n2725), .A2(n2890), .ZN(\mult_22/ab[25][59] ) );
  NOR2_X1 U11598 ( .A1(n2620), .A2(n3002), .ZN(\mult_22/ab[44][40] ) );
  NOR2_X1 U11599 ( .A1(n2632), .A2(n2991), .ZN(\mult_22/ab[42][42] ) );
  NOR2_X1 U11600 ( .A1(n2644), .A2(n2979), .ZN(\mult_22/ab[40][44] ) );
  NOR2_X1 U11601 ( .A1(n2656), .A2(n2967), .ZN(\mult_22/ab[38][46] ) );
  NOR2_X1 U11602 ( .A1(n2668), .A2(n2955), .ZN(\mult_22/ab[36][48] ) );
  NOR2_X1 U11603 ( .A1(n2681), .A2(n2943), .ZN(\mult_22/ab[34][50] ) );
  NOR2_X1 U11604 ( .A1(n2691), .A2(n2931), .ZN(\mult_22/ab[32][52] ) );
  NOR2_X1 U11605 ( .A1(n2712), .A2(n2908), .ZN(\mult_22/ab[28][56] ) );
  NOR2_X1 U11606 ( .A1(n2720), .A2(n2896), .ZN(\mult_22/ab[26][58] ) );
  NOR2_X1 U11607 ( .A1(n2732), .A2(n2884), .ZN(\mult_22/ab[24][60] ) );
  NOR2_X1 U11608 ( .A1(n2739), .A2(n2878), .ZN(\mult_22/ab[23][61] ) );
  NOR2_X1 U11609 ( .A1(n2584), .A2(n3044), .ZN(\mult_22/ab[51][34] ) );
  NOR2_X1 U11610 ( .A1(n2578), .A2(n3050), .ZN(\mult_22/ab[52][33] ) );
  NOR2_X1 U11611 ( .A1(n2590), .A2(n3038), .ZN(\mult_22/ab[50][35] ) );
  NOR2_X1 U11612 ( .A1(n2602), .A2(n3026), .ZN(\mult_22/ab[48][37] ) );
  NOR2_X1 U11613 ( .A1(n2596), .A2(n3032), .ZN(\mult_22/ab[49][36] ) );
  NOR2_X1 U11614 ( .A1(n2608), .A2(n3020), .ZN(\mult_22/ab[47][38] ) );
  NOR2_X1 U11615 ( .A1(n2590), .A2(n3044), .ZN(\mult_22/ab[51][35] ) );
  NOR2_X1 U11616 ( .A1(n2602), .A2(n3032), .ZN(\mult_22/ab[49][37] ) );
  NOR2_X1 U11617 ( .A1(n2584), .A2(n3050), .ZN(\mult_22/ab[52][34] ) );
  NOR2_X1 U11618 ( .A1(n2614), .A2(n3014), .ZN(\mult_22/ab[46][39] ) );
  NOR2_X1 U11619 ( .A1(n2627), .A2(n3002), .ZN(\mult_22/ab[44][41] ) );
  NOR2_X1 U11620 ( .A1(n2638), .A2(n2991), .ZN(\mult_22/ab[42][43] ) );
  NOR2_X1 U11621 ( .A1(n2650), .A2(n2979), .ZN(\mult_22/ab[40][45] ) );
  NOR2_X1 U11622 ( .A1(n2662), .A2(n2967), .ZN(\mult_22/ab[38][47] ) );
  NOR2_X1 U11623 ( .A1(n2674), .A2(n2955), .ZN(\mult_22/ab[36][49] ) );
  NOR2_X1 U11624 ( .A1(n2687), .A2(n2943), .ZN(\mult_22/ab[34][51] ) );
  NOR2_X1 U11625 ( .A1(n2700), .A2(n2932), .ZN(\mult_22/ab[32][53] ) );
  NOR2_X1 U11626 ( .A1(n2709), .A2(n2920), .ZN(\mult_22/ab[30][55] ) );
  NOR2_X1 U11627 ( .A1(n2716), .A2(n2908), .ZN(\mult_22/ab[28][57] ) );
  NOR2_X1 U11628 ( .A1(n2726), .A2(n2896), .ZN(\mult_22/ab[26][59] ) );
  NOR2_X1 U11629 ( .A1(n2596), .A2(n3038), .ZN(\mult_22/ab[50][36] ) );
  NOR2_X1 U11630 ( .A1(n2608), .A2(n3026), .ZN(\mult_22/ab[48][38] ) );
  NOR2_X1 U11631 ( .A1(n2620), .A2(n3008), .ZN(\mult_22/ab[45][40] ) );
  NOR2_X1 U11632 ( .A1(n2632), .A2(n2997), .ZN(\mult_22/ab[43][42] ) );
  NOR2_X1 U11633 ( .A1(n2644), .A2(n2985), .ZN(\mult_22/ab[41][44] ) );
  NOR2_X1 U11634 ( .A1(n2656), .A2(n2973), .ZN(\mult_22/ab[39][46] ) );
  NOR2_X1 U11635 ( .A1(n2668), .A2(n2961), .ZN(\mult_22/ab[37][48] ) );
  NOR2_X1 U11636 ( .A1(n2680), .A2(n2949), .ZN(\mult_22/ab[35][50] ) );
  NOR2_X1 U11637 ( .A1(n2692), .A2(n2937), .ZN(\mult_22/ab[33][52] ) );
  NOR2_X1 U11638 ( .A1(n2712), .A2(n2914), .ZN(\mult_22/ab[29][56] ) );
  NOR2_X1 U11639 ( .A1(n2720), .A2(n2902), .ZN(\mult_22/ab[27][58] ) );
  NOR2_X1 U11640 ( .A1(n2732), .A2(n2890), .ZN(\mult_22/ab[25][60] ) );
  NOR2_X1 U11641 ( .A1(n2613), .A2(n3020), .ZN(\mult_22/ab[47][39] ) );
  NOR2_X1 U11642 ( .A1(n2627), .A2(n3008), .ZN(\mult_22/ab[45][41] ) );
  NOR2_X1 U11643 ( .A1(n2638), .A2(n2997), .ZN(\mult_22/ab[43][43] ) );
  NOR2_X1 U11644 ( .A1(n2650), .A2(n2985), .ZN(\mult_22/ab[41][45] ) );
  NOR2_X1 U11645 ( .A1(n2662), .A2(n2973), .ZN(\mult_22/ab[39][47] ) );
  NOR2_X1 U11646 ( .A1(n2674), .A2(n2961), .ZN(\mult_22/ab[37][49] ) );
  NOR2_X1 U11647 ( .A1(n2687), .A2(n2949), .ZN(\mult_22/ab[35][51] ) );
  NOR2_X1 U11648 ( .A1(n2367), .A2(n2937), .ZN(\mult_22/ab[33][53] ) );
  NOR2_X1 U11649 ( .A1(n2709), .A2(n2926), .ZN(\mult_22/ab[31][55] ) );
  NOR2_X1 U11650 ( .A1(n2716), .A2(n2914), .ZN(\mult_22/ab[29][57] ) );
  NOR2_X1 U11651 ( .A1(n2727), .A2(n2902), .ZN(\mult_22/ab[27][59] ) );
  NOR2_X1 U11652 ( .A1(n2596), .A2(n3044), .ZN(\mult_22/ab[51][36] ) );
  NOR2_X1 U11653 ( .A1(n2738), .A2(n2884), .ZN(\mult_22/ab[24][61] ) );
  NOR2_X1 U11654 ( .A1(n2590), .A2(n3050), .ZN(\mult_22/ab[52][35] ) );
  NOR2_X1 U11655 ( .A1(n2602), .A2(n3038), .ZN(\mult_22/ab[50][37] ) );
  NOR2_X1 U11656 ( .A1(n2620), .A2(n3014), .ZN(\mult_22/ab[46][40] ) );
  NOR2_X1 U11657 ( .A1(n2632), .A2(n3003), .ZN(\mult_22/ab[44][42] ) );
  NOR2_X1 U11658 ( .A1(n2644), .A2(n2991), .ZN(\mult_22/ab[42][44] ) );
  NOR2_X1 U11659 ( .A1(n2656), .A2(n2979), .ZN(\mult_22/ab[40][46] ) );
  NOR2_X1 U11660 ( .A1(n2668), .A2(n2967), .ZN(\mult_22/ab[38][48] ) );
  NOR2_X1 U11661 ( .A1(n2680), .A2(n2955), .ZN(\mult_22/ab[36][50] ) );
  NOR2_X1 U11662 ( .A1(n2692), .A2(n2943), .ZN(\mult_22/ab[34][52] ) );
  NOR2_X1 U11663 ( .A1(n2712), .A2(n2920), .ZN(\mult_22/ab[30][56] ) );
  NOR2_X1 U11664 ( .A1(n2720), .A2(n2908), .ZN(\mult_22/ab[28][58] ) );
  NOR2_X1 U11665 ( .A1(n2608), .A2(n3032), .ZN(\mult_22/ab[49][38] ) );
  NOR2_X1 U11666 ( .A1(n2732), .A2(n2896), .ZN(\mult_22/ab[26][60] ) );
  NOR2_X1 U11667 ( .A1(n2739), .A2(n2890), .ZN(\mult_22/ab[25][61] ) );
  NOR2_X1 U11668 ( .A1(n2590), .A2(n3068), .ZN(\mult_22/ab[55][35] ) );
  NOR2_X1 U11669 ( .A1(n2613), .A2(n3026), .ZN(\mult_22/ab[48][39] ) );
  NOR2_X1 U11670 ( .A1(n2627), .A2(n3014), .ZN(\mult_22/ab[46][41] ) );
  NOR2_X1 U11671 ( .A1(n2639), .A2(n3003), .ZN(\mult_22/ab[44][43] ) );
  NOR2_X1 U11672 ( .A1(n2650), .A2(n2991), .ZN(\mult_22/ab[42][45] ) );
  NOR2_X1 U11673 ( .A1(n2662), .A2(n2979), .ZN(\mult_22/ab[40][47] ) );
  NOR2_X1 U11674 ( .A1(n2674), .A2(n2967), .ZN(\mult_22/ab[38][49] ) );
  NOR2_X1 U11675 ( .A1(n2687), .A2(n2955), .ZN(\mult_22/ab[36][51] ) );
  NOR2_X1 U11676 ( .A1(n2699), .A2(n2944), .ZN(\mult_22/ab[34][53] ) );
  NOR2_X1 U11677 ( .A1(n2709), .A2(n2932), .ZN(\mult_22/ab[32][55] ) );
  NOR2_X1 U11678 ( .A1(n2716), .A2(n2920), .ZN(\mult_22/ab[30][57] ) );
  NOR2_X1 U11679 ( .A1(n2728), .A2(n2908), .ZN(\mult_22/ab[28][59] ) );
  NOR2_X1 U11680 ( .A1(n2619), .A2(n3020), .ZN(\mult_22/ab[47][40] ) );
  NOR2_X1 U11681 ( .A1(n2632), .A2(n3009), .ZN(\mult_22/ab[45][42] ) );
  NOR2_X1 U11682 ( .A1(n2644), .A2(n2997), .ZN(\mult_22/ab[43][44] ) );
  NOR2_X1 U11683 ( .A1(n2656), .A2(n2985), .ZN(\mult_22/ab[41][46] ) );
  NOR2_X1 U11684 ( .A1(n2668), .A2(n2973), .ZN(\mult_22/ab[39][48] ) );
  NOR2_X1 U11685 ( .A1(n2680), .A2(n2961), .ZN(\mult_22/ab[37][50] ) );
  NOR2_X1 U11686 ( .A1(n2692), .A2(n2949), .ZN(\mult_22/ab[35][52] ) );
  NOR2_X1 U11687 ( .A1(n2712), .A2(n2926), .ZN(\mult_22/ab[31][56] ) );
  NOR2_X1 U11688 ( .A1(n2720), .A2(n2914), .ZN(\mult_22/ab[29][58] ) );
  NOR2_X1 U11689 ( .A1(n2732), .A2(n2902), .ZN(\mult_22/ab[27][60] ) );
  NOR2_X1 U11690 ( .A1(n2738), .A2(n2896), .ZN(\mult_22/ab[26][61] ) );
  NOR2_X1 U11691 ( .A1(n2590), .A2(n3056), .ZN(\mult_22/ab[53][35] ) );
  NOR2_X1 U11692 ( .A1(n2602), .A2(n3044), .ZN(\mult_22/ab[51][37] ) );
  NOR2_X1 U11693 ( .A1(n2590), .A2(n3074), .ZN(\mult_22/ab[56][35] ) );
  NOR2_X1 U11694 ( .A1(n2596), .A2(n3050), .ZN(\mult_22/ab[52][36] ) );
  NOR2_X1 U11695 ( .A1(n2608), .A2(n3038), .ZN(\mult_22/ab[50][38] ) );
  NOR2_X1 U11696 ( .A1(n2613), .A2(n3032), .ZN(\mult_22/ab[49][39] ) );
  NOR2_X1 U11697 ( .A1(n2627), .A2(n3020), .ZN(\mult_22/ab[47][41] ) );
  NOR2_X1 U11698 ( .A1(n2639), .A2(n3009), .ZN(\mult_22/ab[45][43] ) );
  NOR2_X1 U11699 ( .A1(n2650), .A2(n2997), .ZN(\mult_22/ab[43][45] ) );
  NOR2_X1 U11700 ( .A1(n2662), .A2(n2985), .ZN(\mult_22/ab[41][47] ) );
  NOR2_X1 U11701 ( .A1(n2674), .A2(n2973), .ZN(\mult_22/ab[39][49] ) );
  NOR2_X1 U11702 ( .A1(n2687), .A2(n2961), .ZN(\mult_22/ab[37][51] ) );
  NOR2_X1 U11703 ( .A1(n2696), .A2(n2950), .ZN(\mult_22/ab[35][53] ) );
  NOR2_X1 U11704 ( .A1(n2709), .A2(n2938), .ZN(\mult_22/ab[33][55] ) );
  NOR2_X1 U11705 ( .A1(n2716), .A2(n2926), .ZN(\mult_22/ab[31][57] ) );
  NOR2_X1 U11706 ( .A1(n2729), .A2(n2914), .ZN(\mult_22/ab[29][59] ) );
  NOR2_X1 U11707 ( .A1(n2619), .A2(n3026), .ZN(\mult_22/ab[48][40] ) );
  NOR2_X1 U11708 ( .A1(n2632), .A2(n3015), .ZN(\mult_22/ab[46][42] ) );
  NOR2_X1 U11709 ( .A1(n2644), .A2(n3003), .ZN(\mult_22/ab[44][44] ) );
  NOR2_X1 U11710 ( .A1(n2656), .A2(n2991), .ZN(\mult_22/ab[42][46] ) );
  NOR2_X1 U11711 ( .A1(n2668), .A2(n2979), .ZN(\mult_22/ab[40][48] ) );
  NOR2_X1 U11712 ( .A1(n2680), .A2(n2967), .ZN(\mult_22/ab[38][50] ) );
  NOR2_X1 U11713 ( .A1(n2692), .A2(n2955), .ZN(\mult_22/ab[36][52] ) );
  NOR2_X1 U11714 ( .A1(n2712), .A2(n2932), .ZN(\mult_22/ab[32][56] ) );
  NOR2_X1 U11715 ( .A1(n2720), .A2(n2920), .ZN(\mult_22/ab[30][58] ) );
  NOR2_X1 U11716 ( .A1(n2590), .A2(n3062), .ZN(\mult_22/ab[54][35] ) );
  NOR2_X1 U11717 ( .A1(n2732), .A2(n2908), .ZN(\mult_22/ab[28][60] ) );
  NOR2_X1 U11718 ( .A1(n2739), .A2(n2902), .ZN(\mult_22/ab[27][61] ) );
  NOR2_X1 U11719 ( .A1(n2596), .A2(n3056), .ZN(\mult_22/ab[53][36] ) );
  NOR2_X1 U11720 ( .A1(n2602), .A2(n3050), .ZN(\mult_22/ab[52][37] ) );
  NOR2_X1 U11721 ( .A1(n2608), .A2(n3044), .ZN(\mult_22/ab[51][38] ) );
  NOR2_X1 U11722 ( .A1(n2613), .A2(n3038), .ZN(\mult_22/ab[50][39] ) );
  NOR2_X1 U11723 ( .A1(n2627), .A2(n3026), .ZN(\mult_22/ab[48][41] ) );
  NOR2_X1 U11724 ( .A1(n2639), .A2(n3015), .ZN(\mult_22/ab[46][43] ) );
  NOR2_X1 U11725 ( .A1(n2651), .A2(n3003), .ZN(\mult_22/ab[44][45] ) );
  NOR2_X1 U11726 ( .A1(n2662), .A2(n2991), .ZN(\mult_22/ab[42][47] ) );
  NOR2_X1 U11727 ( .A1(n2674), .A2(n2979), .ZN(\mult_22/ab[40][49] ) );
  NOR2_X1 U11728 ( .A1(n2686), .A2(n2967), .ZN(\mult_22/ab[38][51] ) );
  NOR2_X1 U11729 ( .A1(n2619), .A2(n3032), .ZN(\mult_22/ab[49][40] ) );
  NOR2_X1 U11730 ( .A1(n2697), .A2(n2956), .ZN(\mult_22/ab[36][53] ) );
  NOR2_X1 U11731 ( .A1(n2632), .A2(n3021), .ZN(\mult_22/ab[47][42] ) );
  NOR2_X1 U11732 ( .A1(n2709), .A2(n2944), .ZN(\mult_22/ab[34][55] ) );
  NOR2_X1 U11733 ( .A1(n2644), .A2(n3009), .ZN(\mult_22/ab[45][44] ) );
  NOR2_X1 U11734 ( .A1(n2716), .A2(n2932), .ZN(\mult_22/ab[32][57] ) );
  NOR2_X1 U11735 ( .A1(n2656), .A2(n2997), .ZN(\mult_22/ab[43][46] ) );
  NOR2_X1 U11736 ( .A1(n2730), .A2(n2920), .ZN(\mult_22/ab[30][59] ) );
  NOR2_X1 U11737 ( .A1(n2668), .A2(n2985), .ZN(\mult_22/ab[41][48] ) );
  NOR2_X1 U11738 ( .A1(n2680), .A2(n2973), .ZN(\mult_22/ab[39][50] ) );
  NOR2_X1 U11739 ( .A1(n2692), .A2(n2961), .ZN(\mult_22/ab[37][52] ) );
  NOR2_X1 U11740 ( .A1(n2712), .A2(n2938), .ZN(\mult_22/ab[33][56] ) );
  NOR2_X1 U11741 ( .A1(n2720), .A2(n2926), .ZN(\mult_22/ab[31][58] ) );
  NOR2_X1 U11742 ( .A1(n2732), .A2(n2914), .ZN(\mult_22/ab[29][60] ) );
  NOR2_X1 U11743 ( .A1(n2740), .A2(n2908), .ZN(\mult_22/ab[28][61] ) );
  NOR2_X1 U11744 ( .A1(n2602), .A2(n3056), .ZN(\mult_22/ab[53][37] ) );
  NOR2_X1 U11745 ( .A1(n2596), .A2(n3062), .ZN(\mult_22/ab[54][36] ) );
  NOR2_X1 U11746 ( .A1(n2608), .A2(n3050), .ZN(\mult_22/ab[52][38] ) );
  NOR2_X1 U11747 ( .A1(n2613), .A2(n3044), .ZN(\mult_22/ab[51][39] ) );
  NOR2_X1 U11748 ( .A1(n2627), .A2(n3032), .ZN(\mult_22/ab[49][41] ) );
  NOR2_X1 U11749 ( .A1(n2639), .A2(n3021), .ZN(\mult_22/ab[47][43] ) );
  NOR2_X1 U11750 ( .A1(n2651), .A2(n3009), .ZN(\mult_22/ab[45][45] ) );
  NOR2_X1 U11751 ( .A1(n2662), .A2(n2997), .ZN(\mult_22/ab[43][47] ) );
  NOR2_X1 U11752 ( .A1(n2674), .A2(n2985), .ZN(\mult_22/ab[41][49] ) );
  NOR2_X1 U11753 ( .A1(n2686), .A2(n2973), .ZN(\mult_22/ab[39][51] ) );
  NOR2_X1 U11754 ( .A1(n2700), .A2(n2962), .ZN(\mult_22/ab[37][53] ) );
  NOR2_X1 U11755 ( .A1(n2709), .A2(n2950), .ZN(\mult_22/ab[35][55] ) );
  NOR2_X1 U11756 ( .A1(n2716), .A2(n2938), .ZN(\mult_22/ab[33][57] ) );
  NOR2_X1 U11757 ( .A1(n2725), .A2(n2926), .ZN(\mult_22/ab[31][59] ) );
  NOR2_X1 U11758 ( .A1(n2619), .A2(n3038), .ZN(\mult_22/ab[50][40] ) );
  NOR2_X1 U11759 ( .A1(n2631), .A2(n3027), .ZN(\mult_22/ab[48][42] ) );
  NOR2_X1 U11760 ( .A1(n2644), .A2(n3015), .ZN(\mult_22/ab[46][44] ) );
  NOR2_X1 U11761 ( .A1(n2656), .A2(n3003), .ZN(\mult_22/ab[44][46] ) );
  NOR2_X1 U11762 ( .A1(n2668), .A2(n2991), .ZN(\mult_22/ab[42][48] ) );
  NOR2_X1 U11763 ( .A1(n2680), .A2(n2979), .ZN(\mult_22/ab[40][50] ) );
  NOR2_X1 U11764 ( .A1(n2692), .A2(n2967), .ZN(\mult_22/ab[38][52] ) );
  NOR2_X1 U11765 ( .A1(n2702), .A2(n2956), .ZN(\mult_22/ab[36][54] ) );
  NOR2_X1 U11766 ( .A1(n2712), .A2(n2944), .ZN(\mult_22/ab[34][56] ) );
  NOR2_X1 U11767 ( .A1(n2720), .A2(n2932), .ZN(\mult_22/ab[32][58] ) );
  NOR2_X1 U11768 ( .A1(n2732), .A2(n2920), .ZN(\mult_22/ab[30][60] ) );
  NOR2_X1 U11769 ( .A1(n2738), .A2(n2914), .ZN(\mult_22/ab[29][61] ) );
  NOR2_X1 U11770 ( .A1(n2596), .A2(n3068), .ZN(\mult_22/ab[55][36] ) );
  NOR2_X1 U11771 ( .A1(n2602), .A2(n3062), .ZN(\mult_22/ab[54][37] ) );
  NOR2_X1 U11772 ( .A1(n2608), .A2(n3056), .ZN(\mult_22/ab[53][38] ) );
  NOR2_X1 U11773 ( .A1(n2613), .A2(n3050), .ZN(\mult_22/ab[52][39] ) );
  NOR2_X1 U11774 ( .A1(n2627), .A2(n3038), .ZN(\mult_22/ab[50][41] ) );
  NOR2_X1 U11775 ( .A1(n2639), .A2(n3027), .ZN(\mult_22/ab[48][43] ) );
  NOR2_X1 U11776 ( .A1(n2651), .A2(n3015), .ZN(\mult_22/ab[46][45] ) );
  NOR2_X1 U11777 ( .A1(n2662), .A2(n3003), .ZN(\mult_22/ab[44][47] ) );
  NOR2_X1 U11778 ( .A1(n2674), .A2(n2991), .ZN(\mult_22/ab[42][49] ) );
  NOR2_X1 U11779 ( .A1(n2686), .A2(n2979), .ZN(\mult_22/ab[40][51] ) );
  NOR2_X1 U11780 ( .A1(n2695), .A2(n2968), .ZN(\mult_22/ab[38][53] ) );
  NOR2_X1 U11781 ( .A1(n2709), .A2(n2956), .ZN(\mult_22/ab[36][55] ) );
  NOR2_X1 U11782 ( .A1(n2716), .A2(n2944), .ZN(\mult_22/ab[34][57] ) );
  NOR2_X1 U11783 ( .A1(n2726), .A2(n2932), .ZN(\mult_22/ab[32][59] ) );
  NOR2_X1 U11784 ( .A1(n2619), .A2(n3044), .ZN(\mult_22/ab[51][40] ) );
  NOR2_X1 U11785 ( .A1(n2631), .A2(n3033), .ZN(\mult_22/ab[49][42] ) );
  NOR2_X1 U11786 ( .A1(n2644), .A2(n3021), .ZN(\mult_22/ab[47][44] ) );
  NOR2_X1 U11787 ( .A1(n2656), .A2(n3009), .ZN(\mult_22/ab[45][46] ) );
  NOR2_X1 U11788 ( .A1(n2668), .A2(n2997), .ZN(\mult_22/ab[43][48] ) );
  NOR2_X1 U11789 ( .A1(n2680), .A2(n2985), .ZN(\mult_22/ab[41][50] ) );
  NOR2_X1 U11790 ( .A1(n2692), .A2(n2973), .ZN(\mult_22/ab[39][52] ) );
  NOR2_X1 U11791 ( .A1(n2702), .A2(n2962), .ZN(\mult_22/ab[37][54] ) );
  NOR2_X1 U11792 ( .A1(n2712), .A2(n2950), .ZN(\mult_22/ab[35][56] ) );
  NOR2_X1 U11793 ( .A1(n2721), .A2(n2938), .ZN(\mult_22/ab[33][58] ) );
  NOR2_X1 U11794 ( .A1(n2732), .A2(n2926), .ZN(\mult_22/ab[31][60] ) );
  NOR2_X1 U11795 ( .A1(n2741), .A2(n2920), .ZN(\mult_22/ab[30][61] ) );
  NOR2_X1 U11796 ( .A1(n2542), .A2(n2785), .ZN(\mult_22/ab[8][27] ) );
  NOR2_X1 U11797 ( .A1(n2535), .A2(n2797), .ZN(\mult_22/ab[10][25] ) );
  NOR2_X1 U11798 ( .A1(n2523), .A2(n2809), .ZN(\mult_22/ab[12][23] ) );
  NOR2_X1 U11799 ( .A1(n2510), .A2(n2821), .ZN(\mult_22/ab[14][21] ) );
  NOR2_X1 U11800 ( .A1(n2498), .A2(n2832), .ZN(\mult_22/ab[16][19] ) );
  NOR2_X1 U11801 ( .A1(n2486), .A2(n2844), .ZN(\mult_22/ab[18][17] ) );
  NOR2_X1 U11802 ( .A1(n2474), .A2(n2856), .ZN(\mult_22/ab[20][15] ) );
  NOR2_X1 U11803 ( .A1(n2462), .A2(n2868), .ZN(\mult_22/ab[22][13] ) );
  NOR2_X1 U11804 ( .A1(n2450), .A2(n2880), .ZN(\mult_22/ab[24][11] ) );
  NOR2_X1 U11805 ( .A1(n2437), .A2(n2897), .ZN(\mult_22/ab[26][9] ) );
  NOR2_X1 U11806 ( .A1(n2425), .A2(n2909), .ZN(\mult_22/ab[28][7] ) );
  NOR2_X1 U11807 ( .A1(n2413), .A2(n2920), .ZN(\mult_22/ab[30][5] ) );
  NOR2_X1 U11808 ( .A1(n2536), .A2(n2785), .ZN(\mult_22/ab[8][26] ) );
  NOR2_X1 U11809 ( .A1(n2524), .A2(n2797), .ZN(\mult_22/ab[10][24] ) );
  NOR2_X1 U11810 ( .A1(n2401), .A2(n2930), .ZN(\mult_22/ab[32][3] ) );
  NOR2_X1 U11811 ( .A1(n2517), .A2(n2809), .ZN(\mult_22/ab[12][22] ) );
  NOR2_X1 U11812 ( .A1(n2504), .A2(n2821), .ZN(\mult_22/ab[14][20] ) );
  NOR2_X1 U11813 ( .A1(n2492), .A2(n2832), .ZN(\mult_22/ab[16][18] ) );
  NOR2_X1 U11814 ( .A1(n2480), .A2(n2844), .ZN(\mult_22/ab[18][16] ) );
  NOR2_X1 U11815 ( .A1(n2468), .A2(n2856), .ZN(\mult_22/ab[20][14] ) );
  NOR2_X1 U11816 ( .A1(n2456), .A2(n2868), .ZN(\mult_22/ab[22][12] ) );
  NOR2_X1 U11817 ( .A1(n2441), .A2(n2880), .ZN(\mult_22/ab[24][10] ) );
  NOR2_X1 U11818 ( .A1(n2431), .A2(n2897), .ZN(\mult_22/ab[26][8] ) );
  NOR2_X1 U11819 ( .A1(n2419), .A2(n2908), .ZN(\mult_22/ab[28][6] ) );
  NOR2_X1 U11820 ( .A1(n2548), .A2(n2767), .ZN(\mult_22/ab[5][28] ) );
  NOR2_X1 U11821 ( .A1(n2405), .A2(n2919), .ZN(\mult_22/ab[30][4] ) );
  NOR2_X1 U11822 ( .A1(n2549), .A2(n2761), .ZN(\mult_22/ab[4][28] ) );
  NOR2_X1 U11823 ( .A1(n2388), .A2(n2976), .ZN(\mult_22/ab[40][1] ) );
  NOR2_X1 U11824 ( .A1(n2401), .A2(n2924), .ZN(\mult_22/ab[31][3] ) );
  NOR2_X1 U11825 ( .A1(n2542), .A2(n2773), .ZN(\mult_22/ab[6][27] ) );
  NOR2_X1 U11826 ( .A1(n2530), .A2(n2785), .ZN(\mult_22/ab[8][25] ) );
  NOR2_X1 U11827 ( .A1(n2523), .A2(n2797), .ZN(\mult_22/ab[10][23] ) );
  NOR2_X1 U11828 ( .A1(n2511), .A2(n2809), .ZN(\mult_22/ab[12][21] ) );
  NOR2_X1 U11829 ( .A1(n2498), .A2(n2820), .ZN(\mult_22/ab[14][19] ) );
  NOR2_X1 U11830 ( .A1(n2486), .A2(n2832), .ZN(\mult_22/ab[16][17] ) );
  NOR2_X1 U11831 ( .A1(n2474), .A2(n2844), .ZN(\mult_22/ab[18][15] ) );
  NOR2_X1 U11832 ( .A1(n2462), .A2(n2856), .ZN(\mult_22/ab[20][13] ) );
  NOR2_X1 U11833 ( .A1(n2450), .A2(n2868), .ZN(\mult_22/ab[22][11] ) );
  NOR2_X1 U11834 ( .A1(n2438), .A2(n2885), .ZN(\mult_22/ab[24][9] ) );
  NOR2_X1 U11835 ( .A1(n2425), .A2(n2897), .ZN(\mult_22/ab[26][7] ) );
  NOR2_X1 U11836 ( .A1(n2413), .A2(n2908), .ZN(\mult_22/ab[28][5] ) );
  NOR2_X1 U11837 ( .A1(n2388), .A2(n2970), .ZN(\mult_22/ab[39][1] ) );
  NOR2_X1 U11838 ( .A1(n2536), .A2(n2773), .ZN(\mult_22/ab[6][26] ) );
  NOR2_X1 U11839 ( .A1(n2529), .A2(n2785), .ZN(\mult_22/ab[8][24] ) );
  NOR2_X1 U11840 ( .A1(n2388), .A2(n2964), .ZN(\mult_22/ab[38][1] ) );
  NOR2_X1 U11841 ( .A1(n2517), .A2(n2797), .ZN(\mult_22/ab[10][22] ) );
  NOR2_X1 U11842 ( .A1(n2505), .A2(n2809), .ZN(\mult_22/ab[12][20] ) );
  NOR2_X1 U11843 ( .A1(n2492), .A2(n2820), .ZN(\mult_22/ab[14][18] ) );
  NOR2_X1 U11844 ( .A1(n2480), .A2(n2832), .ZN(\mult_22/ab[16][16] ) );
  NOR2_X1 U11845 ( .A1(n2468), .A2(n2844), .ZN(\mult_22/ab[18][14] ) );
  NOR2_X1 U11846 ( .A1(n2550), .A2(n2755), .ZN(\mult_22/ab[3][28] ) );
  NOR2_X1 U11847 ( .A1(n2456), .A2(n2856), .ZN(\mult_22/ab[20][12] ) );
  NOR2_X1 U11848 ( .A1(n2441), .A2(n2868), .ZN(\mult_22/ab[22][10] ) );
  NOR2_X1 U11849 ( .A1(n2432), .A2(n2885), .ZN(\mult_22/ab[24][8] ) );
  NOR2_X1 U11850 ( .A1(n2419), .A2(n2897), .ZN(\mult_22/ab[26][6] ) );
  NOR2_X1 U11851 ( .A1(n2401), .A2(n2918), .ZN(\mult_22/ab[30][3] ) );
  NOR2_X1 U11852 ( .A1(n2405), .A2(n2907), .ZN(\mult_22/ab[28][4] ) );
  NOR2_X1 U11853 ( .A1(n2543), .A2(n2761), .ZN(\mult_22/ab[4][27] ) );
  NOR2_X1 U11854 ( .A1(n2544), .A2(n2755), .ZN(\mult_22/ab[3][27] ) );
  NOR2_X1 U11855 ( .A1(n2530), .A2(n2773), .ZN(\mult_22/ab[6][25] ) );
  NOR2_X1 U11856 ( .A1(n2530), .A2(n2767), .ZN(\mult_22/ab[5][25] ) );
  NOR2_X1 U11857 ( .A1(n2518), .A2(n2785), .ZN(\mult_22/ab[8][23] ) );
  NOR2_X1 U11858 ( .A1(n2518), .A2(n2779), .ZN(\mult_22/ab[7][23] ) );
  NOR2_X1 U11859 ( .A1(n2511), .A2(n2797), .ZN(\mult_22/ab[10][21] ) );
  NOR2_X1 U11860 ( .A1(n2506), .A2(n2791), .ZN(\mult_22/ab[9][21] ) );
  NOR2_X1 U11861 ( .A1(n2499), .A2(n2808), .ZN(\mult_22/ab[12][19] ) );
  NOR2_X1 U11862 ( .A1(n2499), .A2(n2802), .ZN(\mult_22/ab[11][19] ) );
  NOR2_X1 U11863 ( .A1(n2486), .A2(n2820), .ZN(\mult_22/ab[14][17] ) );
  NOR2_X1 U11864 ( .A1(n2486), .A2(n2814), .ZN(\mult_22/ab[13][17] ) );
  NOR2_X1 U11865 ( .A1(n2474), .A2(n2832), .ZN(\mult_22/ab[16][15] ) );
  NOR2_X1 U11866 ( .A1(n2474), .A2(n2826), .ZN(\mult_22/ab[15][15] ) );
  NOR2_X1 U11867 ( .A1(n2462), .A2(n2844), .ZN(\mult_22/ab[18][13] ) );
  NOR2_X1 U11868 ( .A1(n2462), .A2(n2838), .ZN(\mult_22/ab[17][13] ) );
  NOR2_X1 U11869 ( .A1(n2450), .A2(n2856), .ZN(\mult_22/ab[20][11] ) );
  NOR2_X1 U11870 ( .A1(n2450), .A2(n2850), .ZN(\mult_22/ab[19][11] ) );
  NOR2_X1 U11871 ( .A1(n2438), .A2(n2873), .ZN(\mult_22/ab[22][9] ) );
  NOR2_X1 U11872 ( .A1(n2438), .A2(n2867), .ZN(\mult_22/ab[21][9] ) );
  NOR2_X1 U11873 ( .A1(n2426), .A2(n2885), .ZN(\mult_22/ab[24][7] ) );
  NOR2_X1 U11874 ( .A1(n2426), .A2(n2879), .ZN(\mult_22/ab[23][7] ) );
  NOR2_X1 U11875 ( .A1(n2413), .A2(n2896), .ZN(\mult_22/ab[26][5] ) );
  NOR2_X1 U11876 ( .A1(n2414), .A2(n2890), .ZN(\mult_22/ab[25][5] ) );
  NOR2_X1 U11877 ( .A1(n2395), .A2(n2935), .ZN(\mult_22/ab[33][2] ) );
  NOR2_X1 U11878 ( .A1(n2401), .A2(n2912), .ZN(\mult_22/ab[29][3] ) );
  NOR2_X1 U11879 ( .A1(n2388), .A2(n2958), .ZN(\mult_22/ab[37][1] ) );
  NOR2_X1 U11880 ( .A1(n2401), .A2(n2906), .ZN(\mult_22/ab[28][3] ) );
  NOR2_X1 U11881 ( .A1(n2401), .A2(n2900), .ZN(\mult_22/ab[27][3] ) );
  NOR2_X1 U11882 ( .A1(n2395), .A2(n2929), .ZN(\mult_22/ab[32][2] ) );
  NOR2_X1 U11883 ( .A1(n2389), .A2(n2952), .ZN(\mult_22/ab[36][1] ) );
  NOR2_X1 U11884 ( .A1(n2531), .A2(n2761), .ZN(\mult_22/ab[4][25] ) );
  NOR2_X1 U11885 ( .A1(n2518), .A2(n2773), .ZN(\mult_22/ab[6][23] ) );
  NOR2_X1 U11886 ( .A1(n2506), .A2(n2785), .ZN(\mult_22/ab[8][21] ) );
  NOR2_X1 U11887 ( .A1(n2499), .A2(n2796), .ZN(\mult_22/ab[10][19] ) );
  NOR2_X1 U11888 ( .A1(n2487), .A2(n2808), .ZN(\mult_22/ab[12][17] ) );
  NOR2_X1 U11889 ( .A1(n2474), .A2(n2820), .ZN(\mult_22/ab[14][15] ) );
  NOR2_X1 U11890 ( .A1(n2462), .A2(n2832), .ZN(\mult_22/ab[16][13] ) );
  NOR2_X1 U11891 ( .A1(n2450), .A2(n2844), .ZN(\mult_22/ab[18][11] ) );
  NOR2_X1 U11892 ( .A1(n2438), .A2(n2861), .ZN(\mult_22/ab[20][9] ) );
  NOR2_X1 U11893 ( .A1(n2426), .A2(n2873), .ZN(\mult_22/ab[22][7] ) );
  NOR2_X1 U11894 ( .A1(n2414), .A2(n2884), .ZN(\mult_22/ab[24][5] ) );
  NOR2_X1 U11895 ( .A1(n2532), .A2(n2755), .ZN(\mult_22/ab[3][25] ) );
  NOR2_X1 U11896 ( .A1(n2518), .A2(n2767), .ZN(\mult_22/ab[5][23] ) );
  NOR2_X1 U11897 ( .A1(n2506), .A2(n2779), .ZN(\mult_22/ab[7][21] ) );
  NOR2_X1 U11898 ( .A1(n2494), .A2(n2790), .ZN(\mult_22/ab[9][19] ) );
  NOR2_X1 U11899 ( .A1(n2487), .A2(n2802), .ZN(\mult_22/ab[11][17] ) );
  NOR2_X1 U11900 ( .A1(n2474), .A2(n2814), .ZN(\mult_22/ab[13][15] ) );
  NOR2_X1 U11901 ( .A1(n2462), .A2(n2826), .ZN(\mult_22/ab[15][13] ) );
  NOR2_X1 U11902 ( .A1(n2450), .A2(n2838), .ZN(\mult_22/ab[17][11] ) );
  NOR2_X1 U11903 ( .A1(n2438), .A2(n2855), .ZN(\mult_22/ab[19][9] ) );
  NOR2_X1 U11904 ( .A1(n2426), .A2(n2867), .ZN(\mult_22/ab[21][7] ) );
  NOR2_X1 U11905 ( .A1(n2414), .A2(n2878), .ZN(\mult_22/ab[23][5] ) );
  NOR2_X1 U11906 ( .A1(n2389), .A2(n2946), .ZN(\mult_22/ab[35][1] ) );
  NOR2_X1 U11907 ( .A1(n2401), .A2(n2894), .ZN(\mult_22/ab[26][3] ) );
  NOR2_X1 U11908 ( .A1(n2395), .A2(n2923), .ZN(\mult_22/ab[31][2] ) );
  NOR2_X1 U11909 ( .A1(n2401), .A2(n2888), .ZN(\mult_22/ab[25][3] ) );
  NOR2_X1 U11910 ( .A1(n2395), .A2(n2917), .ZN(\mult_22/ab[30][2] ) );
  NOR2_X1 U11911 ( .A1(n2519), .A2(n2761), .ZN(\mult_22/ab[4][23] ) );
  NOR2_X1 U11912 ( .A1(n2506), .A2(n2773), .ZN(\mult_22/ab[6][21] ) );
  NOR2_X1 U11913 ( .A1(n2494), .A2(n2784), .ZN(\mult_22/ab[8][19] ) );
  NOR2_X1 U11914 ( .A1(n2487), .A2(n2796), .ZN(\mult_22/ab[10][17] ) );
  NOR2_X1 U11915 ( .A1(n2389), .A2(n2940), .ZN(\mult_22/ab[34][1] ) );
  NOR2_X1 U11916 ( .A1(n2475), .A2(n2808), .ZN(\mult_22/ab[12][15] ) );
  NOR2_X1 U11917 ( .A1(n2462), .A2(n2820), .ZN(\mult_22/ab[14][13] ) );
  NOR2_X1 U11918 ( .A1(n2450), .A2(n2832), .ZN(\mult_22/ab[16][11] ) );
  NOR2_X1 U11919 ( .A1(n2438), .A2(n2849), .ZN(\mult_22/ab[18][9] ) );
  NOR2_X1 U11920 ( .A1(n2426), .A2(n2861), .ZN(\mult_22/ab[20][7] ) );
  NOR2_X1 U11921 ( .A1(n2414), .A2(n2872), .ZN(\mult_22/ab[22][5] ) );
  NOR2_X1 U11922 ( .A1(n2395), .A2(n2911), .ZN(\mult_22/ab[29][2] ) );
  NOR2_X1 U11923 ( .A1(n2395), .A2(n2905), .ZN(\mult_22/ab[28][2] ) );
  NOR2_X1 U11924 ( .A1(n2402), .A2(n2882), .ZN(\mult_22/ab[24][3] ) );
  NOR2_X1 U11925 ( .A1(n2389), .A2(n2934), .ZN(\mult_22/ab[33][1] ) );
  NOR2_X1 U11926 ( .A1(n2395), .A2(n2899), .ZN(\mult_22/ab[27][2] ) );
  NOR2_X1 U11927 ( .A1(n2520), .A2(n2755), .ZN(\mult_22/ab[3][23] ) );
  NOR2_X1 U11928 ( .A1(n2506), .A2(n2767), .ZN(\mult_22/ab[5][21] ) );
  NOR2_X1 U11929 ( .A1(n2494), .A2(n2778), .ZN(\mult_22/ab[7][19] ) );
  NOR2_X1 U11930 ( .A1(n2482), .A2(n2790), .ZN(\mult_22/ab[9][17] ) );
  NOR2_X1 U11931 ( .A1(n2475), .A2(n2802), .ZN(\mult_22/ab[11][15] ) );
  NOR2_X1 U11932 ( .A1(n2463), .A2(n2814), .ZN(\mult_22/ab[13][13] ) );
  NOR2_X1 U11933 ( .A1(n2450), .A2(n2826), .ZN(\mult_22/ab[15][11] ) );
  NOR2_X1 U11934 ( .A1(n2438), .A2(n2843), .ZN(\mult_22/ab[17][9] ) );
  NOR2_X1 U11935 ( .A1(n2426), .A2(n2855), .ZN(\mult_22/ab[19][7] ) );
  NOR2_X1 U11936 ( .A1(n2414), .A2(n2866), .ZN(\mult_22/ab[21][5] ) );
  NOR2_X1 U11937 ( .A1(n2395), .A2(n2893), .ZN(\mult_22/ab[26][2] ) );
  NOR2_X1 U11938 ( .A1(n2389), .A2(n2928), .ZN(\mult_22/ab[32][1] ) );
  NOR2_X1 U11939 ( .A1(n2514), .A2(n2755), .ZN(\mult_22/ab[3][22] ) );
  NOR2_X1 U11940 ( .A1(n2500), .A2(n2767), .ZN(\mult_22/ab[5][20] ) );
  NOR2_X1 U11941 ( .A1(n2501), .A2(n2761), .ZN(\mult_22/ab[4][20] ) );
  NOR2_X1 U11942 ( .A1(n2488), .A2(n2778), .ZN(\mult_22/ab[7][18] ) );
  NOR2_X1 U11943 ( .A1(n2488), .A2(n2772), .ZN(\mult_22/ab[6][18] ) );
  NOR2_X1 U11944 ( .A1(n2476), .A2(n2790), .ZN(\mult_22/ab[9][16] ) );
  NOR2_X1 U11945 ( .A1(n2476), .A2(n2784), .ZN(\mult_22/ab[8][16] ) );
  NOR2_X1 U11946 ( .A1(n2469), .A2(n2802), .ZN(\mult_22/ab[11][14] ) );
  NOR2_X1 U11947 ( .A1(n2469), .A2(n2796), .ZN(\mult_22/ab[10][14] ) );
  NOR2_X1 U11948 ( .A1(n2402), .A2(n2876), .ZN(\mult_22/ab[23][3] ) );
  NOR2_X1 U11949 ( .A1(n2456), .A2(n2814), .ZN(\mult_22/ab[13][12] ) );
  NOR2_X1 U11950 ( .A1(n2457), .A2(n2808), .ZN(\mult_22/ab[12][12] ) );
  NOR2_X1 U11951 ( .A1(n2440), .A2(n2826), .ZN(\mult_22/ab[15][10] ) );
  NOR2_X1 U11952 ( .A1(n2440), .A2(n2820), .ZN(\mult_22/ab[14][10] ) );
  NOR2_X1 U11953 ( .A1(n2432), .A2(n2843), .ZN(\mult_22/ab[17][8] ) );
  NOR2_X1 U11954 ( .A1(n2432), .A2(n2837), .ZN(\mult_22/ab[16][8] ) );
  NOR2_X1 U11955 ( .A1(n2420), .A2(n2855), .ZN(\mult_22/ab[19][6] ) );
  NOR2_X1 U11956 ( .A1(n2420), .A2(n2848), .ZN(\mult_22/ab[18][6] ) );
  NOR2_X1 U11957 ( .A1(n2389), .A2(n2922), .ZN(\mult_22/ab[31][1] ) );
  NOR2_X1 U11958 ( .A1(n2404), .A2(n2865), .ZN(\mult_22/ab[21][4] ) );
  NOR2_X1 U11959 ( .A1(n2404), .A2(n2859), .ZN(\mult_22/ab[20][4] ) );
  NOR2_X1 U11960 ( .A1(n2389), .A2(n2916), .ZN(\mult_22/ab[30][1] ) );
  NOR2_X1 U11961 ( .A1(n2389), .A2(n2910), .ZN(\mult_22/ab[29][1] ) );
  NOR2_X1 U11962 ( .A1(n2402), .A2(n2870), .ZN(\mult_22/ab[22][3] ) );
  NOR2_X1 U11963 ( .A1(n2395), .A2(n2887), .ZN(\mult_22/ab[25][2] ) );
  NOR2_X1 U11964 ( .A1(n2402), .A2(n2864), .ZN(\mult_22/ab[21][3] ) );
  NOR2_X1 U11965 ( .A1(n2495), .A2(n2760), .ZN(\mult_22/ab[4][19] ) );
  NOR2_X1 U11966 ( .A1(n2482), .A2(n2772), .ZN(\mult_22/ab[6][17] ) );
  NOR2_X1 U11967 ( .A1(n2470), .A2(n2784), .ZN(\mult_22/ab[8][15] ) );
  NOR2_X1 U11968 ( .A1(n2463), .A2(n2796), .ZN(\mult_22/ab[10][13] ) );
  NOR2_X1 U11969 ( .A1(n2451), .A2(n2808), .ZN(\mult_22/ab[12][11] ) );
  NOR2_X1 U11970 ( .A1(n2438), .A2(n2825), .ZN(\mult_22/ab[14][9] ) );
  NOR2_X1 U11971 ( .A1(n2426), .A2(n2837), .ZN(\mult_22/ab[16][7] ) );
  NOR2_X1 U11972 ( .A1(n2414), .A2(n2848), .ZN(\mult_22/ab[18][5] ) );
  NOR2_X1 U11973 ( .A1(n2402), .A2(n2858), .ZN(\mult_22/ab[20][3] ) );
  NOR2_X1 U11974 ( .A1(n2489), .A2(n2760), .ZN(\mult_22/ab[4][18] ) );
  NOR2_X1 U11975 ( .A1(n2476), .A2(n2772), .ZN(\mult_22/ab[6][16] ) );
  NOR2_X1 U11976 ( .A1(n2464), .A2(n2784), .ZN(\mult_22/ab[8][14] ) );
  NOR2_X1 U11977 ( .A1(n2389), .A2(n2904), .ZN(\mult_22/ab[28][1] ) );
  NOR2_X1 U11978 ( .A1(n2457), .A2(n2796), .ZN(\mult_22/ab[10][12] ) );
  NOR2_X1 U11979 ( .A1(n2440), .A2(n2808), .ZN(\mult_22/ab[12][10] ) );
  NOR2_X1 U11980 ( .A1(n2432), .A2(n2825), .ZN(\mult_22/ab[14][8] ) );
  NOR2_X1 U11981 ( .A1(n2420), .A2(n2837), .ZN(\mult_22/ab[16][6] ) );
  NOR2_X1 U11982 ( .A1(n2404), .A2(n2847), .ZN(\mult_22/ab[18][4] ) );
  NOR2_X1 U11983 ( .A1(n2396), .A2(n2881), .ZN(\mult_22/ab[24][2] ) );
  NOR2_X1 U11984 ( .A1(n2389), .A2(n2898), .ZN(\mult_22/ab[27][1] ) );
  NOR2_X1 U11985 ( .A1(n2402), .A2(n2852), .ZN(\mult_22/ab[19][3] ) );
  NOR2_X1 U11986 ( .A1(n2483), .A2(n2760), .ZN(\mult_22/ab[4][17] ) );
  NOR2_X1 U11987 ( .A1(n2470), .A2(n2772), .ZN(\mult_22/ab[6][15] ) );
  NOR2_X1 U11988 ( .A1(n2458), .A2(n2784), .ZN(\mult_22/ab[8][13] ) );
  NOR2_X1 U11989 ( .A1(n2451), .A2(n2796), .ZN(\mult_22/ab[10][11] ) );
  NOR2_X1 U11990 ( .A1(n2439), .A2(n2813), .ZN(\mult_22/ab[12][9] ) );
  NOR2_X1 U11991 ( .A1(n2426), .A2(n2825), .ZN(\mult_22/ab[14][7] ) );
  NOR2_X1 U11992 ( .A1(n2414), .A2(n2836), .ZN(\mult_22/ab[16][5] ) );
  NOR2_X1 U11993 ( .A1(n2396), .A2(n2875), .ZN(\mult_22/ab[23][2] ) );
  NOR2_X1 U11994 ( .A1(n2396), .A2(n2869), .ZN(\mult_22/ab[22][2] ) );
  NOR2_X1 U11995 ( .A1(n2389), .A2(n2893), .ZN(\mult_22/ab[26][1] ) );
  NOR2_X1 U11996 ( .A1(n2402), .A2(n2846), .ZN(\mult_22/ab[18][3] ) );
  NOR2_X1 U11997 ( .A1(n2477), .A2(n2760), .ZN(\mult_22/ab[4][16] ) );
  NOR2_X1 U11998 ( .A1(n2464), .A2(n2772), .ZN(\mult_22/ab[6][14] ) );
  NOR2_X1 U11999 ( .A1(n2396), .A2(n2863), .ZN(\mult_22/ab[21][2] ) );
  NOR2_X1 U12000 ( .A1(n2452), .A2(n2784), .ZN(\mult_22/ab[8][12] ) );
  NOR2_X1 U12001 ( .A1(n2440), .A2(n2796), .ZN(\mult_22/ab[10][10] ) );
  NOR2_X1 U12002 ( .A1(n2433), .A2(n2813), .ZN(\mult_22/ab[12][8] ) );
  NOR2_X1 U12003 ( .A1(n2420), .A2(n2825), .ZN(\mult_22/ab[14][6] ) );
  NOR2_X1 U12004 ( .A1(n2404), .A2(n2835), .ZN(\mult_22/ab[16][4] ) );
  NOR2_X1 U12005 ( .A1(n2402), .A2(n2840), .ZN(\mult_22/ab[17][3] ) );
  NOR2_X1 U12006 ( .A1(n2396), .A2(n2857), .ZN(\mult_22/ab[20][2] ) );
  NOR2_X1 U12007 ( .A1(n2390), .A2(n2886), .ZN(\mult_22/ab[25][1] ) );
  NOR2_X1 U12008 ( .A1(n2471), .A2(n2760), .ZN(\mult_22/ab[4][15] ) );
  NOR2_X1 U12009 ( .A1(n2458), .A2(n2772), .ZN(\mult_22/ab[6][13] ) );
  NOR2_X1 U12010 ( .A1(n2446), .A2(n2784), .ZN(\mult_22/ab[8][11] ) );
  NOR2_X1 U12011 ( .A1(n2439), .A2(n2801), .ZN(\mult_22/ab[10][9] ) );
  NOR2_X1 U12012 ( .A1(n2427), .A2(n2813), .ZN(\mult_22/ab[12][7] ) );
  NOR2_X1 U12013 ( .A1(n2414), .A2(n2824), .ZN(\mult_22/ab[14][5] ) );
  NOR2_X1 U12014 ( .A1(n2472), .A2(n2754), .ZN(\mult_22/ab[3][15] ) );
  NOR2_X1 U12015 ( .A1(n2458), .A2(n2766), .ZN(\mult_22/ab[5][13] ) );
  NOR2_X1 U12016 ( .A1(n2446), .A2(n2778), .ZN(\mult_22/ab[7][11] ) );
  NOR2_X1 U12017 ( .A1(n2434), .A2(n2795), .ZN(\mult_22/ab[9][9] ) );
  NOR2_X1 U12018 ( .A1(n2459), .A2(n2760), .ZN(\mult_22/ab[4][13] ) );
  NOR2_X1 U12019 ( .A1(n2427), .A2(n2807), .ZN(\mult_22/ab[11][7] ) );
  NOR2_X1 U12020 ( .A1(n2446), .A2(n2772), .ZN(\mult_22/ab[6][11] ) );
  NOR2_X1 U12021 ( .A1(n2415), .A2(n2818), .ZN(\mult_22/ab[13][5] ) );
  NOR2_X1 U12022 ( .A1(n2434), .A2(n2789), .ZN(\mult_22/ab[8][9] ) );
  NOR2_X1 U12023 ( .A1(n2427), .A2(n2801), .ZN(\mult_22/ab[10][7] ) );
  NOR2_X1 U12024 ( .A1(n2415), .A2(n2812), .ZN(\mult_22/ab[12][5] ) );
  NOR2_X1 U12025 ( .A1(n2390), .A2(n2880), .ZN(\mult_22/ab[24][1] ) );
  NOR2_X1 U12026 ( .A1(n2396), .A2(n2851), .ZN(\mult_22/ab[19][2] ) );
  NOR2_X1 U12027 ( .A1(n2402), .A2(n2834), .ZN(\mult_22/ab[16][3] ) );
  NOR2_X1 U12028 ( .A1(n2390), .A2(n2874), .ZN(\mult_22/ab[23][1] ) );
  NOR2_X1 U12029 ( .A1(n2402), .A2(n2828), .ZN(\mult_22/ab[15][3] ) );
  NOR2_X1 U12030 ( .A1(n2402), .A2(n2822), .ZN(\mult_22/ab[14][3] ) );
  NOR2_X1 U12031 ( .A1(n2390), .A2(n2868), .ZN(\mult_22/ab[22][1] ) );
  NOR2_X1 U12032 ( .A1(n2396), .A2(n2845), .ZN(\mult_22/ab[18][2] ) );
  NOR2_X1 U12033 ( .A1(n2453), .A2(n2760), .ZN(\mult_22/ab[4][12] ) );
  NOR2_X1 U12034 ( .A1(n2444), .A2(n2772), .ZN(\mult_22/ab[6][10] ) );
  NOR2_X1 U12035 ( .A1(n2428), .A2(n2789), .ZN(\mult_22/ab[8][8] ) );
  NOR2_X1 U12036 ( .A1(n2421), .A2(n2801), .ZN(\mult_22/ab[10][6] ) );
  NOR2_X1 U12037 ( .A1(n2404), .A2(n2811), .ZN(\mult_22/ab[12][4] ) );
  NOR2_X1 U12038 ( .A1(n2390), .A2(n2863), .ZN(\mult_22/ab[21][1] ) );
  NOR2_X1 U12039 ( .A1(n2402), .A2(n2816), .ZN(\mult_22/ab[13][3] ) );
  NOR2_X1 U12040 ( .A1(n2447), .A2(n2760), .ZN(\mult_22/ab[4][11] ) );
  NOR2_X1 U12041 ( .A1(n2434), .A2(n2777), .ZN(\mult_22/ab[6][9] ) );
  NOR2_X1 U12042 ( .A1(n2422), .A2(n2789), .ZN(\mult_22/ab[8][7] ) );
  NOR2_X1 U12043 ( .A1(n2415), .A2(n2800), .ZN(\mult_22/ab[10][5] ) );
  NOR2_X1 U12044 ( .A1(n2448), .A2(n2754), .ZN(\mult_22/ab[3][11] ) );
  NOR2_X1 U12045 ( .A1(n2434), .A2(n2771), .ZN(\mult_22/ab[5][9] ) );
  NOR2_X1 U12046 ( .A1(n2422), .A2(n2783), .ZN(\mult_22/ab[7][7] ) );
  NOR2_X1 U12047 ( .A1(n2410), .A2(n2794), .ZN(\mult_22/ab[9][5] ) );
  NOR2_X1 U12048 ( .A1(n2396), .A2(n2839), .ZN(\mult_22/ab[17][2] ) );
  NOR2_X1 U12049 ( .A1(n2403), .A2(n2810), .ZN(\mult_22/ab[12][3] ) );
  NOR2_X1 U12050 ( .A1(n2396), .A2(n2833), .ZN(\mult_22/ab[16][2] ) );
  NOR2_X1 U12051 ( .A1(n2435), .A2(n2765), .ZN(\mult_22/ab[4][9] ) );
  NOR2_X1 U12052 ( .A1(n2422), .A2(n2777), .ZN(\mult_22/ab[6][7] ) );
  NOR2_X1 U12053 ( .A1(n2410), .A2(n2788), .ZN(\mult_22/ab[8][5] ) );
  NOR2_X1 U12054 ( .A1(n2396), .A2(n2827), .ZN(\mult_22/ab[15][2] ) );
  NOR2_X1 U12055 ( .A1(n2403), .A2(n2804), .ZN(\mult_22/ab[11][3] ) );
  NOR2_X1 U12056 ( .A1(n2390), .A2(n2856), .ZN(\mult_22/ab[20][1] ) );
  NOR2_X1 U12057 ( .A1(n2403), .A2(n2798), .ZN(\mult_22/ab[10][3] ) );
  NOR2_X1 U12058 ( .A1(n2436), .A2(n2759), .ZN(\mult_22/ab[3][9] ) );
  NOR2_X1 U12059 ( .A1(n2422), .A2(n2771), .ZN(\mult_22/ab[5][7] ) );
  NOR2_X1 U12060 ( .A1(n2410), .A2(n2782), .ZN(\mult_22/ab[7][5] ) );
  NOR2_X1 U12061 ( .A1(n2390), .A2(n2850), .ZN(\mult_22/ab[19][1] ) );
  NOR2_X1 U12062 ( .A1(n2396), .A2(n2821), .ZN(\mult_22/ab[14][2] ) );
  NOR2_X1 U12063 ( .A1(n2398), .A2(n2792), .ZN(\mult_22/ab[9][3] ) );
  NOR2_X1 U12064 ( .A1(n2396), .A2(n2815), .ZN(\mult_22/ab[13][2] ) );
  NOR2_X1 U12065 ( .A1(n2423), .A2(n2765), .ZN(\mult_22/ab[4][7] ) );
  NOR2_X1 U12066 ( .A1(n2410), .A2(n2776), .ZN(\mult_22/ab[6][5] ) );
  NOR2_X1 U12067 ( .A1(n2397), .A2(n2809), .ZN(\mult_22/ab[12][2] ) );
  NOR2_X1 U12068 ( .A1(n2390), .A2(n2844), .ZN(\mult_22/ab[18][1] ) );
  NOR2_X1 U12069 ( .A1(n2398), .A2(n2786), .ZN(\mult_22/ab[8][3] ) );
  NOR2_X1 U12070 ( .A1(n2390), .A2(n2838), .ZN(\mult_22/ab[17][1] ) );
  NOR2_X1 U12071 ( .A1(n2417), .A2(n2764), .ZN(\mult_22/ab[4][6] ) );
  NOR2_X1 U12072 ( .A1(n2390), .A2(n2832), .ZN(\mult_22/ab[16][1] ) );
  NOR2_X1 U12073 ( .A1(n2397), .A2(n2803), .ZN(\mult_22/ab[11][2] ) );
  NOR2_X1 U12074 ( .A1(n2408), .A2(n2775), .ZN(\mult_22/ab[6][4] ) );
  NOR2_X1 U12075 ( .A1(n2398), .A2(n2780), .ZN(\mult_22/ab[7][3] ) );
  NOR2_X1 U12076 ( .A1(n2418), .A2(n2758), .ZN(\mult_22/ab[3][6] ) );
  NOR2_X1 U12077 ( .A1(n2397), .A2(n2797), .ZN(\mult_22/ab[10][2] ) );
  NOR2_X1 U12078 ( .A1(n2408), .A2(n2769), .ZN(\mult_22/ab[5][4] ) );
  NOR2_X1 U12079 ( .A1(n2407), .A2(n2763), .ZN(\mult_22/ab[4][4] ) );
  NOR2_X1 U12080 ( .A1(n2390), .A2(n2826), .ZN(\mult_22/ab[15][1] ) );
  NOR2_X1 U12081 ( .A1(n2398), .A2(n2774), .ZN(\mult_22/ab[6][3] ) );
  NOR2_X1 U12082 ( .A1(n2398), .A2(n2768), .ZN(\mult_22/ab[5][3] ) );
  NOR2_X1 U12083 ( .A1(n2390), .A2(n2820), .ZN(\mult_22/ab[14][1] ) );
  NOR2_X1 U12084 ( .A1(n2392), .A2(n2791), .ZN(\mult_22/ab[9][2] ) );
  NOR2_X1 U12085 ( .A1(n2391), .A2(n2814), .ZN(\mult_22/ab[13][1] ) );
  NOR2_X1 U12086 ( .A1(n2392), .A2(n2785), .ZN(\mult_22/ab[8][2] ) );
  NOR2_X1 U12087 ( .A1(n2391), .A2(n2808), .ZN(\mult_22/ab[12][1] ) );
  NOR2_X1 U12088 ( .A1(n2399), .A2(n2762), .ZN(\mult_22/ab[4][3] ) );
  NOR2_X1 U12089 ( .A1(n2400), .A2(n2756), .ZN(\mult_22/ab[3][3] ) );
  NOR2_X1 U12090 ( .A1(n2391), .A2(n2802), .ZN(\mult_22/ab[11][1] ) );
  NOR2_X1 U12091 ( .A1(n2392), .A2(n2779), .ZN(\mult_22/ab[7][2] ) );
  NOR2_X1 U12092 ( .A1(n2392), .A2(n2773), .ZN(\mult_22/ab[6][2] ) );
  NOR2_X1 U12093 ( .A1(n2391), .A2(n2796), .ZN(\mult_22/ab[10][1] ) );
  NOR2_X1 U12094 ( .A1(n2392), .A2(n2767), .ZN(\mult_22/ab[5][2] ) );
  NOR2_X1 U12095 ( .A1(n2386), .A2(n2790), .ZN(\mult_22/ab[9][1] ) );
  NOR2_X1 U12096 ( .A1(n2393), .A2(n2761), .ZN(\mult_22/ab[4][2] ) );
  NOR2_X1 U12097 ( .A1(n2394), .A2(n2755), .ZN(\mult_22/ab[3][2] ) );
  NOR2_X1 U12098 ( .A1(n2386), .A2(n2784), .ZN(\mult_22/ab[8][1] ) );
  NOR2_X1 U12099 ( .A1(n2386), .A2(n2778), .ZN(\mult_22/ab[7][1] ) );
  NOR2_X1 U12100 ( .A1(n2386), .A2(n2772), .ZN(\mult_22/ab[6][1] ) );
  NOR2_X1 U12101 ( .A1(n2386), .A2(n2766), .ZN(\mult_22/ab[5][1] ) );
  NOR2_X1 U12102 ( .A1(n2387), .A2(n2760), .ZN(\mult_22/ab[4][1] ) );
  NOR2_X1 U12103 ( .A1(n2388), .A2(n2754), .ZN(\mult_22/ab[3][1] ) );
  NOR2_X1 U12104 ( .A1(n2384), .A2(n3066), .ZN(\mult_22/ab[55][0] ) );
  NOR2_X1 U12105 ( .A1(n2384), .A2(n3060), .ZN(\mult_22/ab[54][0] ) );
  NOR2_X1 U12106 ( .A1(n2383), .A2(n3054), .ZN(\mult_22/ab[53][0] ) );
  NOR2_X1 U12107 ( .A1(n2383), .A2(n3048), .ZN(\mult_22/ab[52][0] ) );
  NOR2_X1 U12108 ( .A1(n2383), .A2(n3042), .ZN(\mult_22/ab[51][0] ) );
  NOR2_X1 U12109 ( .A1(n2383), .A2(n3036), .ZN(\mult_22/ab[50][0] ) );
  NOR2_X1 U12110 ( .A1(n2383), .A2(n3030), .ZN(\mult_22/ab[49][0] ) );
  NOR2_X1 U12111 ( .A1(n2383), .A2(n3024), .ZN(\mult_22/ab[48][0] ) );
  NOR2_X1 U12112 ( .A1(n2383), .A2(n3018), .ZN(\mult_22/ab[47][0] ) );
  NOR2_X1 U12113 ( .A1(n2383), .A2(n3012), .ZN(\mult_22/ab[46][0] ) );
  NOR2_X1 U12114 ( .A1(n2383), .A2(n3006), .ZN(\mult_22/ab[45][0] ) );
  NOR2_X1 U12115 ( .A1(n2383), .A2(n3000), .ZN(\mult_22/ab[44][0] ) );
  NOR2_X1 U12116 ( .A1(n2383), .A2(n2994), .ZN(\mult_22/ab[43][0] ) );
  NOR2_X1 U12117 ( .A1(n2382), .A2(n2988), .ZN(\mult_22/ab[42][0] ) );
  NOR2_X1 U12118 ( .A1(n2382), .A2(n2982), .ZN(\mult_22/ab[41][0] ) );
  NOR2_X1 U12119 ( .A1(n2382), .A2(n2976), .ZN(\mult_22/ab[40][0] ) );
  NOR2_X1 U12120 ( .A1(n2382), .A2(n2970), .ZN(\mult_22/ab[39][0] ) );
  NOR2_X1 U12121 ( .A1(n2382), .A2(n2964), .ZN(\mult_22/ab[38][0] ) );
  NOR2_X1 U12122 ( .A1(n2382), .A2(n2958), .ZN(\mult_22/ab[37][0] ) );
  NOR2_X1 U12123 ( .A1(n2382), .A2(n2952), .ZN(\mult_22/ab[36][0] ) );
  NOR2_X1 U12124 ( .A1(n2382), .A2(n2946), .ZN(\mult_22/ab[35][0] ) );
  NOR2_X1 U12125 ( .A1(n2382), .A2(n2940), .ZN(\mult_22/ab[34][0] ) );
  NOR2_X1 U12126 ( .A1(n2382), .A2(n2934), .ZN(\mult_22/ab[33][0] ) );
  NOR2_X1 U12127 ( .A1(n2382), .A2(n2928), .ZN(\mult_22/ab[32][0] ) );
  NOR2_X1 U12128 ( .A1(n2381), .A2(n2922), .ZN(\mult_22/ab[31][0] ) );
  NOR2_X1 U12129 ( .A1(n2381), .A2(n2916), .ZN(\mult_22/ab[30][0] ) );
  NOR2_X1 U12130 ( .A1(n2381), .A2(n2910), .ZN(\mult_22/ab[29][0] ) );
  NOR2_X1 U12131 ( .A1(n2381), .A2(n2904), .ZN(\mult_22/ab[28][0] ) );
  NOR2_X1 U12132 ( .A1(n2381), .A2(n2898), .ZN(\mult_22/ab[27][0] ) );
  NOR2_X1 U12133 ( .A1(n2381), .A2(n2892), .ZN(\mult_22/ab[26][0] ) );
  NOR2_X1 U12134 ( .A1(n2381), .A2(n2886), .ZN(\mult_22/ab[25][0] ) );
  NOR2_X1 U12135 ( .A1(n2381), .A2(n2880), .ZN(\mult_22/ab[24][0] ) );
  NOR2_X1 U12136 ( .A1(n2381), .A2(n2874), .ZN(\mult_22/ab[23][0] ) );
  NOR2_X1 U12137 ( .A1(n2381), .A2(n2868), .ZN(\mult_22/ab[22][0] ) );
  NOR2_X1 U12138 ( .A1(n2381), .A2(n2862), .ZN(\mult_22/ab[21][0] ) );
  NOR2_X1 U12139 ( .A1(n2380), .A2(n2856), .ZN(\mult_22/ab[20][0] ) );
  NOR2_X1 U12140 ( .A1(n2380), .A2(n2850), .ZN(\mult_22/ab[19][0] ) );
  NOR2_X1 U12141 ( .A1(n2380), .A2(n2844), .ZN(\mult_22/ab[18][0] ) );
  NOR2_X1 U12142 ( .A1(n2380), .A2(n2838), .ZN(\mult_22/ab[17][0] ) );
  NOR2_X1 U12143 ( .A1(n2380), .A2(n2832), .ZN(\mult_22/ab[16][0] ) );
  NOR2_X1 U12144 ( .A1(n2380), .A2(n2826), .ZN(\mult_22/ab[15][0] ) );
  NOR2_X1 U12145 ( .A1(n2380), .A2(n2820), .ZN(\mult_22/ab[14][0] ) );
  NOR2_X1 U12146 ( .A1(n2380), .A2(n2814), .ZN(\mult_22/ab[13][0] ) );
  NOR2_X1 U12147 ( .A1(n2380), .A2(n2808), .ZN(\mult_22/ab[12][0] ) );
  NOR2_X1 U12148 ( .A1(n2380), .A2(n2802), .ZN(\mult_22/ab[11][0] ) );
  NOR2_X1 U12149 ( .A1(n2380), .A2(n2796), .ZN(\mult_22/ab[10][0] ) );
  NOR2_X1 U12150 ( .A1(n2385), .A2(n2790), .ZN(\mult_22/ab[9][0] ) );
  NOR2_X1 U12151 ( .A1(n2385), .A2(n2784), .ZN(\mult_22/ab[8][0] ) );
  NOR2_X1 U12152 ( .A1(n2385), .A2(n2778), .ZN(\mult_22/ab[7][0] ) );
  NOR2_X1 U12153 ( .A1(n2384), .A2(n2772), .ZN(\mult_22/ab[6][0] ) );
  NOR2_X1 U12154 ( .A1(n2384), .A2(n2766), .ZN(\mult_22/ab[5][0] ) );
  NOR2_X1 U12155 ( .A1(n2383), .A2(n2760), .ZN(\mult_22/ab[4][0] ) );
  NOR2_X1 U12156 ( .A1(n2382), .A2(n2754), .ZN(\mult_22/ab[3][0] ) );
  NOR2_X1 U12157 ( .A1(n2560), .A2(n3115), .ZN(\mult_22/ab[63][30] ) );
  AOI21_X1 U12158 ( .B1(\mult_22/CARRYB[63][53] ), .B2(\mult_22/SUMB[63][54] ), 
        .A(n1330), .ZN(n1327) );
  NOR2_X1 U12159 ( .A1(n2723), .A2(n3118), .ZN(\mult_22/ab[63][58] ) );
  AOI21_X1 U12160 ( .B1(\mult_22/CARRYB[63][52] ), .B2(\mult_22/SUMB[63][53] ), 
        .A(n1338), .ZN(n1331) );
  AOI21_X1 U12161 ( .B1(\mult_22/CARRYB[63][54] ), .B2(\mult_22/SUMB[63][55] ), 
        .A(n1328), .ZN(n1321) );
  NOR2_X1 U12162 ( .A1(n2642), .A2(n3117), .ZN(\mult_22/ab[63][44] ) );
  NOR2_X1 U12163 ( .A1(n2666), .A2(n3117), .ZN(\mult_22/ab[63][48] ) );
  NOR2_X1 U12164 ( .A1(n2654), .A2(n3117), .ZN(\mult_22/ab[63][46] ) );
  NOR2_X1 U12165 ( .A1(n2618), .A2(n3116), .ZN(\mult_22/ab[63][40] ) );
  NOR2_X1 U12166 ( .A1(n2576), .A2(n3116), .ZN(\mult_22/ab[63][32] ) );
  NOR2_X1 U12167 ( .A1(n2694), .A2(n3117), .ZN(\mult_22/ab[63][52] ) );
  NOR2_X1 U12168 ( .A1(n2712), .A2(n3118), .ZN(\mult_22/ab[63][56] ) );
  NOR2_X1 U12169 ( .A1(n2735), .A2(n3118), .ZN(\mult_22/ab[63][60] ) );
  NOR2_X1 U12170 ( .A1(n2660), .A2(n3117), .ZN(\mult_22/ab[63][47] ) );
  NOR2_X1 U12171 ( .A1(n2607), .A2(n3116), .ZN(\mult_22/ab[63][38] ) );
  NOR2_X1 U12172 ( .A1(n2612), .A2(n3116), .ZN(\mult_22/ab[63][39] ) );
  NOR2_X1 U12173 ( .A1(n2601), .A2(n3116), .ZN(\mult_22/ab[63][37] ) );
  NOR2_X1 U12174 ( .A1(n2652), .A2(n3117), .ZN(\mult_22/ab[63][45] ) );
  NOR2_X1 U12175 ( .A1(n2640), .A2(n3117), .ZN(\mult_22/ab[63][43] ) );
  NOR2_X1 U12176 ( .A1(n2630), .A2(n3117), .ZN(\mult_22/ab[63][42] ) );
  NOR2_X1 U12177 ( .A1(n2589), .A2(n3116), .ZN(\mult_22/ab[63][35] ) );
  NOR2_X1 U12178 ( .A1(n2628), .A2(n3116), .ZN(\mult_22/ab[63][41] ) );
  NOR2_X1 U12179 ( .A1(n2676), .A2(n3117), .ZN(\mult_22/ab[63][49] ) );
  NOR2_X1 U12180 ( .A1(n2566), .A2(n3116), .ZN(\mult_22/ab[63][31] ) );
  NOR2_X1 U12181 ( .A1(n2684), .A2(n3117), .ZN(\mult_22/ab[63][51] ) );
  NOR2_X1 U12182 ( .A1(n2678), .A2(n3117), .ZN(\mult_22/ab[63][50] ) );
  NOR2_X1 U12183 ( .A1(n2595), .A2(n3116), .ZN(\mult_22/ab[63][36] ) );
  NOR2_X1 U12184 ( .A1(n2577), .A2(n3116), .ZN(\mult_22/ab[63][33] ) );
  NOR2_X1 U12185 ( .A1(n2583), .A2(n3116), .ZN(\mult_22/ab[63][34] ) );
  NOR2_X1 U12186 ( .A1(n2554), .A2(n3115), .ZN(\mult_22/ab[63][29] ) );
  NOR2_X1 U12187 ( .A1(n2718), .A2(n3118), .ZN(\mult_22/ab[63][57] ) );
  NOR2_X1 U12188 ( .A1(n2600), .A2(n2862), .ZN(n952) );
  NOR2_X1 U12189 ( .A1(n2727), .A2(n3118), .ZN(\mult_22/ab[63][59] ) );
  NOR2_X1 U12190 ( .A1(n2186), .A2(n2920), .ZN(\mult_22/ab[30][62] ) );
  NOR2_X1 U12191 ( .A1(n2751), .A2(n2914), .ZN(\mult_22/ab[29][63] ) );
  NOR2_X1 U12192 ( .A1(n2185), .A2(n2926), .ZN(\mult_22/ab[31][62] ) );
  NOR2_X1 U12193 ( .A1(n2751), .A2(n2920), .ZN(\mult_22/ab[30][63] ) );
  NOR2_X1 U12194 ( .A1(n2744), .A2(n2932), .ZN(\mult_22/ab[32][62] ) );
  NOR2_X1 U12195 ( .A1(n2751), .A2(n2926), .ZN(\mult_22/ab[31][63] ) );
  NOR2_X1 U12196 ( .A1(n2751), .A2(n2932), .ZN(\mult_22/ab[32][63] ) );
  NOR2_X1 U12197 ( .A1(n2745), .A2(n2938), .ZN(\mult_22/ab[33][62] ) );
  NOR2_X1 U12198 ( .A1(n2186), .A2(n2944), .ZN(\mult_22/ab[34][62] ) );
  NOR2_X1 U12199 ( .A1(n2751), .A2(n2938), .ZN(\mult_22/ab[33][63] ) );
  NOR2_X1 U12200 ( .A1(n2185), .A2(n2950), .ZN(\mult_22/ab[35][62] ) );
  NOR2_X1 U12201 ( .A1(n2751), .A2(n2944), .ZN(\mult_22/ab[34][63] ) );
  NOR2_X1 U12202 ( .A1(n2751), .A2(n2950), .ZN(\mult_22/ab[35][63] ) );
  NOR2_X1 U12203 ( .A1(n2745), .A2(n2956), .ZN(\mult_22/ab[36][62] ) );
  NOR2_X1 U12204 ( .A1(n2748), .A2(n3088), .ZN(\mult_22/ab[58][63] ) );
  NOR2_X1 U12205 ( .A1(n2745), .A2(n3094), .ZN(\mult_22/ab[59][62] ) );
  NOR2_X1 U12206 ( .A1(n2748), .A2(n3094), .ZN(\mult_22/ab[59][63] ) );
  NOR2_X1 U12207 ( .A1(n2746), .A2(n3100), .ZN(\mult_22/ab[60][62] ) );
  NOR2_X1 U12208 ( .A1(n2744), .A2(n2962), .ZN(\mult_22/ab[37][62] ) );
  NOR2_X1 U12209 ( .A1(n2750), .A2(n2956), .ZN(\mult_22/ab[36][63] ) );
  NOR2_X1 U12210 ( .A1(n2186), .A2(n2968), .ZN(\mult_22/ab[38][62] ) );
  NOR2_X1 U12211 ( .A1(n2750), .A2(n2962), .ZN(\mult_22/ab[37][63] ) );
  NOR2_X1 U12212 ( .A1(n2185), .A2(n2974), .ZN(\mult_22/ab[39][62] ) );
  NOR2_X1 U12213 ( .A1(n2750), .A2(n2968), .ZN(\mult_22/ab[38][63] ) );
  NOR2_X1 U12214 ( .A1(n2745), .A2(n2980), .ZN(\mult_22/ab[40][62] ) );
  NOR2_X1 U12215 ( .A1(n2750), .A2(n2974), .ZN(\mult_22/ab[39][63] ) );
  NOR2_X1 U12216 ( .A1(n2745), .A2(n3028), .ZN(\mult_22/ab[48][62] ) );
  NOR2_X1 U12217 ( .A1(n2749), .A2(n3022), .ZN(\mult_22/ab[47][63] ) );
  NOR2_X1 U12218 ( .A1(n2746), .A2(n2986), .ZN(\mult_22/ab[41][62] ) );
  NOR2_X1 U12219 ( .A1(n2750), .A2(n2980), .ZN(\mult_22/ab[40][63] ) );
  NOR2_X1 U12220 ( .A1(n2185), .A2(n3022), .ZN(\mult_22/ab[47][62] ) );
  NOR2_X1 U12221 ( .A1(n2749), .A2(n3016), .ZN(\mult_22/ab[46][63] ) );
  NOR2_X1 U12222 ( .A1(n2747), .A2(n2992), .ZN(\mult_22/ab[42][62] ) );
  NOR2_X1 U12223 ( .A1(n2750), .A2(n2986), .ZN(\mult_22/ab[41][63] ) );
  NOR2_X1 U12224 ( .A1(n2744), .A2(n3034), .ZN(\mult_22/ab[49][62] ) );
  NOR2_X1 U12225 ( .A1(n2749), .A2(n3028), .ZN(\mult_22/ab[48][63] ) );
  NOR2_X1 U12226 ( .A1(n2743), .A2(n2998), .ZN(\mult_22/ab[43][62] ) );
  NOR2_X1 U12227 ( .A1(n2750), .A2(n2992), .ZN(\mult_22/ab[42][63] ) );
  NOR2_X1 U12228 ( .A1(n2744), .A2(n3004), .ZN(\mult_22/ab[44][62] ) );
  NOR2_X1 U12229 ( .A1(n2750), .A2(n2998), .ZN(\mult_22/ab[43][63] ) );
  NOR2_X1 U12230 ( .A1(n2186), .A2(n3010), .ZN(\mult_22/ab[45][62] ) );
  NOR2_X1 U12231 ( .A1(n2750), .A2(n3004), .ZN(\mult_22/ab[44][63] ) );
  NOR2_X1 U12232 ( .A1(n2744), .A2(n3016), .ZN(\mult_22/ab[46][62] ) );
  NOR2_X1 U12233 ( .A1(n2750), .A2(n3010), .ZN(\mult_22/ab[45][63] ) );
  NOR2_X1 U12234 ( .A1(n2186), .A2(n3040), .ZN(\mult_22/ab[50][62] ) );
  NOR2_X1 U12235 ( .A1(n2749), .A2(n3034), .ZN(\mult_22/ab[49][63] ) );
  NOR2_X1 U12236 ( .A1(n2185), .A2(n3046), .ZN(\mult_22/ab[51][62] ) );
  NOR2_X1 U12237 ( .A1(n2749), .A2(n3040), .ZN(\mult_22/ab[50][63] ) );
  NOR2_X1 U12238 ( .A1(n2745), .A2(n3052), .ZN(\mult_22/ab[52][62] ) );
  NOR2_X1 U12239 ( .A1(n2749), .A2(n3046), .ZN(\mult_22/ab[51][63] ) );
  NOR2_X1 U12240 ( .A1(n2746), .A2(n3058), .ZN(\mult_22/ab[53][62] ) );
  NOR2_X1 U12241 ( .A1(n2749), .A2(n3052), .ZN(\mult_22/ab[52][63] ) );
  NOR2_X1 U12242 ( .A1(n2747), .A2(n3064), .ZN(\mult_22/ab[54][62] ) );
  NOR2_X1 U12243 ( .A1(n2749), .A2(n3058), .ZN(\mult_22/ab[53][63] ) );
  NOR2_X1 U12244 ( .A1(n2743), .A2(n3070), .ZN(\mult_22/ab[55][62] ) );
  NOR2_X1 U12245 ( .A1(n2749), .A2(n3064), .ZN(\mult_22/ab[54][63] ) );
  NOR2_X1 U12246 ( .A1(n2186), .A2(n3076), .ZN(\mult_22/ab[56][62] ) );
  NOR2_X1 U12247 ( .A1(n2749), .A2(n3070), .ZN(\mult_22/ab[55][63] ) );
  NOR2_X1 U12248 ( .A1(n2185), .A2(n3082), .ZN(\mult_22/ab[57][62] ) );
  NOR2_X1 U12249 ( .A1(n2749), .A2(n3076), .ZN(\mult_22/ab[56][63] ) );
  NOR2_X1 U12250 ( .A1(n2748), .A2(n3082), .ZN(\mult_22/ab[57][63] ) );
  NOR2_X1 U12251 ( .A1(n2744), .A2(n3088), .ZN(\mult_22/ab[58][62] ) );
  NOR2_X1 U12252 ( .A1(n2560), .A2(n3109), .ZN(\mult_22/ab[62][30] ) );
  NOR2_X1 U12253 ( .A1(n2607), .A2(n3110), .ZN(\mult_22/ab[62][38] ) );
  NOR2_X1 U12254 ( .A1(n2612), .A2(n3110), .ZN(\mult_22/ab[62][39] ) );
  NOR2_X1 U12255 ( .A1(n2566), .A2(n3104), .ZN(\mult_22/ab[61][31] ) );
  NOR2_X1 U12256 ( .A1(n2566), .A2(n3110), .ZN(\mult_22/ab[62][31] ) );
  NOR2_X1 U12257 ( .A1(n2601), .A2(n3110), .ZN(\mult_22/ab[62][37] ) );
  NOR2_X1 U12258 ( .A1(n2618), .A2(n3110), .ZN(\mult_22/ab[62][40] ) );
  NOR2_X1 U12259 ( .A1(n2595), .A2(n3110), .ZN(\mult_22/ab[62][36] ) );
  NOR2_X1 U12260 ( .A1(n2666), .A2(n3111), .ZN(\mult_22/ab[62][48] ) );
  NOR2_X1 U12261 ( .A1(n2660), .A2(n3111), .ZN(\mult_22/ab[62][47] ) );
  NOR2_X1 U12262 ( .A1(n2628), .A2(n3110), .ZN(\mult_22/ab[62][41] ) );
  NOR2_X1 U12263 ( .A1(n2652), .A2(n3111), .ZN(\mult_22/ab[62][45] ) );
  NOR2_X1 U12264 ( .A1(n2676), .A2(n3111), .ZN(\mult_22/ab[62][49] ) );
  NOR2_X1 U12265 ( .A1(n2642), .A2(n3111), .ZN(\mult_22/ab[62][44] ) );
  NOR2_X1 U12266 ( .A1(n2576), .A2(n3098), .ZN(\mult_22/ab[60][32] ) );
  NOR2_X1 U12267 ( .A1(n2601), .A2(n3104), .ZN(\mult_22/ab[61][37] ) );
  NOR2_X1 U12268 ( .A1(n2612), .A2(n3104), .ZN(\mult_22/ab[61][39] ) );
  NOR2_X1 U12269 ( .A1(n2607), .A2(n3104), .ZN(\mult_22/ab[61][38] ) );
  NOR2_X1 U12270 ( .A1(n2576), .A2(n3104), .ZN(\mult_22/ab[61][32] ) );
  NOR2_X1 U12271 ( .A1(n2576), .A2(n3110), .ZN(\mult_22/ab[62][32] ) );
  NOR2_X1 U12272 ( .A1(n2640), .A2(n3111), .ZN(\mult_22/ab[62][43] ) );
  NOR2_X1 U12273 ( .A1(n2630), .A2(n3111), .ZN(\mult_22/ab[62][42] ) );
  NOR2_X1 U12274 ( .A1(n2618), .A2(n3104), .ZN(\mult_22/ab[61][40] ) );
  NOR2_X1 U12275 ( .A1(n2654), .A2(n3111), .ZN(\mult_22/ab[62][46] ) );
  NOR2_X1 U12276 ( .A1(n2601), .A2(n3098), .ZN(\mult_22/ab[60][37] ) );
  NOR2_X1 U12277 ( .A1(n2607), .A2(n3098), .ZN(\mult_22/ab[60][38] ) );
  NOR2_X1 U12278 ( .A1(n2577), .A2(n3092), .ZN(\mult_22/ab[59][33] ) );
  NOR2_X1 U12279 ( .A1(n2676), .A2(n3105), .ZN(\mult_22/ab[61][49] ) );
  NOR2_X1 U12280 ( .A1(n2612), .A2(n3098), .ZN(\mult_22/ab[60][39] ) );
  NOR2_X1 U12281 ( .A1(n2630), .A2(n3105), .ZN(\mult_22/ab[61][42] ) );
  NOR2_X1 U12282 ( .A1(n2666), .A2(n3105), .ZN(\mult_22/ab[61][48] ) );
  NOR2_X1 U12283 ( .A1(n2618), .A2(n3098), .ZN(\mult_22/ab[60][40] ) );
  NOR2_X1 U12284 ( .A1(n2601), .A2(n3092), .ZN(\mult_22/ab[59][37] ) );
  NOR2_X1 U12285 ( .A1(n2607), .A2(n3092), .ZN(\mult_22/ab[59][38] ) );
  NOR2_X1 U12286 ( .A1(n2678), .A2(n3111), .ZN(\mult_22/ab[62][50] ) );
  NOR2_X1 U12287 ( .A1(n2628), .A2(n3098), .ZN(\mult_22/ab[60][41] ) );
  NOR2_X1 U12288 ( .A1(n2612), .A2(n3092), .ZN(\mult_22/ab[59][39] ) );
  NOR2_X1 U12289 ( .A1(n2652), .A2(n3105), .ZN(\mult_22/ab[61][45] ) );
  NOR2_X1 U12290 ( .A1(n2678), .A2(n3105), .ZN(\mult_22/ab[61][50] ) );
  NOR2_X1 U12291 ( .A1(n2640), .A2(n3105), .ZN(\mult_22/ab[61][43] ) );
  NOR2_X1 U12292 ( .A1(n2642), .A2(n3105), .ZN(\mult_22/ab[61][44] ) );
  NOR2_X1 U12293 ( .A1(n2601), .A2(n3086), .ZN(\mult_22/ab[58][37] ) );
  NOR2_X1 U12294 ( .A1(n2654), .A2(n3105), .ZN(\mult_22/ab[61][46] ) );
  NOR2_X1 U12295 ( .A1(n2630), .A2(n3099), .ZN(\mult_22/ab[60][42] ) );
  NOR2_X1 U12296 ( .A1(n2618), .A2(n3092), .ZN(\mult_22/ab[59][40] ) );
  NOR2_X1 U12297 ( .A1(n2612), .A2(n3086), .ZN(\mult_22/ab[58][39] ) );
  NOR2_X1 U12298 ( .A1(n2660), .A2(n3105), .ZN(\mult_22/ab[61][47] ) );
  NOR2_X1 U12299 ( .A1(n2628), .A2(n3092), .ZN(\mult_22/ab[59][41] ) );
  NOR2_X1 U12300 ( .A1(n2602), .A2(n3080), .ZN(\mult_22/ab[57][37] ) );
  NOR2_X1 U12301 ( .A1(n2678), .A2(n3099), .ZN(\mult_22/ab[60][50] ) );
  NOR2_X1 U12302 ( .A1(n2602), .A2(n3068), .ZN(\mult_22/ab[55][37] ) );
  NOR2_X1 U12303 ( .A1(n2602), .A2(n3074), .ZN(\mult_22/ab[56][37] ) );
  NOR2_X1 U12304 ( .A1(n2640), .A2(n3099), .ZN(\mult_22/ab[60][43] ) );
  NOR2_X1 U12305 ( .A1(n2628), .A2(n3068), .ZN(\mult_22/ab[55][41] ) );
  NOR2_X1 U12306 ( .A1(n2674), .A2(n2997), .ZN(\mult_22/ab[43][49] ) );
  NOR2_X1 U12307 ( .A1(n2662), .A2(n3015), .ZN(\mult_22/ab[46][47] ) );
  NOR2_X1 U12308 ( .A1(n2651), .A2(n3033), .ZN(\mult_22/ab[49][45] ) );
  NOR2_X1 U12309 ( .A1(n2639), .A2(n3051), .ZN(\mult_22/ab[52][43] ) );
  NOR2_X1 U12310 ( .A1(n2628), .A2(n3074), .ZN(\mult_22/ab[56][41] ) );
  NOR2_X1 U12311 ( .A1(n2662), .A2(n3021), .ZN(\mult_22/ab[47][47] ) );
  NOR2_X1 U12312 ( .A1(n2651), .A2(n3039), .ZN(\mult_22/ab[50][45] ) );
  NOR2_X1 U12313 ( .A1(n2639), .A2(n3057), .ZN(\mult_22/ab[53][43] ) );
  NOR2_X1 U12314 ( .A1(n2686), .A2(n2985), .ZN(\mult_22/ab[41][51] ) );
  NOR2_X1 U12315 ( .A1(n2675), .A2(n3003), .ZN(\mult_22/ab[44][49] ) );
  NOR2_X1 U12316 ( .A1(n2675), .A2(n3009), .ZN(\mult_22/ab[45][49] ) );
  NOR2_X1 U12317 ( .A1(n2661), .A2(n3027), .ZN(\mult_22/ab[48][47] ) );
  NOR2_X1 U12318 ( .A1(n2651), .A2(n3045), .ZN(\mult_22/ab[51][45] ) );
  NOR2_X1 U12319 ( .A1(n2639), .A2(n3063), .ZN(\mult_22/ab[54][43] ) );
  NOR2_X1 U12320 ( .A1(n2367), .A2(n2974), .ZN(\mult_22/ab[39][53] ) );
  NOR2_X1 U12321 ( .A1(n2686), .A2(n2991), .ZN(\mult_22/ab[42][51] ) );
  NOR2_X1 U12322 ( .A1(n2675), .A2(n3015), .ZN(\mult_22/ab[46][49] ) );
  NOR2_X1 U12323 ( .A1(n2661), .A2(n3033), .ZN(\mult_22/ab[49][47] ) );
  NOR2_X1 U12324 ( .A1(n2651), .A2(n3051), .ZN(\mult_22/ab[52][45] ) );
  NOR2_X1 U12325 ( .A1(n2708), .A2(n2962), .ZN(\mult_22/ab[37][55] ) );
  NOR2_X1 U12326 ( .A1(n2699), .A2(n2980), .ZN(\mult_22/ab[40][53] ) );
  NOR2_X1 U12327 ( .A1(n2686), .A2(n2997), .ZN(\mult_22/ab[43][51] ) );
  NOR2_X1 U12328 ( .A1(n2675), .A2(n3021), .ZN(\mult_22/ab[47][49] ) );
  NOR2_X1 U12329 ( .A1(n2661), .A2(n3039), .ZN(\mult_22/ab[50][47] ) );
  NOR2_X1 U12330 ( .A1(n2716), .A2(n2950), .ZN(\mult_22/ab[35][57] ) );
  NOR2_X1 U12331 ( .A1(n2708), .A2(n2968), .ZN(\mult_22/ab[38][55] ) );
  NOR2_X1 U12332 ( .A1(n2700), .A2(n2986), .ZN(\mult_22/ab[41][53] ) );
  NOR2_X1 U12333 ( .A1(n2686), .A2(n3003), .ZN(\mult_22/ab[44][51] ) );
  NOR2_X1 U12334 ( .A1(n2686), .A2(n3009), .ZN(\mult_22/ab[45][51] ) );
  NOR2_X1 U12335 ( .A1(n2675), .A2(n3027), .ZN(\mult_22/ab[48][49] ) );
  NOR2_X1 U12336 ( .A1(n2716), .A2(n2956), .ZN(\mult_22/ab[36][57] ) );
  NOR2_X1 U12337 ( .A1(n2708), .A2(n2974), .ZN(\mult_22/ab[39][55] ) );
  NOR2_X1 U12338 ( .A1(n2696), .A2(n2992), .ZN(\mult_22/ab[42][53] ) );
  NOR2_X1 U12339 ( .A1(n2727), .A2(n2938), .ZN(\mult_22/ab[33][59] ) );
  NOR2_X1 U12340 ( .A1(n2686), .A2(n3015), .ZN(\mult_22/ab[46][51] ) );
  NOR2_X1 U12341 ( .A1(n2728), .A2(n2944), .ZN(\mult_22/ab[34][59] ) );
  NOR2_X1 U12342 ( .A1(n2716), .A2(n2962), .ZN(\mult_22/ab[37][57] ) );
  NOR2_X1 U12343 ( .A1(n2708), .A2(n2980), .ZN(\mult_22/ab[40][55] ) );
  NOR2_X1 U12344 ( .A1(n2697), .A2(n2998), .ZN(\mult_22/ab[43][53] ) );
  NOR2_X1 U12345 ( .A1(n2708), .A2(n2986), .ZN(\mult_22/ab[41][55] ) );
  NOR2_X1 U12346 ( .A1(n2695), .A2(n3004), .ZN(\mult_22/ab[44][53] ) );
  NOR2_X1 U12347 ( .A1(n2729), .A2(n2950), .ZN(\mult_22/ab[35][59] ) );
  NOR2_X1 U12348 ( .A1(n2716), .A2(n2968), .ZN(\mult_22/ab[38][57] ) );
  NOR2_X1 U12349 ( .A1(n2708), .A2(n2992), .ZN(\mult_22/ab[42][55] ) );
  NOR2_X1 U12350 ( .A1(n2730), .A2(n2956), .ZN(\mult_22/ab[36][59] ) );
  NOR2_X1 U12351 ( .A1(n2716), .A2(n2974), .ZN(\mult_22/ab[39][57] ) );
  NOR2_X1 U12352 ( .A1(n2725), .A2(n2962), .ZN(\mult_22/ab[37][59] ) );
  NOR2_X1 U12353 ( .A1(n2716), .A2(n2980), .ZN(\mult_22/ab[40][57] ) );
  NOR2_X1 U12354 ( .A1(n2726), .A2(n2968), .ZN(\mult_22/ab[38][59] ) );
  NOR2_X1 U12355 ( .A1(n2656), .A2(n3015), .ZN(\mult_22/ab[46][46] ) );
  NOR2_X1 U12356 ( .A1(n2643), .A2(n3027), .ZN(\mult_22/ab[48][44] ) );
  NOR2_X1 U12357 ( .A1(n2631), .A2(n3039), .ZN(\mult_22/ab[50][42] ) );
  NOR2_X1 U12358 ( .A1(n2619), .A2(n3050), .ZN(\mult_22/ab[52][40] ) );
  NOR2_X1 U12359 ( .A1(n2643), .A2(n3033), .ZN(\mult_22/ab[49][44] ) );
  NOR2_X1 U12360 ( .A1(n2631), .A2(n3045), .ZN(\mult_22/ab[51][42] ) );
  NOR2_X1 U12361 ( .A1(n2631), .A2(n3051), .ZN(\mult_22/ab[52][42] ) );
  NOR2_X1 U12362 ( .A1(n2619), .A2(n3056), .ZN(\mult_22/ab[53][40] ) );
  NOR2_X1 U12363 ( .A1(n2619), .A2(n3062), .ZN(\mult_22/ab[54][40] ) );
  NOR2_X1 U12364 ( .A1(n2619), .A2(n3068), .ZN(\mult_22/ab[55][40] ) );
  NOR2_X1 U12365 ( .A1(n2668), .A2(n3003), .ZN(\mult_22/ab[44][48] ) );
  NOR2_X1 U12366 ( .A1(n2655), .A2(n3021), .ZN(\mult_22/ab[47][46] ) );
  NOR2_X1 U12367 ( .A1(n2643), .A2(n3039), .ZN(\mult_22/ab[50][44] ) );
  NOR2_X1 U12368 ( .A1(n2631), .A2(n3057), .ZN(\mult_22/ab[53][42] ) );
  NOR2_X1 U12369 ( .A1(n2619), .A2(n3074), .ZN(\mult_22/ab[56][40] ) );
  NOR2_X1 U12370 ( .A1(n2619), .A2(n3080), .ZN(\mult_22/ab[57][40] ) );
  NOR2_X1 U12371 ( .A1(n2655), .A2(n3027), .ZN(\mult_22/ab[48][46] ) );
  NOR2_X1 U12372 ( .A1(n2643), .A2(n3045), .ZN(\mult_22/ab[51][44] ) );
  NOR2_X1 U12373 ( .A1(n2631), .A2(n3063), .ZN(\mult_22/ab[54][42] ) );
  NOR2_X1 U12374 ( .A1(n2680), .A2(n2991), .ZN(\mult_22/ab[42][50] ) );
  NOR2_X1 U12375 ( .A1(n2668), .A2(n3009), .ZN(\mult_22/ab[45][48] ) );
  NOR2_X1 U12376 ( .A1(n2668), .A2(n3015), .ZN(\mult_22/ab[46][48] ) );
  NOR2_X1 U12377 ( .A1(n2655), .A2(n3033), .ZN(\mult_22/ab[49][46] ) );
  NOR2_X1 U12378 ( .A1(n2643), .A2(n3051), .ZN(\mult_22/ab[52][44] ) );
  NOR2_X1 U12379 ( .A1(n2631), .A2(n3069), .ZN(\mult_22/ab[55][42] ) );
  NOR2_X1 U12380 ( .A1(n2692), .A2(n2979), .ZN(\mult_22/ab[40][52] ) );
  NOR2_X1 U12381 ( .A1(n2680), .A2(n2997), .ZN(\mult_22/ab[43][50] ) );
  NOR2_X1 U12382 ( .A1(n2667), .A2(n3021), .ZN(\mult_22/ab[47][48] ) );
  NOR2_X1 U12383 ( .A1(n2655), .A2(n3039), .ZN(\mult_22/ab[50][46] ) );
  NOR2_X1 U12384 ( .A1(n2643), .A2(n3057), .ZN(\mult_22/ab[53][44] ) );
  NOR2_X1 U12385 ( .A1(n2702), .A2(n2968), .ZN(\mult_22/ab[38][54] ) );
  NOR2_X1 U12386 ( .A1(n2692), .A2(n2985), .ZN(\mult_22/ab[41][52] ) );
  NOR2_X1 U12387 ( .A1(n2680), .A2(n3003), .ZN(\mult_22/ab[44][50] ) );
  NOR2_X1 U12388 ( .A1(n2692), .A2(n2991), .ZN(\mult_22/ab[42][52] ) );
  NOR2_X1 U12389 ( .A1(n2680), .A2(n3009), .ZN(\mult_22/ab[45][50] ) );
  NOR2_X1 U12390 ( .A1(n2667), .A2(n3027), .ZN(\mult_22/ab[48][48] ) );
  NOR2_X1 U12391 ( .A1(n2655), .A2(n3045), .ZN(\mult_22/ab[51][46] ) );
  NOR2_X1 U12392 ( .A1(n2712), .A2(n2956), .ZN(\mult_22/ab[36][56] ) );
  NOR2_X1 U12393 ( .A1(n2702), .A2(n2974), .ZN(\mult_22/ab[39][54] ) );
  NOR2_X1 U12394 ( .A1(n2679), .A2(n3015), .ZN(\mult_22/ab[46][50] ) );
  NOR2_X1 U12395 ( .A1(n2667), .A2(n3033), .ZN(\mult_22/ab[49][48] ) );
  NOR2_X1 U12396 ( .A1(n2721), .A2(n2944), .ZN(\mult_22/ab[34][58] ) );
  NOR2_X1 U12397 ( .A1(n2712), .A2(n2962), .ZN(\mult_22/ab[37][56] ) );
  NOR2_X1 U12398 ( .A1(n2702), .A2(n2980), .ZN(\mult_22/ab[40][54] ) );
  NOR2_X1 U12399 ( .A1(n2692), .A2(n2997), .ZN(\mult_22/ab[43][52] ) );
  NOR2_X1 U12400 ( .A1(n2693), .A2(n3003), .ZN(\mult_22/ab[44][52] ) );
  NOR2_X1 U12401 ( .A1(n2679), .A2(n3021), .ZN(\mult_22/ab[47][50] ) );
  NOR2_X1 U12402 ( .A1(n2702), .A2(n2986), .ZN(\mult_22/ab[41][54] ) );
  NOR2_X1 U12403 ( .A1(n2721), .A2(n2950), .ZN(\mult_22/ab[35][58] ) );
  NOR2_X1 U12404 ( .A1(n2712), .A2(n2968), .ZN(\mult_22/ab[38][56] ) );
  NOR2_X1 U12405 ( .A1(n2693), .A2(n3009), .ZN(\mult_22/ab[45][52] ) );
  NOR2_X1 U12406 ( .A1(n2721), .A2(n2956), .ZN(\mult_22/ab[36][58] ) );
  NOR2_X1 U12407 ( .A1(n2712), .A2(n2974), .ZN(\mult_22/ab[39][56] ) );
  NOR2_X1 U12408 ( .A1(n2702), .A2(n2992), .ZN(\mult_22/ab[42][54] ) );
  NOR2_X1 U12409 ( .A1(n2712), .A2(n2980), .ZN(\mult_22/ab[40][56] ) );
  NOR2_X1 U12410 ( .A1(n2702), .A2(n2998), .ZN(\mult_22/ab[43][54] ) );
  NOR2_X1 U12411 ( .A1(n2721), .A2(n2962), .ZN(\mult_22/ab[37][58] ) );
  NOR2_X1 U12412 ( .A1(n2721), .A2(n2968), .ZN(\mult_22/ab[38][58] ) );
  NOR2_X1 U12413 ( .A1(n2712), .A2(n2986), .ZN(\mult_22/ab[41][56] ) );
  NOR2_X1 U12414 ( .A1(n2721), .A2(n2974), .ZN(\mult_22/ab[39][58] ) );
  NOR2_X1 U12415 ( .A1(n2732), .A2(n2932), .ZN(\mult_22/ab[32][60] ) );
  NOR2_X1 U12416 ( .A1(n2733), .A2(n2938), .ZN(\mult_22/ab[33][60] ) );
  NOR2_X1 U12417 ( .A1(n2733), .A2(n2944), .ZN(\mult_22/ab[34][60] ) );
  NOR2_X1 U12418 ( .A1(n2733), .A2(n2950), .ZN(\mult_22/ab[35][60] ) );
  NOR2_X1 U12419 ( .A1(n2733), .A2(n2956), .ZN(\mult_22/ab[36][60] ) );
  NOR2_X1 U12420 ( .A1(n2733), .A2(n2962), .ZN(\mult_22/ab[37][60] ) );
  NOR2_X1 U12421 ( .A1(n2739), .A2(n2926), .ZN(\mult_22/ab[31][61] ) );
  NOR2_X1 U12422 ( .A1(n2738), .A2(n2932), .ZN(\mult_22/ab[32][61] ) );
  NOR2_X1 U12423 ( .A1(n2739), .A2(n2938), .ZN(\mult_22/ab[33][61] ) );
  NOR2_X1 U12424 ( .A1(n2737), .A2(n2944), .ZN(\mult_22/ab[34][61] ) );
  NOR2_X1 U12425 ( .A1(n2740), .A2(n2950), .ZN(\mult_22/ab[35][61] ) );
  NOR2_X1 U12426 ( .A1(n2741), .A2(n2956), .ZN(\mult_22/ab[36][61] ) );
  NOR2_X1 U12427 ( .A1(n2618), .A2(n3086), .ZN(\mult_22/ab[58][40] ) );
  NOR2_X1 U12428 ( .A1(n2676), .A2(n3099), .ZN(\mult_22/ab[60][49] ) );
  NOR2_X1 U12429 ( .A1(n2630), .A2(n3093), .ZN(\mult_22/ab[59][42] ) );
  NOR2_X1 U12430 ( .A1(n2628), .A2(n3080), .ZN(\mult_22/ab[57][41] ) );
  NOR2_X1 U12431 ( .A1(n2640), .A2(n3069), .ZN(\mult_22/ab[55][43] ) );
  NOR2_X1 U12432 ( .A1(n2651), .A2(n3057), .ZN(\mult_22/ab[53][45] ) );
  NOR2_X1 U12433 ( .A1(n2661), .A2(n3045), .ZN(\mult_22/ab[51][47] ) );
  NOR2_X1 U12434 ( .A1(n2675), .A2(n3033), .ZN(\mult_22/ab[49][49] ) );
  NOR2_X1 U12435 ( .A1(n2686), .A2(n3021), .ZN(\mult_22/ab[47][51] ) );
  NOR2_X1 U12436 ( .A1(n2700), .A2(n3010), .ZN(\mult_22/ab[45][53] ) );
  NOR2_X1 U12437 ( .A1(n2708), .A2(n2998), .ZN(\mult_22/ab[43][55] ) );
  NOR2_X1 U12438 ( .A1(n2716), .A2(n2986), .ZN(\mult_22/ab[41][57] ) );
  NOR2_X1 U12439 ( .A1(n2727), .A2(n2974), .ZN(\mult_22/ab[39][59] ) );
  NOR2_X1 U12440 ( .A1(n2631), .A2(n3075), .ZN(\mult_22/ab[56][42] ) );
  NOR2_X1 U12441 ( .A1(n2643), .A2(n3063), .ZN(\mult_22/ab[54][44] ) );
  NOR2_X1 U12442 ( .A1(n2655), .A2(n3051), .ZN(\mult_22/ab[52][46] ) );
  NOR2_X1 U12443 ( .A1(n2667), .A2(n3039), .ZN(\mult_22/ab[50][48] ) );
  NOR2_X1 U12444 ( .A1(n2679), .A2(n3027), .ZN(\mult_22/ab[48][50] ) );
  NOR2_X1 U12445 ( .A1(n2693), .A2(n3015), .ZN(\mult_22/ab[46][52] ) );
  NOR2_X1 U12446 ( .A1(n2702), .A2(n3004), .ZN(\mult_22/ab[44][54] ) );
  NOR2_X1 U12447 ( .A1(n2712), .A2(n2992), .ZN(\mult_22/ab[42][56] ) );
  NOR2_X1 U12448 ( .A1(n2721), .A2(n2980), .ZN(\mult_22/ab[40][58] ) );
  NOR2_X1 U12449 ( .A1(n2733), .A2(n2968), .ZN(\mult_22/ab[38][60] ) );
  NOR2_X1 U12450 ( .A1(n2738), .A2(n2962), .ZN(\mult_22/ab[37][61] ) );
  NOR2_X1 U12451 ( .A1(n2628), .A2(n3086), .ZN(\mult_22/ab[58][41] ) );
  NOR2_X1 U12452 ( .A1(n2640), .A2(n3075), .ZN(\mult_22/ab[56][43] ) );
  NOR2_X1 U12453 ( .A1(n2651), .A2(n3063), .ZN(\mult_22/ab[54][45] ) );
  NOR2_X1 U12454 ( .A1(n2661), .A2(n3051), .ZN(\mult_22/ab[52][47] ) );
  NOR2_X1 U12455 ( .A1(n2675), .A2(n3039), .ZN(\mult_22/ab[50][49] ) );
  NOR2_X1 U12456 ( .A1(n2685), .A2(n3027), .ZN(\mult_22/ab[48][51] ) );
  NOR2_X1 U12457 ( .A1(n2367), .A2(n3016), .ZN(\mult_22/ab[46][53] ) );
  NOR2_X1 U12458 ( .A1(n2708), .A2(n3004), .ZN(\mult_22/ab[44][55] ) );
  NOR2_X1 U12459 ( .A1(n2716), .A2(n2992), .ZN(\mult_22/ab[42][57] ) );
  NOR2_X1 U12460 ( .A1(n2728), .A2(n2980), .ZN(\mult_22/ab[40][59] ) );
  NOR2_X1 U12461 ( .A1(n2631), .A2(n3081), .ZN(\mult_22/ab[57][42] ) );
  NOR2_X1 U12462 ( .A1(n2643), .A2(n3069), .ZN(\mult_22/ab[55][44] ) );
  NOR2_X1 U12463 ( .A1(n2655), .A2(n3057), .ZN(\mult_22/ab[53][46] ) );
  NOR2_X1 U12464 ( .A1(n2667), .A2(n3045), .ZN(\mult_22/ab[51][48] ) );
  NOR2_X1 U12465 ( .A1(n2679), .A2(n3033), .ZN(\mult_22/ab[49][50] ) );
  NOR2_X1 U12466 ( .A1(n2693), .A2(n3021), .ZN(\mult_22/ab[47][52] ) );
  NOR2_X1 U12467 ( .A1(n2702), .A2(n3010), .ZN(\mult_22/ab[45][54] ) );
  NOR2_X1 U12468 ( .A1(n2712), .A2(n2998), .ZN(\mult_22/ab[43][56] ) );
  NOR2_X1 U12469 ( .A1(n2721), .A2(n2986), .ZN(\mult_22/ab[41][58] ) );
  NOR2_X1 U12470 ( .A1(n2733), .A2(n2974), .ZN(\mult_22/ab[39][60] ) );
  NOR2_X1 U12471 ( .A1(n2737), .A2(n2968), .ZN(\mult_22/ab[38][61] ) );
  NOR2_X1 U12472 ( .A1(n2640), .A2(n3081), .ZN(\mult_22/ab[57][43] ) );
  NOR2_X1 U12473 ( .A1(n2652), .A2(n3069), .ZN(\mult_22/ab[55][45] ) );
  NOR2_X1 U12474 ( .A1(n2661), .A2(n3057), .ZN(\mult_22/ab[53][47] ) );
  NOR2_X1 U12475 ( .A1(n2675), .A2(n3045), .ZN(\mult_22/ab[51][49] ) );
  NOR2_X1 U12476 ( .A1(n2685), .A2(n3033), .ZN(\mult_22/ab[49][51] ) );
  NOR2_X1 U12477 ( .A1(n2699), .A2(n3022), .ZN(\mult_22/ab[47][53] ) );
  NOR2_X1 U12478 ( .A1(n2631), .A2(n3087), .ZN(\mult_22/ab[58][42] ) );
  NOR2_X1 U12479 ( .A1(n2708), .A2(n3010), .ZN(\mult_22/ab[45][55] ) );
  NOR2_X1 U12480 ( .A1(n2716), .A2(n2998), .ZN(\mult_22/ab[43][57] ) );
  NOR2_X1 U12481 ( .A1(n2729), .A2(n2986), .ZN(\mult_22/ab[41][59] ) );
  NOR2_X1 U12482 ( .A1(n2643), .A2(n3075), .ZN(\mult_22/ab[56][44] ) );
  NOR2_X1 U12483 ( .A1(n2655), .A2(n3063), .ZN(\mult_22/ab[54][46] ) );
  NOR2_X1 U12484 ( .A1(n2667), .A2(n3051), .ZN(\mult_22/ab[52][48] ) );
  NOR2_X1 U12485 ( .A1(n2679), .A2(n3039), .ZN(\mult_22/ab[50][50] ) );
  NOR2_X1 U12486 ( .A1(n2693), .A2(n3027), .ZN(\mult_22/ab[48][52] ) );
  NOR2_X1 U12487 ( .A1(n2702), .A2(n3016), .ZN(\mult_22/ab[46][54] ) );
  NOR2_X1 U12488 ( .A1(n2712), .A2(n3004), .ZN(\mult_22/ab[44][56] ) );
  NOR2_X1 U12489 ( .A1(n2721), .A2(n2992), .ZN(\mult_22/ab[42][58] ) );
  NOR2_X1 U12490 ( .A1(n2733), .A2(n2980), .ZN(\mult_22/ab[40][60] ) );
  NOR2_X1 U12491 ( .A1(n2739), .A2(n2974), .ZN(\mult_22/ab[39][61] ) );
  NOR2_X1 U12492 ( .A1(n2640), .A2(n3093), .ZN(\mult_22/ab[59][43] ) );
  NOR2_X1 U12493 ( .A1(n2642), .A2(n3099), .ZN(\mult_22/ab[60][44] ) );
  NOR2_X1 U12494 ( .A1(n2684), .A2(n3099), .ZN(\mult_22/ab[60][51] ) );
  NOR2_X1 U12495 ( .A1(n2640), .A2(n3087), .ZN(\mult_22/ab[58][43] ) );
  NOR2_X1 U12496 ( .A1(n2652), .A2(n3075), .ZN(\mult_22/ab[56][45] ) );
  NOR2_X1 U12497 ( .A1(n2661), .A2(n3063), .ZN(\mult_22/ab[54][47] ) );
  NOR2_X1 U12498 ( .A1(n2675), .A2(n3051), .ZN(\mult_22/ab[52][49] ) );
  NOR2_X1 U12499 ( .A1(n2685), .A2(n3039), .ZN(\mult_22/ab[50][51] ) );
  NOR2_X1 U12500 ( .A1(n2696), .A2(n3028), .ZN(\mult_22/ab[48][53] ) );
  NOR2_X1 U12501 ( .A1(n2708), .A2(n3016), .ZN(\mult_22/ab[46][55] ) );
  NOR2_X1 U12502 ( .A1(n2716), .A2(n3004), .ZN(\mult_22/ab[44][57] ) );
  NOR2_X1 U12503 ( .A1(n2730), .A2(n2992), .ZN(\mult_22/ab[42][59] ) );
  NOR2_X1 U12504 ( .A1(n2643), .A2(n3081), .ZN(\mult_22/ab[57][44] ) );
  NOR2_X1 U12505 ( .A1(n2655), .A2(n3069), .ZN(\mult_22/ab[55][46] ) );
  NOR2_X1 U12506 ( .A1(n2667), .A2(n3057), .ZN(\mult_22/ab[53][48] ) );
  NOR2_X1 U12507 ( .A1(n2679), .A2(n3045), .ZN(\mult_22/ab[51][50] ) );
  NOR2_X1 U12508 ( .A1(n2693), .A2(n3033), .ZN(\mult_22/ab[49][52] ) );
  NOR2_X1 U12509 ( .A1(n2701), .A2(n3022), .ZN(\mult_22/ab[47][54] ) );
  NOR2_X1 U12510 ( .A1(n2712), .A2(n3010), .ZN(\mult_22/ab[45][56] ) );
  NOR2_X1 U12511 ( .A1(n2721), .A2(n2998), .ZN(\mult_22/ab[43][58] ) );
  NOR2_X1 U12512 ( .A1(n2733), .A2(n2986), .ZN(\mult_22/ab[41][60] ) );
  NOR2_X1 U12513 ( .A1(n2740), .A2(n2980), .ZN(\mult_22/ab[40][61] ) );
  NOR2_X1 U12514 ( .A1(n2684), .A2(n3105), .ZN(\mult_22/ab[61][51] ) );
  NOR2_X1 U12515 ( .A1(n2652), .A2(n3099), .ZN(\mult_22/ab[60][45] ) );
  NOR2_X1 U12516 ( .A1(n2652), .A2(n3081), .ZN(\mult_22/ab[57][45] ) );
  NOR2_X1 U12517 ( .A1(n2661), .A2(n3069), .ZN(\mult_22/ab[55][47] ) );
  NOR2_X1 U12518 ( .A1(n2675), .A2(n3057), .ZN(\mult_22/ab[53][49] ) );
  NOR2_X1 U12519 ( .A1(n2685), .A2(n3045), .ZN(\mult_22/ab[51][51] ) );
  NOR2_X1 U12520 ( .A1(n2697), .A2(n3034), .ZN(\mult_22/ab[49][53] ) );
  NOR2_X1 U12521 ( .A1(n2707), .A2(n3022), .ZN(\mult_22/ab[47][55] ) );
  NOR2_X1 U12522 ( .A1(n2716), .A2(n3010), .ZN(\mult_22/ab[45][57] ) );
  NOR2_X1 U12523 ( .A1(n2725), .A2(n2998), .ZN(\mult_22/ab[43][59] ) );
  NOR2_X1 U12524 ( .A1(n2643), .A2(n3087), .ZN(\mult_22/ab[58][44] ) );
  NOR2_X1 U12525 ( .A1(n2655), .A2(n3075), .ZN(\mult_22/ab[56][46] ) );
  NOR2_X1 U12526 ( .A1(n2667), .A2(n3063), .ZN(\mult_22/ab[54][48] ) );
  NOR2_X1 U12527 ( .A1(n2679), .A2(n3051), .ZN(\mult_22/ab[52][50] ) );
  NOR2_X1 U12528 ( .A1(n2693), .A2(n3039), .ZN(\mult_22/ab[50][52] ) );
  NOR2_X1 U12529 ( .A1(n2701), .A2(n3028), .ZN(\mult_22/ab[48][54] ) );
  NOR2_X1 U12530 ( .A1(n2712), .A2(n3016), .ZN(\mult_22/ab[46][56] ) );
  NOR2_X1 U12531 ( .A1(n2722), .A2(n3004), .ZN(\mult_22/ab[44][58] ) );
  NOR2_X1 U12532 ( .A1(n2738), .A2(n2986), .ZN(\mult_22/ab[41][61] ) );
  NOR2_X1 U12533 ( .A1(n2733), .A2(n2992), .ZN(\mult_22/ab[42][60] ) );
  NOR2_X1 U12534 ( .A1(n2654), .A2(n3099), .ZN(\mult_22/ab[60][46] ) );
  NOR2_X1 U12535 ( .A1(n2652), .A2(n3087), .ZN(\mult_22/ab[58][45] ) );
  NOR2_X1 U12536 ( .A1(n2661), .A2(n3075), .ZN(\mult_22/ab[56][47] ) );
  NOR2_X1 U12537 ( .A1(n2675), .A2(n3063), .ZN(\mult_22/ab[54][49] ) );
  NOR2_X1 U12538 ( .A1(n2685), .A2(n3051), .ZN(\mult_22/ab[52][51] ) );
  NOR2_X1 U12539 ( .A1(n2695), .A2(n3040), .ZN(\mult_22/ab[50][53] ) );
  NOR2_X1 U12540 ( .A1(n2707), .A2(n3028), .ZN(\mult_22/ab[48][55] ) );
  NOR2_X1 U12541 ( .A1(n2718), .A2(n3016), .ZN(\mult_22/ab[46][57] ) );
  NOR2_X1 U12542 ( .A1(n2726), .A2(n3004), .ZN(\mult_22/ab[44][59] ) );
  NOR2_X1 U12543 ( .A1(n2642), .A2(n3093), .ZN(\mult_22/ab[59][44] ) );
  NOR2_X1 U12544 ( .A1(n2655), .A2(n3081), .ZN(\mult_22/ab[57][46] ) );
  NOR2_X1 U12545 ( .A1(n2667), .A2(n3069), .ZN(\mult_22/ab[55][48] ) );
  NOR2_X1 U12546 ( .A1(n2679), .A2(n3057), .ZN(\mult_22/ab[53][50] ) );
  NOR2_X1 U12547 ( .A1(n2693), .A2(n3045), .ZN(\mult_22/ab[51][52] ) );
  NOR2_X1 U12548 ( .A1(n2701), .A2(n3034), .ZN(\mult_22/ab[49][54] ) );
  NOR2_X1 U12549 ( .A1(n2712), .A2(n3022), .ZN(\mult_22/ab[47][56] ) );
  NOR2_X1 U12550 ( .A1(n2722), .A2(n3010), .ZN(\mult_22/ab[45][58] ) );
  NOR2_X1 U12551 ( .A1(n2733), .A2(n2998), .ZN(\mult_22/ab[43][60] ) );
  NOR2_X1 U12552 ( .A1(n2737), .A2(n3034), .ZN(\mult_22/ab[49][61] ) );
  NOR2_X1 U12553 ( .A1(n2734), .A2(n3040), .ZN(\mult_22/ab[50][60] ) );
  NOR2_X1 U12554 ( .A1(n2727), .A2(n3046), .ZN(\mult_22/ab[51][59] ) );
  NOR2_X1 U12555 ( .A1(n2722), .A2(n3052), .ZN(\mult_22/ab[52][58] ) );
  NOR2_X1 U12556 ( .A1(n2738), .A2(n3040), .ZN(\mult_22/ab[50][61] ) );
  NOR2_X1 U12557 ( .A1(n2718), .A2(n3058), .ZN(\mult_22/ab[53][57] ) );
  NOR2_X1 U12558 ( .A1(n2734), .A2(n3046), .ZN(\mult_22/ab[51][60] ) );
  NOR2_X1 U12559 ( .A1(n2712), .A2(n3064), .ZN(\mult_22/ab[54][56] ) );
  NOR2_X1 U12560 ( .A1(n2728), .A2(n3052), .ZN(\mult_22/ab[52][59] ) );
  NOR2_X1 U12561 ( .A1(n2707), .A2(n3070), .ZN(\mult_22/ab[55][55] ) );
  NOR2_X1 U12562 ( .A1(n2722), .A2(n3058), .ZN(\mult_22/ab[53][58] ) );
  NOR2_X1 U12563 ( .A1(n2701), .A2(n3076), .ZN(\mult_22/ab[56][54] ) );
  NOR2_X1 U12564 ( .A1(n2716), .A2(n3064), .ZN(\mult_22/ab[54][57] ) );
  NOR2_X1 U12565 ( .A1(n2700), .A2(n3082), .ZN(\mult_22/ab[57][53] ) );
  NOR2_X1 U12566 ( .A1(n2712), .A2(n3070), .ZN(\mult_22/ab[55][56] ) );
  NOR2_X1 U12567 ( .A1(n2694), .A2(n3087), .ZN(\mult_22/ab[58][52] ) );
  NOR2_X1 U12568 ( .A1(n2707), .A2(n3076), .ZN(\mult_22/ab[56][55] ) );
  NOR2_X1 U12569 ( .A1(n2685), .A2(n3093), .ZN(\mult_22/ab[59][51] ) );
  NOR2_X1 U12570 ( .A1(n2701), .A2(n3082), .ZN(\mult_22/ab[57][54] ) );
  NOR2_X1 U12571 ( .A1(n2367), .A2(n3088), .ZN(\mult_22/ab[58][53] ) );
  NOR2_X1 U12572 ( .A1(n2694), .A2(n3093), .ZN(\mult_22/ab[59][52] ) );
  NOR2_X1 U12573 ( .A1(n2741), .A2(n2992), .ZN(\mult_22/ab[42][61] ) );
  NOR2_X1 U12574 ( .A1(n2660), .A2(n3099), .ZN(\mult_22/ab[60][47] ) );
  NOR2_X1 U12575 ( .A1(n2652), .A2(n3093), .ZN(\mult_22/ab[59][45] ) );
  NOR2_X1 U12576 ( .A1(n2661), .A2(n3081), .ZN(\mult_22/ab[57][47] ) );
  NOR2_X1 U12577 ( .A1(n2676), .A2(n3069), .ZN(\mult_22/ab[55][49] ) );
  NOR2_X1 U12578 ( .A1(n2685), .A2(n3057), .ZN(\mult_22/ab[53][51] ) );
  NOR2_X1 U12579 ( .A1(n2700), .A2(n3046), .ZN(\mult_22/ab[51][53] ) );
  NOR2_X1 U12580 ( .A1(n2707), .A2(n3034), .ZN(\mult_22/ab[49][55] ) );
  NOR2_X1 U12581 ( .A1(n2716), .A2(n3022), .ZN(\mult_22/ab[47][57] ) );
  NOR2_X1 U12582 ( .A1(n2727), .A2(n3010), .ZN(\mult_22/ab[45][59] ) );
  NOR2_X1 U12583 ( .A1(n2666), .A2(n3099), .ZN(\mult_22/ab[60][48] ) );
  NOR2_X1 U12584 ( .A1(n2654), .A2(n3087), .ZN(\mult_22/ab[58][46] ) );
  NOR2_X1 U12585 ( .A1(n2667), .A2(n3075), .ZN(\mult_22/ab[56][48] ) );
  NOR2_X1 U12586 ( .A1(n2679), .A2(n3063), .ZN(\mult_22/ab[54][50] ) );
  NOR2_X1 U12587 ( .A1(n2693), .A2(n3051), .ZN(\mult_22/ab[52][52] ) );
  NOR2_X1 U12588 ( .A1(n2701), .A2(n3040), .ZN(\mult_22/ab[50][54] ) );
  NOR2_X1 U12589 ( .A1(n2712), .A2(n3028), .ZN(\mult_22/ab[48][56] ) );
  NOR2_X1 U12590 ( .A1(n2722), .A2(n3016), .ZN(\mult_22/ab[46][58] ) );
  NOR2_X1 U12591 ( .A1(n2734), .A2(n3004), .ZN(\mult_22/ab[44][60] ) );
  NOR2_X1 U12592 ( .A1(n2739), .A2(n2998), .ZN(\mult_22/ab[43][61] ) );
  NOR2_X1 U12593 ( .A1(n2685), .A2(n3087), .ZN(\mult_22/ab[58][51] ) );
  NOR2_X1 U12594 ( .A1(n2678), .A2(n3093), .ZN(\mult_22/ab[59][50] ) );
  NOR2_X1 U12595 ( .A1(n2695), .A2(n3076), .ZN(\mult_22/ab[56][53] ) );
  NOR2_X1 U12596 ( .A1(n2694), .A2(n3081), .ZN(\mult_22/ab[57][52] ) );
  NOR2_X1 U12597 ( .A1(n2707), .A2(n3064), .ZN(\mult_22/ab[54][55] ) );
  NOR2_X1 U12598 ( .A1(n2701), .A2(n3070), .ZN(\mult_22/ab[55][54] ) );
  NOR2_X1 U12599 ( .A1(n2716), .A2(n3052), .ZN(\mult_22/ab[52][57] ) );
  NOR2_X1 U12600 ( .A1(n2715), .A2(n3058), .ZN(\mult_22/ab[53][56] ) );
  NOR2_X1 U12601 ( .A1(n2726), .A2(n3040), .ZN(\mult_22/ab[50][59] ) );
  NOR2_X1 U12602 ( .A1(n2722), .A2(n3046), .ZN(\mult_22/ab[51][58] ) );
  NOR2_X1 U12603 ( .A1(n2741), .A2(n3028), .ZN(\mult_22/ab[48][61] ) );
  NOR2_X1 U12604 ( .A1(n2734), .A2(n3034), .ZN(\mult_22/ab[49][60] ) );
  NOR2_X1 U12605 ( .A1(n2661), .A2(n3087), .ZN(\mult_22/ab[58][47] ) );
  NOR2_X1 U12606 ( .A1(n2676), .A2(n3075), .ZN(\mult_22/ab[56][49] ) );
  NOR2_X1 U12607 ( .A1(n2686), .A2(n3063), .ZN(\mult_22/ab[54][51] ) );
  NOR2_X1 U12608 ( .A1(n2367), .A2(n3052), .ZN(\mult_22/ab[52][53] ) );
  NOR2_X1 U12609 ( .A1(n2707), .A2(n3040), .ZN(\mult_22/ab[50][55] ) );
  NOR2_X1 U12610 ( .A1(n2716), .A2(n3028), .ZN(\mult_22/ab[48][57] ) );
  NOR2_X1 U12611 ( .A1(n2728), .A2(n3016), .ZN(\mult_22/ab[46][59] ) );
  NOR2_X1 U12612 ( .A1(n2660), .A2(n3093), .ZN(\mult_22/ab[59][47] ) );
  NOR2_X1 U12613 ( .A1(n2676), .A2(n3081), .ZN(\mult_22/ab[57][49] ) );
  NOR2_X1 U12614 ( .A1(n2685), .A2(n3069), .ZN(\mult_22/ab[55][51] ) );
  NOR2_X1 U12615 ( .A1(n2699), .A2(n3058), .ZN(\mult_22/ab[53][53] ) );
  NOR2_X1 U12616 ( .A1(n2707), .A2(n3046), .ZN(\mult_22/ab[51][55] ) );
  NOR2_X1 U12617 ( .A1(n2718), .A2(n3034), .ZN(\mult_22/ab[49][57] ) );
  NOR2_X1 U12618 ( .A1(n2729), .A2(n3022), .ZN(\mult_22/ab[47][59] ) );
  NOR2_X1 U12619 ( .A1(n2654), .A2(n3093), .ZN(\mult_22/ab[59][46] ) );
  NOR2_X1 U12620 ( .A1(n2667), .A2(n3081), .ZN(\mult_22/ab[57][48] ) );
  NOR2_X1 U12621 ( .A1(n2679), .A2(n3069), .ZN(\mult_22/ab[55][50] ) );
  NOR2_X1 U12622 ( .A1(n2693), .A2(n3057), .ZN(\mult_22/ab[53][52] ) );
  NOR2_X1 U12623 ( .A1(n2701), .A2(n3046), .ZN(\mult_22/ab[51][54] ) );
  NOR2_X1 U12624 ( .A1(n2666), .A2(n3087), .ZN(\mult_22/ab[58][48] ) );
  NOR2_X1 U12625 ( .A1(n2712), .A2(n3034), .ZN(\mult_22/ab[49][56] ) );
  NOR2_X1 U12626 ( .A1(n2679), .A2(n3075), .ZN(\mult_22/ab[56][50] ) );
  NOR2_X1 U12627 ( .A1(n2722), .A2(n3022), .ZN(\mult_22/ab[47][58] ) );
  NOR2_X1 U12628 ( .A1(n2693), .A2(n3063), .ZN(\mult_22/ab[54][52] ) );
  NOR2_X1 U12629 ( .A1(n2701), .A2(n3052), .ZN(\mult_22/ab[52][54] ) );
  NOR2_X1 U12630 ( .A1(n2712), .A2(n3040), .ZN(\mult_22/ab[50][56] ) );
  NOR2_X1 U12631 ( .A1(n2722), .A2(n3028), .ZN(\mult_22/ab[48][58] ) );
  NOR2_X1 U12632 ( .A1(n2737), .A2(n3004), .ZN(\mult_22/ab[44][61] ) );
  NOR2_X1 U12633 ( .A1(n2739), .A2(n3046), .ZN(\mult_22/ab[51][61] ) );
  NOR2_X1 U12634 ( .A1(n2734), .A2(n3052), .ZN(\mult_22/ab[52][60] ) );
  NOR2_X1 U12635 ( .A1(n2729), .A2(n3058), .ZN(\mult_22/ab[53][59] ) );
  NOR2_X1 U12636 ( .A1(n2722), .A2(n3064), .ZN(\mult_22/ab[54][58] ) );
  NOR2_X1 U12637 ( .A1(n2718), .A2(n3070), .ZN(\mult_22/ab[55][57] ) );
  NOR2_X1 U12638 ( .A1(n2715), .A2(n3076), .ZN(\mult_22/ab[56][56] ) );
  NOR2_X1 U12639 ( .A1(n2707), .A2(n3082), .ZN(\mult_22/ab[57][55] ) );
  NOR2_X1 U12640 ( .A1(n2694), .A2(n3099), .ZN(\mult_22/ab[60][52] ) );
  NOR2_X1 U12641 ( .A1(n2738), .A2(n3010), .ZN(\mult_22/ab[45][61] ) );
  NOR2_X1 U12642 ( .A1(n2734), .A2(n3010), .ZN(\mult_22/ab[45][60] ) );
  NOR2_X1 U12643 ( .A1(n2734), .A2(n3016), .ZN(\mult_22/ab[46][60] ) );
  NOR2_X1 U12644 ( .A1(n2676), .A2(n3087), .ZN(\mult_22/ab[58][49] ) );
  NOR2_X1 U12645 ( .A1(n2685), .A2(n3075), .ZN(\mult_22/ab[56][51] ) );
  NOR2_X1 U12646 ( .A1(n2696), .A2(n3064), .ZN(\mult_22/ab[54][53] ) );
  NOR2_X1 U12647 ( .A1(n2707), .A2(n3052), .ZN(\mult_22/ab[52][55] ) );
  NOR2_X1 U12648 ( .A1(n2716), .A2(n3040), .ZN(\mult_22/ab[50][57] ) );
  NOR2_X1 U12649 ( .A1(n2730), .A2(n3028), .ZN(\mult_22/ab[48][59] ) );
  NOR2_X1 U12650 ( .A1(n2666), .A2(n3093), .ZN(\mult_22/ab[59][48] ) );
  NOR2_X1 U12651 ( .A1(n2678), .A2(n3081), .ZN(\mult_22/ab[57][50] ) );
  NOR2_X1 U12652 ( .A1(n2693), .A2(n3069), .ZN(\mult_22/ab[55][52] ) );
  NOR2_X1 U12653 ( .A1(n2701), .A2(n3058), .ZN(\mult_22/ab[53][54] ) );
  NOR2_X1 U12654 ( .A1(n2712), .A2(n3046), .ZN(\mult_22/ab[51][56] ) );
  NOR2_X1 U12655 ( .A1(n2722), .A2(n3034), .ZN(\mult_22/ab[49][58] ) );
  NOR2_X1 U12656 ( .A1(n2734), .A2(n3022), .ZN(\mult_22/ab[47][60] ) );
  NOR2_X1 U12657 ( .A1(n2739), .A2(n3016), .ZN(\mult_22/ab[46][61] ) );
  NOR2_X1 U12658 ( .A1(n2676), .A2(n3093), .ZN(\mult_22/ab[59][49] ) );
  NOR2_X1 U12659 ( .A1(n2685), .A2(n3081), .ZN(\mult_22/ab[57][51] ) );
  NOR2_X1 U12660 ( .A1(n2697), .A2(n3070), .ZN(\mult_22/ab[55][53] ) );
  NOR2_X1 U12661 ( .A1(n2707), .A2(n3058), .ZN(\mult_22/ab[53][55] ) );
  NOR2_X1 U12662 ( .A1(n2718), .A2(n3046), .ZN(\mult_22/ab[51][57] ) );
  NOR2_X1 U12663 ( .A1(n2725), .A2(n3034), .ZN(\mult_22/ab[49][59] ) );
  NOR2_X1 U12664 ( .A1(n2678), .A2(n3087), .ZN(\mult_22/ab[58][50] ) );
  NOR2_X1 U12665 ( .A1(n2694), .A2(n3075), .ZN(\mult_22/ab[56][52] ) );
  NOR2_X1 U12666 ( .A1(n2701), .A2(n3064), .ZN(\mult_22/ab[54][54] ) );
  NOR2_X1 U12667 ( .A1(n2712), .A2(n3052), .ZN(\mult_22/ab[52][56] ) );
  NOR2_X1 U12668 ( .A1(n2722), .A2(n3040), .ZN(\mult_22/ab[50][58] ) );
  NOR2_X1 U12669 ( .A1(n2734), .A2(n3028), .ZN(\mult_22/ab[48][60] ) );
  NOR2_X1 U12670 ( .A1(n2740), .A2(n3022), .ZN(\mult_22/ab[47][61] ) );
  NOR2_X1 U12671 ( .A1(n2738), .A2(n3052), .ZN(\mult_22/ab[52][61] ) );
  NOR2_X1 U12672 ( .A1(n2739), .A2(n3058), .ZN(\mult_22/ab[53][61] ) );
  NOR2_X1 U12673 ( .A1(n2734), .A2(n3058), .ZN(\mult_22/ab[53][60] ) );
  NOR2_X1 U12674 ( .A1(n2734), .A2(n3064), .ZN(\mult_22/ab[54][60] ) );
  NOR2_X1 U12675 ( .A1(n2730), .A2(n3064), .ZN(\mult_22/ab[54][59] ) );
  NOR2_X1 U12676 ( .A1(n2725), .A2(n3070), .ZN(\mult_22/ab[55][59] ) );
  NOR2_X1 U12677 ( .A1(n2723), .A2(n3070), .ZN(\mult_22/ab[55][58] ) );
  NOR2_X1 U12678 ( .A1(n2723), .A2(n3076), .ZN(\mult_22/ab[56][58] ) );
  NOR2_X1 U12679 ( .A1(n2716), .A2(n3076), .ZN(\mult_22/ab[56][57] ) );
  NOR2_X1 U12680 ( .A1(n2740), .A2(n3064), .ZN(\mult_22/ab[54][61] ) );
  NOR2_X1 U12681 ( .A1(n2718), .A2(n3082), .ZN(\mult_22/ab[57][57] ) );
  NOR2_X1 U12682 ( .A1(n2712), .A2(n3082), .ZN(\mult_22/ab[57][56] ) );
  NOR2_X1 U12683 ( .A1(n2741), .A2(n3070), .ZN(\mult_22/ab[55][61] ) );
  NOR2_X1 U12684 ( .A1(n2735), .A2(n3070), .ZN(\mult_22/ab[55][60] ) );
  NOR2_X1 U12685 ( .A1(n2712), .A2(n3088), .ZN(\mult_22/ab[58][56] ) );
  NOR2_X1 U12686 ( .A1(n2735), .A2(n3076), .ZN(\mult_22/ab[56][60] ) );
  NOR2_X1 U12687 ( .A1(n2726), .A2(n3076), .ZN(\mult_22/ab[56][59] ) );
  NOR2_X1 U12688 ( .A1(n2727), .A2(n3082), .ZN(\mult_22/ab[57][59] ) );
  NOR2_X1 U12689 ( .A1(n2723), .A2(n3082), .ZN(\mult_22/ab[57][58] ) );
  NOR2_X1 U12690 ( .A1(n2723), .A2(n3088), .ZN(\mult_22/ab[58][58] ) );
  NOR2_X1 U12691 ( .A1(n2716), .A2(n3088), .ZN(\mult_22/ab[58][57] ) );
  NOR2_X1 U12692 ( .A1(n2737), .A2(n3076), .ZN(\mult_22/ab[56][61] ) );
  NOR2_X1 U12693 ( .A1(n2694), .A2(n3105), .ZN(\mult_22/ab[61][52] ) );
  NOR2_X1 U12694 ( .A1(n2716), .A2(n3094), .ZN(\mult_22/ab[59][57] ) );
  NOR2_X1 U12695 ( .A1(n2715), .A2(n3094), .ZN(\mult_22/ab[59][56] ) );
  NOR2_X1 U12696 ( .A1(n2738), .A2(n3082), .ZN(\mult_22/ab[57][61] ) );
  NOR2_X1 U12697 ( .A1(n2735), .A2(n3082), .ZN(\mult_22/ab[57][60] ) );
  NOR2_X1 U12698 ( .A1(n2694), .A2(n3111), .ZN(\mult_22/ab[62][52] ) );
  NOR2_X1 U12699 ( .A1(n2684), .A2(n3111), .ZN(\mult_22/ab[62][51] ) );
  NOR2_X1 U12700 ( .A1(n2712), .A2(n3100), .ZN(\mult_22/ab[60][56] ) );
  NOR2_X1 U12701 ( .A1(n2739), .A2(n3088), .ZN(\mult_22/ab[58][61] ) );
  NOR2_X1 U12702 ( .A1(n2735), .A2(n3088), .ZN(\mult_22/ab[58][60] ) );
  NOR2_X1 U12703 ( .A1(n2728), .A2(n3088), .ZN(\mult_22/ab[58][59] ) );
  NOR2_X1 U12704 ( .A1(n2740), .A2(n3094), .ZN(\mult_22/ab[59][61] ) );
  NOR2_X1 U12705 ( .A1(n2735), .A2(n3094), .ZN(\mult_22/ab[59][60] ) );
  NOR2_X1 U12706 ( .A1(n2729), .A2(n3094), .ZN(\mult_22/ab[59][59] ) );
  NOR2_X1 U12707 ( .A1(n2723), .A2(n3094), .ZN(\mult_22/ab[59][58] ) );
  NOR2_X1 U12708 ( .A1(n2735), .A2(n3100), .ZN(\mult_22/ab[60][60] ) );
  NOR2_X1 U12709 ( .A1(n2718), .A2(n3100), .ZN(\mult_22/ab[60][57] ) );
  NOR2_X1 U12710 ( .A1(n2730), .A2(n3100), .ZN(\mult_22/ab[60][59] ) );
  NOR2_X1 U12711 ( .A1(n2723), .A2(n3100), .ZN(\mult_22/ab[60][58] ) );
  NOR2_X1 U12712 ( .A1(n2712), .A2(n3106), .ZN(\mult_22/ab[61][56] ) );
  NOR2_X1 U12713 ( .A1(n2725), .A2(n3106), .ZN(\mult_22/ab[61][59] ) );
  NOR2_X1 U12714 ( .A1(n2718), .A2(n3106), .ZN(\mult_22/ab[61][57] ) );
  NOR2_X1 U12715 ( .A1(n2723), .A2(n3106), .ZN(\mult_22/ab[61][58] ) );
  NOR2_X1 U12716 ( .A1(n2715), .A2(n3112), .ZN(\mult_22/ab[62][56] ) );
  NOR2_X1 U12717 ( .A1(n2723), .A2(n3112), .ZN(\mult_22/ab[62][58] ) );
  NOR2_X1 U12718 ( .A1(n2718), .A2(n3112), .ZN(\mult_22/ab[62][57] ) );
  NOR2_X1 U12719 ( .A1(n2741), .A2(n3100), .ZN(\mult_22/ab[60][61] ) );
  NOR2_X1 U12720 ( .A1(n2735), .A2(n3106), .ZN(\mult_22/ab[61][60] ) );
  NOR2_X1 U12721 ( .A1(n2726), .A2(n3112), .ZN(\mult_22/ab[62][59] ) );
  NOR2_X1 U12722 ( .A1(n2737), .A2(n3106), .ZN(\mult_22/ab[61][61] ) );
  NOR2_X1 U12723 ( .A1(n2735), .A2(n3112), .ZN(\mult_22/ab[62][60] ) );
  NOR2_X1 U12724 ( .A1(n2589), .A2(n3110), .ZN(\mult_22/ab[62][35] ) );
  NOR2_X1 U12725 ( .A1(n2583), .A2(n3110), .ZN(\mult_22/ab[62][34] ) );
  NOR2_X1 U12726 ( .A1(n2577), .A2(n3110), .ZN(\mult_22/ab[62][33] ) );
  NOR2_X1 U12727 ( .A1(n2595), .A2(n3104), .ZN(\mult_22/ab[61][36] ) );
  NOR2_X1 U12728 ( .A1(n2589), .A2(n3104), .ZN(\mult_22/ab[61][35] ) );
  NOR2_X1 U12729 ( .A1(n2583), .A2(n3104), .ZN(\mult_22/ab[61][34] ) );
  NOR2_X1 U12730 ( .A1(n2577), .A2(n3104), .ZN(\mult_22/ab[61][33] ) );
  NOR2_X1 U12731 ( .A1(n2595), .A2(n3098), .ZN(\mult_22/ab[60][36] ) );
  NOR2_X1 U12732 ( .A1(n2628), .A2(n3104), .ZN(\mult_22/ab[61][41] ) );
  NOR2_X1 U12733 ( .A1(n2589), .A2(n3098), .ZN(\mult_22/ab[60][35] ) );
  NOR2_X1 U12734 ( .A1(n2577), .A2(n3098), .ZN(\mult_22/ab[60][33] ) );
  NOR2_X1 U12735 ( .A1(n2583), .A2(n3098), .ZN(\mult_22/ab[60][34] ) );
  NOR2_X1 U12736 ( .A1(n2595), .A2(n3092), .ZN(\mult_22/ab[59][36] ) );
  NOR2_X1 U12737 ( .A1(n2589), .A2(n3092), .ZN(\mult_22/ab[59][35] ) );
  NOR2_X1 U12738 ( .A1(n2583), .A2(n3092), .ZN(\mult_22/ab[59][34] ) );
  NOR2_X1 U12739 ( .A1(n2583), .A2(n3086), .ZN(\mult_22/ab[58][34] ) );
  NOR2_X1 U12740 ( .A1(n2607), .A2(n3086), .ZN(\mult_22/ab[58][38] ) );
  NOR2_X1 U12741 ( .A1(n2595), .A2(n3086), .ZN(\mult_22/ab[58][36] ) );
  NOR2_X1 U12742 ( .A1(n2589), .A2(n3086), .ZN(\mult_22/ab[58][35] ) );
  NOR2_X1 U12743 ( .A1(n2590), .A2(n3080), .ZN(\mult_22/ab[57][35] ) );
  NOR2_X1 U12744 ( .A1(n2608), .A2(n3080), .ZN(\mult_22/ab[57][38] ) );
  NOR2_X1 U12745 ( .A1(n2613), .A2(n3080), .ZN(\mult_22/ab[57][39] ) );
  NOR2_X1 U12746 ( .A1(n2596), .A2(n3080), .ZN(\mult_22/ab[57][36] ) );
  NOR2_X1 U12747 ( .A1(n2608), .A2(n3062), .ZN(\mult_22/ab[54][38] ) );
  NOR2_X1 U12748 ( .A1(n2608), .A2(n3068), .ZN(\mult_22/ab[55][38] ) );
  NOR2_X1 U12749 ( .A1(n2608), .A2(n3074), .ZN(\mult_22/ab[56][38] ) );
  NOR2_X1 U12750 ( .A1(n2596), .A2(n3074), .ZN(\mult_22/ab[56][36] ) );
  NOR2_X1 U12751 ( .A1(n2627), .A2(n3044), .ZN(\mult_22/ab[51][41] ) );
  NOR2_X1 U12752 ( .A1(n2662), .A2(n3009), .ZN(\mult_22/ab[45][47] ) );
  NOR2_X1 U12753 ( .A1(n2651), .A2(n3021), .ZN(\mult_22/ab[47][45] ) );
  NOR2_X1 U12754 ( .A1(n2639), .A2(n3033), .ZN(\mult_22/ab[49][43] ) );
  NOR2_X1 U12755 ( .A1(n2651), .A2(n3027), .ZN(\mult_22/ab[48][45] ) );
  NOR2_X1 U12756 ( .A1(n2613), .A2(n3056), .ZN(\mult_22/ab[53][39] ) );
  NOR2_X1 U12757 ( .A1(n2639), .A2(n3039), .ZN(\mult_22/ab[50][43] ) );
  NOR2_X1 U12758 ( .A1(n2639), .A2(n3045), .ZN(\mult_22/ab[51][43] ) );
  NOR2_X1 U12759 ( .A1(n2627), .A2(n3050), .ZN(\mult_22/ab[52][41] ) );
  NOR2_X1 U12760 ( .A1(n2627), .A2(n3056), .ZN(\mult_22/ab[53][41] ) );
  NOR2_X1 U12761 ( .A1(n2613), .A2(n3062), .ZN(\mult_22/ab[54][39] ) );
  NOR2_X1 U12762 ( .A1(n2613), .A2(n3068), .ZN(\mult_22/ab[55][39] ) );
  NOR2_X1 U12763 ( .A1(n2627), .A2(n3062), .ZN(\mult_22/ab[54][41] ) );
  NOR2_X1 U12764 ( .A1(n2613), .A2(n3074), .ZN(\mult_22/ab[56][39] ) );
  AND3_X1 U12765 ( .A1(\mult_22/CARRYB[63][53] ), .A2(n1330), .A3(
        \mult_22/SUMB[63][54] ), .ZN(n1326) );
  NOR2_X1 U12766 ( .A1(n2748), .A2(n3112), .ZN(\mult_22/ab[62][63] ) );
  NOR2_X1 U12767 ( .A1(n2744), .A2(n3118), .ZN(\mult_22/ab[63][62] ) );
  NOR2_X1 U12768 ( .A1(n2739), .A2(n3118), .ZN(\mult_22/ab[63][61] ) );
  NOR2_X1 U12769 ( .A1(n2748), .A2(n3100), .ZN(\mult_22/ab[60][63] ) );
  NOR2_X1 U12770 ( .A1(n2747), .A2(n3106), .ZN(\mult_22/ab[61][62] ) );
  NOR2_X1 U12771 ( .A1(n2748), .A2(n3106), .ZN(\mult_22/ab[61][63] ) );
  NOR2_X1 U12772 ( .A1(n2743), .A2(n3112), .ZN(\mult_22/ab[62][62] ) );
  NOR2_X1 U12773 ( .A1(n2738), .A2(n3112), .ZN(\mult_22/ab[62][61] ) );
  INV_X1 U12774 ( .A(n3523), .ZN(n3516) );
  INV_X1 U12775 ( .A(n3534), .ZN(n3527) );
  NOR2_X1 U12776 ( .A1(n3417), .A2(n3395), .ZN(\mult_20/ab[31][7] ) );
  NOR2_X1 U12777 ( .A1(n3231), .A2(n3209), .ZN(\mult_19/ab[31][7] ) );
  NOR2_X1 U12778 ( .A1(n3429), .A2(n3393), .ZN(\mult_20/ab[31][11] ) );
  NOR2_X1 U12779 ( .A1(n3243), .A2(n3207), .ZN(\mult_19/ab[31][11] ) );
  NOR2_X1 U12780 ( .A1(n3219), .A2(n3209), .ZN(\mult_19/ab[31][3] ) );
  NOR2_X1 U12781 ( .A1(n3420), .A2(n3395), .ZN(\mult_20/ab[31][8] ) );
  NOR2_X1 U12782 ( .A1(n3234), .A2(n3209), .ZN(\mult_19/ab[31][8] ) );
  NOR2_X1 U12783 ( .A1(n3432), .A2(n3393), .ZN(\mult_20/ab[31][12] ) );
  NOR2_X1 U12784 ( .A1(n3246), .A2(n3207), .ZN(\mult_19/ab[31][12] ) );
  NOR2_X1 U12785 ( .A1(n3435), .A2(n3393), .ZN(\mult_20/ab[31][13] ) );
  NOR2_X1 U12786 ( .A1(n3249), .A2(n3207), .ZN(\mult_19/ab[31][13] ) );
  NOR2_X1 U12787 ( .A1(n3426), .A2(n3393), .ZN(\mult_20/ab[31][10] ) );
  NOR2_X1 U12788 ( .A1(n3240), .A2(n3207), .ZN(\mult_19/ab[31][10] ) );
  NOR2_X1 U12789 ( .A1(n3397), .A2(n3393), .ZN(\mult_20/ab[31][0] ) );
  NOR2_X1 U12790 ( .A1(n3211), .A2(n3207), .ZN(\mult_19/ab[31][0] ) );
  NOR2_X1 U12791 ( .A1(n3411), .A2(n3395), .ZN(\mult_20/ab[31][5] ) );
  NOR2_X1 U12792 ( .A1(n3225), .A2(n3209), .ZN(\mult_19/ab[31][5] ) );
  NOR2_X1 U12793 ( .A1(n3222), .A2(n3209), .ZN(\mult_19/ab[31][4] ) );
  NOR2_X1 U12794 ( .A1(n3405), .A2(n3395), .ZN(\mult_20/ab[31][3] ) );
  NOR2_X1 U12795 ( .A1(n3408), .A2(n3395), .ZN(\mult_20/ab[31][4] ) );
  NOR2_X1 U12796 ( .A1(n3414), .A2(n3395), .ZN(\mult_20/ab[31][6] ) );
  NOR2_X1 U12797 ( .A1(n3216), .A2(n3208), .ZN(\mult_19/ab[31][2] ) );
  NOR2_X1 U12798 ( .A1(n3228), .A2(n3209), .ZN(\mult_19/ab[31][6] ) );
  NOR2_X1 U12799 ( .A1(n3423), .A2(n3395), .ZN(\mult_20/ab[31][9] ) );
  NOR2_X1 U12800 ( .A1(n3237), .A2(n3209), .ZN(\mult_19/ab[31][9] ) );
  NOR2_X1 U12801 ( .A1(n3213), .A2(n3207), .ZN(\mult_19/ab[31][1] ) );
  NOR2_X1 U12802 ( .A1(n3402), .A2(n3394), .ZN(\mult_20/ab[31][2] ) );
  NOR2_X1 U12803 ( .A1(n3399), .A2(n3393), .ZN(\mult_20/ab[31][1] ) );
  NOR2_X1 U12804 ( .A1(n3490), .A2(n3308), .ZN(\mult_20/ab[2][31] ) );
  NOR2_X1 U12805 ( .A1(n3486), .A2(n3310), .ZN(\mult_20/ab[3][30] ) );
  NOR2_X1 U12806 ( .A1(n3304), .A2(n3122), .ZN(\mult_19/ab[2][31] ) );
  NOR2_X1 U12807 ( .A1(n3300), .A2(n3124), .ZN(\mult_19/ab[3][30] ) );
  NOR2_X1 U12808 ( .A1(n3491), .A2(n3311), .ZN(\mult_20/ab[3][31] ) );
  NOR2_X1 U12809 ( .A1(n3486), .A2(n3313), .ZN(\mult_20/ab[4][30] ) );
  NOR2_X1 U12810 ( .A1(n3305), .A2(n3125), .ZN(\mult_19/ab[3][31] ) );
  NOR2_X1 U12811 ( .A1(n3300), .A2(n3127), .ZN(\mult_19/ab[4][30] ) );
  NOR2_X1 U12812 ( .A1(n3491), .A2(n3314), .ZN(\mult_20/ab[4][31] ) );
  NOR2_X1 U12813 ( .A1(n3486), .A2(n3316), .ZN(\mult_20/ab[5][30] ) );
  NOR2_X1 U12814 ( .A1(n3305), .A2(n3128), .ZN(\mult_19/ab[4][31] ) );
  NOR2_X1 U12815 ( .A1(n3300), .A2(n3130), .ZN(\mult_19/ab[5][30] ) );
  NOR2_X1 U12816 ( .A1(n3491), .A2(n3317), .ZN(\mult_20/ab[5][31] ) );
  NOR2_X1 U12817 ( .A1(n3486), .A2(n3319), .ZN(\mult_20/ab[6][30] ) );
  NOR2_X1 U12818 ( .A1(n3305), .A2(n3131), .ZN(\mult_19/ab[5][31] ) );
  NOR2_X1 U12819 ( .A1(n3300), .A2(n3133), .ZN(\mult_19/ab[6][30] ) );
  NOR2_X1 U12820 ( .A1(n3491), .A2(n3320), .ZN(\mult_20/ab[6][31] ) );
  NOR2_X1 U12821 ( .A1(n3486), .A2(n3322), .ZN(\mult_20/ab[7][30] ) );
  NOR2_X1 U12822 ( .A1(n3305), .A2(n3134), .ZN(\mult_19/ab[6][31] ) );
  NOR2_X1 U12823 ( .A1(n3300), .A2(n3136), .ZN(\mult_19/ab[7][30] ) );
  NOR2_X1 U12824 ( .A1(n3491), .A2(n3323), .ZN(\mult_20/ab[7][31] ) );
  NOR2_X1 U12825 ( .A1(n3486), .A2(n3325), .ZN(\mult_20/ab[8][30] ) );
  NOR2_X1 U12826 ( .A1(n3305), .A2(n3137), .ZN(\mult_19/ab[7][31] ) );
  NOR2_X1 U12827 ( .A1(n3300), .A2(n3139), .ZN(\mult_19/ab[8][30] ) );
  NOR2_X1 U12828 ( .A1(n3491), .A2(n3326), .ZN(\mult_20/ab[8][31] ) );
  NOR2_X1 U12829 ( .A1(n3486), .A2(n3328), .ZN(\mult_20/ab[9][30] ) );
  NOR2_X1 U12830 ( .A1(n3305), .A2(n3140), .ZN(\mult_19/ab[8][31] ) );
  NOR2_X1 U12831 ( .A1(n3300), .A2(n3142), .ZN(\mult_19/ab[9][30] ) );
  NOR2_X1 U12832 ( .A1(n3489), .A2(n3329), .ZN(\mult_20/ab[9][31] ) );
  NOR2_X1 U12833 ( .A1(n3488), .A2(n3331), .ZN(\mult_20/ab[10][30] ) );
  NOR2_X1 U12834 ( .A1(n3303), .A2(n3143), .ZN(\mult_19/ab[9][31] ) );
  NOR2_X1 U12835 ( .A1(n3302), .A2(n3145), .ZN(\mult_19/ab[10][30] ) );
  NOR2_X1 U12836 ( .A1(n3490), .A2(n3332), .ZN(\mult_20/ab[10][31] ) );
  NOR2_X1 U12837 ( .A1(n3488), .A2(n3334), .ZN(\mult_20/ab[11][30] ) );
  NOR2_X1 U12838 ( .A1(n3304), .A2(n3146), .ZN(\mult_19/ab[10][31] ) );
  NOR2_X1 U12839 ( .A1(n3302), .A2(n3148), .ZN(\mult_19/ab[11][30] ) );
  NOR2_X1 U12840 ( .A1(n3489), .A2(n3335), .ZN(\mult_20/ab[11][31] ) );
  NOR2_X1 U12841 ( .A1(n3488), .A2(n3337), .ZN(\mult_20/ab[12][30] ) );
  NOR2_X1 U12842 ( .A1(n3303), .A2(n3149), .ZN(\mult_19/ab[11][31] ) );
  NOR2_X1 U12843 ( .A1(n3302), .A2(n3151), .ZN(\mult_19/ab[12][30] ) );
  NOR2_X1 U12844 ( .A1(n3488), .A2(n3340), .ZN(\mult_20/ab[13][30] ) );
  NOR2_X1 U12845 ( .A1(n3489), .A2(n3338), .ZN(\mult_20/ab[12][31] ) );
  NOR2_X1 U12846 ( .A1(n3302), .A2(n3154), .ZN(\mult_19/ab[13][30] ) );
  NOR2_X1 U12847 ( .A1(n3303), .A2(n3152), .ZN(\mult_19/ab[12][31] ) );
  NOR2_X1 U12848 ( .A1(n3484), .A2(n3310), .ZN(\mult_20/ab[3][29] ) );
  NOR2_X1 U12849 ( .A1(n3480), .A2(n3310), .ZN(\mult_20/ab[3][28] ) );
  NOR2_X1 U12850 ( .A1(n3477), .A2(n3310), .ZN(\mult_20/ab[3][27] ) );
  NOR2_X1 U12851 ( .A1(n3474), .A2(n3310), .ZN(\mult_20/ab[3][26] ) );
  NOR2_X1 U12852 ( .A1(n3471), .A2(n3310), .ZN(\mult_20/ab[3][25] ) );
  NOR2_X1 U12853 ( .A1(n3468), .A2(n3310), .ZN(\mult_20/ab[3][24] ) );
  NOR2_X1 U12854 ( .A1(n3465), .A2(n3310), .ZN(\mult_20/ab[3][23] ) );
  NOR2_X1 U12855 ( .A1(n3462), .A2(n3310), .ZN(\mult_20/ab[3][22] ) );
  NOR2_X1 U12856 ( .A1(n3459), .A2(n3310), .ZN(\mult_20/ab[3][21] ) );
  NOR2_X1 U12857 ( .A1(n3453), .A2(n3309), .ZN(\mult_20/ab[3][19] ) );
  NOR2_X1 U12858 ( .A1(n3447), .A2(n3309), .ZN(\mult_20/ab[3][17] ) );
  NOR2_X1 U12859 ( .A1(n3441), .A2(n3309), .ZN(\mult_20/ab[3][15] ) );
  NOR2_X1 U12860 ( .A1(n3435), .A2(n3309), .ZN(\mult_20/ab[3][13] ) );
  NOR2_X1 U12861 ( .A1(n3429), .A2(n3309), .ZN(\mult_20/ab[3][11] ) );
  NOR2_X1 U12862 ( .A1(n3298), .A2(n3124), .ZN(\mult_19/ab[3][29] ) );
  NOR2_X1 U12863 ( .A1(n3294), .A2(n3124), .ZN(\mult_19/ab[3][28] ) );
  NOR2_X1 U12864 ( .A1(n3291), .A2(n3124), .ZN(\mult_19/ab[3][27] ) );
  NOR2_X1 U12865 ( .A1(n3288), .A2(n3124), .ZN(\mult_19/ab[3][26] ) );
  NOR2_X1 U12866 ( .A1(n3285), .A2(n3124), .ZN(\mult_19/ab[3][25] ) );
  NOR2_X1 U12867 ( .A1(n3282), .A2(n3124), .ZN(\mult_19/ab[3][24] ) );
  NOR2_X1 U12868 ( .A1(n3279), .A2(n3124), .ZN(\mult_19/ab[3][23] ) );
  NOR2_X1 U12869 ( .A1(n3273), .A2(n3124), .ZN(\mult_19/ab[3][21] ) );
  NOR2_X1 U12870 ( .A1(n3270), .A2(n3124), .ZN(\mult_19/ab[3][20] ) );
  NOR2_X1 U12871 ( .A1(n3267), .A2(n3123), .ZN(\mult_19/ab[3][19] ) );
  NOR2_X1 U12872 ( .A1(n3264), .A2(n3123), .ZN(\mult_19/ab[3][18] ) );
  NOR2_X1 U12873 ( .A1(n3261), .A2(n3123), .ZN(\mult_19/ab[3][17] ) );
  NOR2_X1 U12874 ( .A1(n3258), .A2(n3123), .ZN(\mult_19/ab[3][16] ) );
  NOR2_X1 U12875 ( .A1(n3255), .A2(n3123), .ZN(\mult_19/ab[3][15] ) );
  NOR2_X1 U12876 ( .A1(n3252), .A2(n3123), .ZN(\mult_19/ab[3][14] ) );
  NOR2_X1 U12877 ( .A1(n3249), .A2(n3123), .ZN(\mult_19/ab[3][13] ) );
  NOR2_X1 U12878 ( .A1(n3246), .A2(n3123), .ZN(\mult_19/ab[3][12] ) );
  NOR2_X1 U12879 ( .A1(n3243), .A2(n3123), .ZN(\mult_19/ab[3][11] ) );
  NOR2_X1 U12880 ( .A1(n3240), .A2(n3123), .ZN(\mult_19/ab[3][10] ) );
  NOR2_X1 U12881 ( .A1(n3483), .A2(n3313), .ZN(\mult_20/ab[4][29] ) );
  NOR2_X1 U12882 ( .A1(n3480), .A2(n3313), .ZN(\mult_20/ab[4][28] ) );
  NOR2_X1 U12883 ( .A1(n3477), .A2(n3313), .ZN(\mult_20/ab[4][27] ) );
  NOR2_X1 U12884 ( .A1(n3474), .A2(n3313), .ZN(\mult_20/ab[4][26] ) );
  NOR2_X1 U12885 ( .A1(n3471), .A2(n3313), .ZN(\mult_20/ab[4][25] ) );
  NOR2_X1 U12886 ( .A1(n3468), .A2(n3313), .ZN(\mult_20/ab[4][24] ) );
  NOR2_X1 U12887 ( .A1(n3465), .A2(n3313), .ZN(\mult_20/ab[4][23] ) );
  NOR2_X1 U12888 ( .A1(n3462), .A2(n3313), .ZN(\mult_20/ab[4][22] ) );
  NOR2_X1 U12889 ( .A1(n3459), .A2(n3313), .ZN(\mult_20/ab[4][21] ) );
  NOR2_X1 U12890 ( .A1(n3456), .A2(n3313), .ZN(\mult_20/ab[4][20] ) );
  NOR2_X1 U12891 ( .A1(n3453), .A2(n3312), .ZN(\mult_20/ab[4][19] ) );
  NOR2_X1 U12892 ( .A1(n3447), .A2(n3312), .ZN(\mult_20/ab[4][17] ) );
  NOR2_X1 U12893 ( .A1(n3441), .A2(n3312), .ZN(\mult_20/ab[4][15] ) );
  NOR2_X1 U12894 ( .A1(n3435), .A2(n3312), .ZN(\mult_20/ab[4][13] ) );
  NOR2_X1 U12895 ( .A1(n3429), .A2(n3312), .ZN(\mult_20/ab[4][11] ) );
  NOR2_X1 U12896 ( .A1(n3297), .A2(n3127), .ZN(\mult_19/ab[4][29] ) );
  NOR2_X1 U12897 ( .A1(n3294), .A2(n3127), .ZN(\mult_19/ab[4][28] ) );
  NOR2_X1 U12898 ( .A1(n3291), .A2(n3127), .ZN(\mult_19/ab[4][27] ) );
  NOR2_X1 U12899 ( .A1(n3288), .A2(n3127), .ZN(\mult_19/ab[4][26] ) );
  NOR2_X1 U12900 ( .A1(n3285), .A2(n3127), .ZN(\mult_19/ab[4][25] ) );
  NOR2_X1 U12901 ( .A1(n3282), .A2(n3127), .ZN(\mult_19/ab[4][24] ) );
  NOR2_X1 U12902 ( .A1(n3279), .A2(n3127), .ZN(\mult_19/ab[4][23] ) );
  NOR2_X1 U12903 ( .A1(n3276), .A2(n3127), .ZN(\mult_19/ab[4][22] ) );
  NOR2_X1 U12904 ( .A1(n3273), .A2(n3127), .ZN(\mult_19/ab[4][21] ) );
  NOR2_X1 U12905 ( .A1(n3483), .A2(n3316), .ZN(\mult_20/ab[5][29] ) );
  NOR2_X1 U12906 ( .A1(n3480), .A2(n3316), .ZN(\mult_20/ab[5][28] ) );
  NOR2_X1 U12907 ( .A1(n3477), .A2(n3316), .ZN(\mult_20/ab[5][27] ) );
  NOR2_X1 U12908 ( .A1(n3474), .A2(n3316), .ZN(\mult_20/ab[5][26] ) );
  NOR2_X1 U12909 ( .A1(n3471), .A2(n3316), .ZN(\mult_20/ab[5][25] ) );
  NOR2_X1 U12910 ( .A1(n3468), .A2(n3316), .ZN(\mult_20/ab[5][24] ) );
  NOR2_X1 U12911 ( .A1(n3465), .A2(n3316), .ZN(\mult_20/ab[5][23] ) );
  NOR2_X1 U12912 ( .A1(n3462), .A2(n3316), .ZN(\mult_20/ab[5][22] ) );
  NOR2_X1 U12913 ( .A1(n3459), .A2(n3316), .ZN(\mult_20/ab[5][21] ) );
  NOR2_X1 U12914 ( .A1(n3453), .A2(n3315), .ZN(\mult_20/ab[5][19] ) );
  NOR2_X1 U12915 ( .A1(n3447), .A2(n3315), .ZN(\mult_20/ab[5][17] ) );
  NOR2_X1 U12916 ( .A1(n3441), .A2(n3315), .ZN(\mult_20/ab[5][15] ) );
  NOR2_X1 U12917 ( .A1(n3435), .A2(n3315), .ZN(\mult_20/ab[5][13] ) );
  NOR2_X1 U12918 ( .A1(n3429), .A2(n3315), .ZN(\mult_20/ab[5][11] ) );
  NOR2_X1 U12919 ( .A1(n3297), .A2(n3130), .ZN(\mult_19/ab[5][29] ) );
  NOR2_X1 U12920 ( .A1(n3294), .A2(n3130), .ZN(\mult_19/ab[5][28] ) );
  NOR2_X1 U12921 ( .A1(n3291), .A2(n3130), .ZN(\mult_19/ab[5][27] ) );
  NOR2_X1 U12922 ( .A1(n3288), .A2(n3130), .ZN(\mult_19/ab[5][26] ) );
  NOR2_X1 U12923 ( .A1(n3285), .A2(n3130), .ZN(\mult_19/ab[5][25] ) );
  NOR2_X1 U12924 ( .A1(n3282), .A2(n3130), .ZN(\mult_19/ab[5][24] ) );
  NOR2_X1 U12925 ( .A1(n3279), .A2(n3130), .ZN(\mult_19/ab[5][23] ) );
  NOR2_X1 U12926 ( .A1(n3276), .A2(n3130), .ZN(\mult_19/ab[5][22] ) );
  NOR2_X1 U12927 ( .A1(n3267), .A2(n3129), .ZN(\mult_19/ab[5][19] ) );
  NOR2_X1 U12928 ( .A1(n3264), .A2(n3129), .ZN(\mult_19/ab[5][18] ) );
  NOR2_X1 U12929 ( .A1(n3261), .A2(n3129), .ZN(\mult_19/ab[5][17] ) );
  NOR2_X1 U12930 ( .A1(n3258), .A2(n3129), .ZN(\mult_19/ab[5][16] ) );
  NOR2_X1 U12931 ( .A1(n3255), .A2(n3129), .ZN(\mult_19/ab[5][15] ) );
  NOR2_X1 U12932 ( .A1(n3252), .A2(n3129), .ZN(\mult_19/ab[5][14] ) );
  NOR2_X1 U12933 ( .A1(n3249), .A2(n3129), .ZN(\mult_19/ab[5][13] ) );
  NOR2_X1 U12934 ( .A1(n3246), .A2(n3129), .ZN(\mult_19/ab[5][12] ) );
  NOR2_X1 U12935 ( .A1(n3243), .A2(n3129), .ZN(\mult_19/ab[5][11] ) );
  NOR2_X1 U12936 ( .A1(n3240), .A2(n3129), .ZN(\mult_19/ab[5][10] ) );
  NOR2_X1 U12937 ( .A1(n3483), .A2(n3319), .ZN(\mult_20/ab[6][29] ) );
  NOR2_X1 U12938 ( .A1(n3480), .A2(n3319), .ZN(\mult_20/ab[6][28] ) );
  NOR2_X1 U12939 ( .A1(n3477), .A2(n3319), .ZN(\mult_20/ab[6][27] ) );
  NOR2_X1 U12940 ( .A1(n3474), .A2(n3319), .ZN(\mult_20/ab[6][26] ) );
  NOR2_X1 U12941 ( .A1(n3471), .A2(n3319), .ZN(\mult_20/ab[6][25] ) );
  NOR2_X1 U12942 ( .A1(n3468), .A2(n3319), .ZN(\mult_20/ab[6][24] ) );
  NOR2_X1 U12943 ( .A1(n3465), .A2(n3319), .ZN(\mult_20/ab[6][23] ) );
  NOR2_X1 U12944 ( .A1(n3462), .A2(n3319), .ZN(\mult_20/ab[6][22] ) );
  NOR2_X1 U12945 ( .A1(n3459), .A2(n3319), .ZN(\mult_20/ab[6][21] ) );
  NOR2_X1 U12946 ( .A1(n3456), .A2(n3319), .ZN(\mult_20/ab[6][20] ) );
  NOR2_X1 U12947 ( .A1(n3453), .A2(n3318), .ZN(\mult_20/ab[6][19] ) );
  NOR2_X1 U12948 ( .A1(n3447), .A2(n3318), .ZN(\mult_20/ab[6][17] ) );
  NOR2_X1 U12949 ( .A1(n3441), .A2(n3318), .ZN(\mult_20/ab[6][15] ) );
  NOR2_X1 U12950 ( .A1(n3435), .A2(n3318), .ZN(\mult_20/ab[6][13] ) );
  NOR2_X1 U12951 ( .A1(n3429), .A2(n3318), .ZN(\mult_20/ab[6][11] ) );
  NOR2_X1 U12952 ( .A1(n3297), .A2(n3133), .ZN(\mult_19/ab[6][29] ) );
  NOR2_X1 U12953 ( .A1(n3294), .A2(n3133), .ZN(\mult_19/ab[6][28] ) );
  NOR2_X1 U12954 ( .A1(n3291), .A2(n3133), .ZN(\mult_19/ab[6][27] ) );
  NOR2_X1 U12955 ( .A1(n3288), .A2(n3133), .ZN(\mult_19/ab[6][26] ) );
  NOR2_X1 U12956 ( .A1(n3285), .A2(n3133), .ZN(\mult_19/ab[6][25] ) );
  NOR2_X1 U12957 ( .A1(n3282), .A2(n3133), .ZN(\mult_19/ab[6][24] ) );
  NOR2_X1 U12958 ( .A1(n3279), .A2(n3133), .ZN(\mult_19/ab[6][23] ) );
  NOR2_X1 U12959 ( .A1(n3276), .A2(n3133), .ZN(\mult_19/ab[6][22] ) );
  NOR2_X1 U12960 ( .A1(n3273), .A2(n3133), .ZN(\mult_19/ab[6][21] ) );
  NOR2_X1 U12961 ( .A1(n3270), .A2(n3133), .ZN(\mult_19/ab[6][20] ) );
  NOR2_X1 U12962 ( .A1(n3267), .A2(n3132), .ZN(\mult_19/ab[6][19] ) );
  NOR2_X1 U12963 ( .A1(n3483), .A2(n3322), .ZN(\mult_20/ab[7][29] ) );
  NOR2_X1 U12964 ( .A1(n3480), .A2(n3322), .ZN(\mult_20/ab[7][28] ) );
  NOR2_X1 U12965 ( .A1(n3477), .A2(n3322), .ZN(\mult_20/ab[7][27] ) );
  NOR2_X1 U12966 ( .A1(n3474), .A2(n3322), .ZN(\mult_20/ab[7][26] ) );
  NOR2_X1 U12967 ( .A1(n3471), .A2(n3322), .ZN(\mult_20/ab[7][25] ) );
  NOR2_X1 U12968 ( .A1(n3468), .A2(n3322), .ZN(\mult_20/ab[7][24] ) );
  NOR2_X1 U12969 ( .A1(n3465), .A2(n3322), .ZN(\mult_20/ab[7][23] ) );
  NOR2_X1 U12970 ( .A1(n3462), .A2(n3322), .ZN(\mult_20/ab[7][22] ) );
  NOR2_X1 U12971 ( .A1(n3459), .A2(n3322), .ZN(\mult_20/ab[7][21] ) );
  NOR2_X1 U12972 ( .A1(n3456), .A2(n3322), .ZN(\mult_20/ab[7][20] ) );
  NOR2_X1 U12973 ( .A1(n3453), .A2(n3321), .ZN(\mult_20/ab[7][19] ) );
  NOR2_X1 U12974 ( .A1(n3450), .A2(n3321), .ZN(\mult_20/ab[7][18] ) );
  NOR2_X1 U12975 ( .A1(n3447), .A2(n3321), .ZN(\mult_20/ab[7][17] ) );
  NOR2_X1 U12976 ( .A1(n3441), .A2(n3321), .ZN(\mult_20/ab[7][15] ) );
  NOR2_X1 U12977 ( .A1(n3435), .A2(n3321), .ZN(\mult_20/ab[7][13] ) );
  NOR2_X1 U12978 ( .A1(n3429), .A2(n3321), .ZN(\mult_20/ab[7][11] ) );
  NOR2_X1 U12979 ( .A1(n3297), .A2(n3136), .ZN(\mult_19/ab[7][29] ) );
  NOR2_X1 U12980 ( .A1(n3294), .A2(n3136), .ZN(\mult_19/ab[7][28] ) );
  NOR2_X1 U12981 ( .A1(n3291), .A2(n3136), .ZN(\mult_19/ab[7][27] ) );
  NOR2_X1 U12982 ( .A1(n3288), .A2(n3136), .ZN(\mult_19/ab[7][26] ) );
  NOR2_X1 U12983 ( .A1(n3285), .A2(n3136), .ZN(\mult_19/ab[7][25] ) );
  NOR2_X1 U12984 ( .A1(n3282), .A2(n3136), .ZN(\mult_19/ab[7][24] ) );
  NOR2_X1 U12985 ( .A1(n3279), .A2(n3136), .ZN(\mult_19/ab[7][23] ) );
  NOR2_X1 U12986 ( .A1(n3276), .A2(n3136), .ZN(\mult_19/ab[7][22] ) );
  NOR2_X1 U12987 ( .A1(n3273), .A2(n3136), .ZN(\mult_19/ab[7][21] ) );
  NOR2_X1 U12988 ( .A1(n3270), .A2(n3136), .ZN(\mult_19/ab[7][20] ) );
  NOR2_X1 U12989 ( .A1(n3267), .A2(n3135), .ZN(\mult_19/ab[7][19] ) );
  NOR2_X1 U12990 ( .A1(n3261), .A2(n3135), .ZN(\mult_19/ab[7][17] ) );
  NOR2_X1 U12991 ( .A1(n3258), .A2(n3135), .ZN(\mult_19/ab[7][16] ) );
  NOR2_X1 U12992 ( .A1(n3255), .A2(n3135), .ZN(\mult_19/ab[7][15] ) );
  NOR2_X1 U12993 ( .A1(n3252), .A2(n3135), .ZN(\mult_19/ab[7][14] ) );
  NOR2_X1 U12994 ( .A1(n3249), .A2(n3135), .ZN(\mult_19/ab[7][13] ) );
  NOR2_X1 U12995 ( .A1(n3246), .A2(n3135), .ZN(\mult_19/ab[7][12] ) );
  NOR2_X1 U12996 ( .A1(n3243), .A2(n3135), .ZN(\mult_19/ab[7][11] ) );
  NOR2_X1 U12997 ( .A1(n3240), .A2(n3135), .ZN(\mult_19/ab[7][10] ) );
  NOR2_X1 U12998 ( .A1(n3483), .A2(n3325), .ZN(\mult_20/ab[8][29] ) );
  NOR2_X1 U12999 ( .A1(n3480), .A2(n3325), .ZN(\mult_20/ab[8][28] ) );
  NOR2_X1 U13000 ( .A1(n3477), .A2(n3325), .ZN(\mult_20/ab[8][27] ) );
  NOR2_X1 U13001 ( .A1(n3474), .A2(n3325), .ZN(\mult_20/ab[8][26] ) );
  NOR2_X1 U13002 ( .A1(n3471), .A2(n3325), .ZN(\mult_20/ab[8][25] ) );
  NOR2_X1 U13003 ( .A1(n3468), .A2(n3325), .ZN(\mult_20/ab[8][24] ) );
  NOR2_X1 U13004 ( .A1(n3465), .A2(n3325), .ZN(\mult_20/ab[8][23] ) );
  NOR2_X1 U13005 ( .A1(n3462), .A2(n3325), .ZN(\mult_20/ab[8][22] ) );
  NOR2_X1 U13006 ( .A1(n3459), .A2(n3325), .ZN(\mult_20/ab[8][21] ) );
  NOR2_X1 U13007 ( .A1(n3456), .A2(n3325), .ZN(\mult_20/ab[8][20] ) );
  NOR2_X1 U13008 ( .A1(n3453), .A2(n3324), .ZN(\mult_20/ab[8][19] ) );
  NOR2_X1 U13009 ( .A1(n3450), .A2(n3324), .ZN(\mult_20/ab[8][18] ) );
  NOR2_X1 U13010 ( .A1(n3447), .A2(n3324), .ZN(\mult_20/ab[8][17] ) );
  NOR2_X1 U13011 ( .A1(n3441), .A2(n3324), .ZN(\mult_20/ab[8][15] ) );
  NOR2_X1 U13012 ( .A1(n3435), .A2(n3324), .ZN(\mult_20/ab[8][13] ) );
  NOR2_X1 U13013 ( .A1(n3429), .A2(n3324), .ZN(\mult_20/ab[8][11] ) );
  NOR2_X1 U13014 ( .A1(n3297), .A2(n3139), .ZN(\mult_19/ab[8][29] ) );
  NOR2_X1 U13015 ( .A1(n3294), .A2(n3139), .ZN(\mult_19/ab[8][28] ) );
  NOR2_X1 U13016 ( .A1(n3291), .A2(n3139), .ZN(\mult_19/ab[8][27] ) );
  NOR2_X1 U13017 ( .A1(n3288), .A2(n3139), .ZN(\mult_19/ab[8][26] ) );
  NOR2_X1 U13018 ( .A1(n3285), .A2(n3139), .ZN(\mult_19/ab[8][25] ) );
  NOR2_X1 U13019 ( .A1(n3282), .A2(n3139), .ZN(\mult_19/ab[8][24] ) );
  NOR2_X1 U13020 ( .A1(n3279), .A2(n3139), .ZN(\mult_19/ab[8][23] ) );
  NOR2_X1 U13021 ( .A1(n3276), .A2(n3139), .ZN(\mult_19/ab[8][22] ) );
  NOR2_X1 U13022 ( .A1(n3273), .A2(n3139), .ZN(\mult_19/ab[8][21] ) );
  NOR2_X1 U13023 ( .A1(n3270), .A2(n3139), .ZN(\mult_19/ab[8][20] ) );
  NOR2_X1 U13024 ( .A1(n3267), .A2(n3138), .ZN(\mult_19/ab[8][19] ) );
  NOR2_X1 U13025 ( .A1(n3264), .A2(n3138), .ZN(\mult_19/ab[8][18] ) );
  NOR2_X1 U13026 ( .A1(n3261), .A2(n3138), .ZN(\mult_19/ab[8][17] ) );
  NOR2_X1 U13027 ( .A1(n3483), .A2(n3328), .ZN(\mult_20/ab[9][29] ) );
  NOR2_X1 U13028 ( .A1(n3480), .A2(n3328), .ZN(\mult_20/ab[9][28] ) );
  NOR2_X1 U13029 ( .A1(n3477), .A2(n3328), .ZN(\mult_20/ab[9][27] ) );
  NOR2_X1 U13030 ( .A1(n3474), .A2(n3328), .ZN(\mult_20/ab[9][26] ) );
  NOR2_X1 U13031 ( .A1(n3471), .A2(n3328), .ZN(\mult_20/ab[9][25] ) );
  NOR2_X1 U13032 ( .A1(n3468), .A2(n3328), .ZN(\mult_20/ab[9][24] ) );
  NOR2_X1 U13033 ( .A1(n3465), .A2(n3328), .ZN(\mult_20/ab[9][23] ) );
  NOR2_X1 U13034 ( .A1(n3462), .A2(n3328), .ZN(\mult_20/ab[9][22] ) );
  NOR2_X1 U13035 ( .A1(n3459), .A2(n3328), .ZN(\mult_20/ab[9][21] ) );
  NOR2_X1 U13036 ( .A1(n3456), .A2(n3328), .ZN(\mult_20/ab[9][20] ) );
  NOR2_X1 U13037 ( .A1(n3453), .A2(n3327), .ZN(\mult_20/ab[9][19] ) );
  NOR2_X1 U13038 ( .A1(n3450), .A2(n3327), .ZN(\mult_20/ab[9][18] ) );
  NOR2_X1 U13039 ( .A1(n3447), .A2(n3327), .ZN(\mult_20/ab[9][17] ) );
  NOR2_X1 U13040 ( .A1(n3441), .A2(n3327), .ZN(\mult_20/ab[9][15] ) );
  NOR2_X1 U13041 ( .A1(n3435), .A2(n3327), .ZN(\mult_20/ab[9][13] ) );
  NOR2_X1 U13042 ( .A1(n3429), .A2(n3327), .ZN(\mult_20/ab[9][11] ) );
  NOR2_X1 U13043 ( .A1(n3297), .A2(n3142), .ZN(\mult_19/ab[9][29] ) );
  NOR2_X1 U13044 ( .A1(n3294), .A2(n3142), .ZN(\mult_19/ab[9][28] ) );
  NOR2_X1 U13045 ( .A1(n3291), .A2(n3142), .ZN(\mult_19/ab[9][27] ) );
  NOR2_X1 U13046 ( .A1(n3288), .A2(n3142), .ZN(\mult_19/ab[9][26] ) );
  NOR2_X1 U13047 ( .A1(n3285), .A2(n3142), .ZN(\mult_19/ab[9][25] ) );
  NOR2_X1 U13048 ( .A1(n3282), .A2(n3142), .ZN(\mult_19/ab[9][24] ) );
  NOR2_X1 U13049 ( .A1(n3279), .A2(n3142), .ZN(\mult_19/ab[9][23] ) );
  NOR2_X1 U13050 ( .A1(n3276), .A2(n3142), .ZN(\mult_19/ab[9][22] ) );
  NOR2_X1 U13051 ( .A1(n3273), .A2(n3142), .ZN(\mult_19/ab[9][21] ) );
  NOR2_X1 U13052 ( .A1(n3270), .A2(n3142), .ZN(\mult_19/ab[9][20] ) );
  NOR2_X1 U13053 ( .A1(n3267), .A2(n3141), .ZN(\mult_19/ab[9][19] ) );
  NOR2_X1 U13054 ( .A1(n3264), .A2(n3141), .ZN(\mult_19/ab[9][18] ) );
  NOR2_X1 U13055 ( .A1(n3255), .A2(n3141), .ZN(\mult_19/ab[9][15] ) );
  NOR2_X1 U13056 ( .A1(n3252), .A2(n3141), .ZN(\mult_19/ab[9][14] ) );
  NOR2_X1 U13057 ( .A1(n3249), .A2(n3141), .ZN(\mult_19/ab[9][13] ) );
  NOR2_X1 U13058 ( .A1(n3246), .A2(n3141), .ZN(\mult_19/ab[9][12] ) );
  NOR2_X1 U13059 ( .A1(n3243), .A2(n3141), .ZN(\mult_19/ab[9][11] ) );
  NOR2_X1 U13060 ( .A1(n3240), .A2(n3141), .ZN(\mult_19/ab[9][10] ) );
  NOR2_X1 U13061 ( .A1(n3483), .A2(n3331), .ZN(\mult_20/ab[10][29] ) );
  NOR2_X1 U13062 ( .A1(n3482), .A2(n3331), .ZN(\mult_20/ab[10][28] ) );
  NOR2_X1 U13063 ( .A1(n3479), .A2(n3331), .ZN(\mult_20/ab[10][27] ) );
  NOR2_X1 U13064 ( .A1(n3476), .A2(n3331), .ZN(\mult_20/ab[10][26] ) );
  NOR2_X1 U13065 ( .A1(n3473), .A2(n3331), .ZN(\mult_20/ab[10][25] ) );
  NOR2_X1 U13066 ( .A1(n3470), .A2(n3331), .ZN(\mult_20/ab[10][24] ) );
  NOR2_X1 U13067 ( .A1(n3467), .A2(n3331), .ZN(\mult_20/ab[10][23] ) );
  NOR2_X1 U13068 ( .A1(n3464), .A2(n3331), .ZN(\mult_20/ab[10][22] ) );
  NOR2_X1 U13069 ( .A1(n3461), .A2(n3331), .ZN(\mult_20/ab[10][21] ) );
  NOR2_X1 U13070 ( .A1(n3458), .A2(n3331), .ZN(\mult_20/ab[10][20] ) );
  NOR2_X1 U13071 ( .A1(n3455), .A2(n3330), .ZN(\mult_20/ab[10][19] ) );
  NOR2_X1 U13072 ( .A1(n3449), .A2(n3330), .ZN(\mult_20/ab[10][17] ) );
  NOR2_X1 U13073 ( .A1(n3443), .A2(n3330), .ZN(\mult_20/ab[10][15] ) );
  NOR2_X1 U13074 ( .A1(n3437), .A2(n3330), .ZN(\mult_20/ab[10][13] ) );
  NOR2_X1 U13075 ( .A1(n3431), .A2(n3330), .ZN(\mult_20/ab[10][11] ) );
  NOR2_X1 U13076 ( .A1(n3297), .A2(n3145), .ZN(\mult_19/ab[10][29] ) );
  NOR2_X1 U13077 ( .A1(n3296), .A2(n3145), .ZN(\mult_19/ab[10][28] ) );
  NOR2_X1 U13078 ( .A1(n3293), .A2(n3145), .ZN(\mult_19/ab[10][27] ) );
  NOR2_X1 U13079 ( .A1(n3290), .A2(n3145), .ZN(\mult_19/ab[10][26] ) );
  NOR2_X1 U13080 ( .A1(n3287), .A2(n3145), .ZN(\mult_19/ab[10][25] ) );
  NOR2_X1 U13081 ( .A1(n3284), .A2(n3145), .ZN(\mult_19/ab[10][24] ) );
  NOR2_X1 U13082 ( .A1(n3281), .A2(n3145), .ZN(\mult_19/ab[10][23] ) );
  NOR2_X1 U13083 ( .A1(n3278), .A2(n3145), .ZN(\mult_19/ab[10][22] ) );
  NOR2_X1 U13084 ( .A1(n3275), .A2(n3145), .ZN(\mult_19/ab[10][21] ) );
  NOR2_X1 U13085 ( .A1(n3272), .A2(n3145), .ZN(\mult_19/ab[10][20] ) );
  NOR2_X1 U13086 ( .A1(n3269), .A2(n3144), .ZN(\mult_19/ab[10][19] ) );
  NOR2_X1 U13087 ( .A1(n3266), .A2(n3144), .ZN(\mult_19/ab[10][18] ) );
  NOR2_X1 U13088 ( .A1(n3263), .A2(n3144), .ZN(\mult_19/ab[10][17] ) );
  NOR2_X1 U13089 ( .A1(n3260), .A2(n3144), .ZN(\mult_19/ab[10][16] ) );
  NOR2_X1 U13090 ( .A1(n3257), .A2(n3144), .ZN(\mult_19/ab[10][15] ) );
  NOR2_X1 U13091 ( .A1(n3485), .A2(n3334), .ZN(\mult_20/ab[11][29] ) );
  NOR2_X1 U13092 ( .A1(n3482), .A2(n3334), .ZN(\mult_20/ab[11][28] ) );
  NOR2_X1 U13093 ( .A1(n3479), .A2(n3334), .ZN(\mult_20/ab[11][27] ) );
  NOR2_X1 U13094 ( .A1(n3476), .A2(n3334), .ZN(\mult_20/ab[11][26] ) );
  NOR2_X1 U13095 ( .A1(n3473), .A2(n3334), .ZN(\mult_20/ab[11][25] ) );
  NOR2_X1 U13096 ( .A1(n3470), .A2(n3334), .ZN(\mult_20/ab[11][24] ) );
  NOR2_X1 U13097 ( .A1(n3467), .A2(n3334), .ZN(\mult_20/ab[11][23] ) );
  NOR2_X1 U13098 ( .A1(n3464), .A2(n3334), .ZN(\mult_20/ab[11][22] ) );
  NOR2_X1 U13099 ( .A1(n3461), .A2(n3334), .ZN(\mult_20/ab[11][21] ) );
  NOR2_X1 U13100 ( .A1(n3455), .A2(n3333), .ZN(\mult_20/ab[11][19] ) );
  NOR2_X1 U13101 ( .A1(n3449), .A2(n3333), .ZN(\mult_20/ab[11][17] ) );
  NOR2_X1 U13102 ( .A1(n3443), .A2(n3333), .ZN(\mult_20/ab[11][15] ) );
  NOR2_X1 U13103 ( .A1(n3437), .A2(n3333), .ZN(\mult_20/ab[11][13] ) );
  NOR2_X1 U13104 ( .A1(n3431), .A2(n3333), .ZN(\mult_20/ab[11][11] ) );
  NOR2_X1 U13105 ( .A1(n3299), .A2(n3148), .ZN(\mult_19/ab[11][29] ) );
  NOR2_X1 U13106 ( .A1(n3296), .A2(n3148), .ZN(\mult_19/ab[11][28] ) );
  NOR2_X1 U13107 ( .A1(n3293), .A2(n3148), .ZN(\mult_19/ab[11][27] ) );
  NOR2_X1 U13108 ( .A1(n3290), .A2(n3148), .ZN(\mult_19/ab[11][26] ) );
  NOR2_X1 U13109 ( .A1(n3287), .A2(n3148), .ZN(\mult_19/ab[11][25] ) );
  NOR2_X1 U13110 ( .A1(n3284), .A2(n3148), .ZN(\mult_19/ab[11][24] ) );
  NOR2_X1 U13111 ( .A1(n3281), .A2(n3148), .ZN(\mult_19/ab[11][23] ) );
  NOR2_X1 U13112 ( .A1(n3278), .A2(n3148), .ZN(\mult_19/ab[11][22] ) );
  NOR2_X1 U13113 ( .A1(n3272), .A2(n3148), .ZN(\mult_19/ab[11][20] ) );
  NOR2_X1 U13114 ( .A1(n3251), .A2(n3147), .ZN(\mult_19/ab[11][13] ) );
  NOR2_X1 U13115 ( .A1(n3248), .A2(n3147), .ZN(\mult_19/ab[11][12] ) );
  NOR2_X1 U13116 ( .A1(n3245), .A2(n3147), .ZN(\mult_19/ab[11][11] ) );
  NOR2_X1 U13117 ( .A1(n3242), .A2(n3147), .ZN(\mult_19/ab[11][10] ) );
  NOR2_X1 U13118 ( .A1(n3485), .A2(n3337), .ZN(\mult_20/ab[12][29] ) );
  NOR2_X1 U13119 ( .A1(n3482), .A2(n3337), .ZN(\mult_20/ab[12][28] ) );
  NOR2_X1 U13120 ( .A1(n3479), .A2(n3337), .ZN(\mult_20/ab[12][27] ) );
  NOR2_X1 U13121 ( .A1(n3476), .A2(n3337), .ZN(\mult_20/ab[12][26] ) );
  NOR2_X1 U13122 ( .A1(n3473), .A2(n3337), .ZN(\mult_20/ab[12][25] ) );
  NOR2_X1 U13123 ( .A1(n3470), .A2(n3337), .ZN(\mult_20/ab[12][24] ) );
  NOR2_X1 U13124 ( .A1(n3467), .A2(n3337), .ZN(\mult_20/ab[12][23] ) );
  NOR2_X1 U13125 ( .A1(n3464), .A2(n3337), .ZN(\mult_20/ab[12][22] ) );
  NOR2_X1 U13126 ( .A1(n3461), .A2(n3337), .ZN(\mult_20/ab[12][21] ) );
  NOR2_X1 U13127 ( .A1(n3458), .A2(n3337), .ZN(\mult_20/ab[12][20] ) );
  NOR2_X1 U13128 ( .A1(n3455), .A2(n3336), .ZN(\mult_20/ab[12][19] ) );
  NOR2_X1 U13129 ( .A1(n3449), .A2(n3336), .ZN(\mult_20/ab[12][17] ) );
  NOR2_X1 U13130 ( .A1(n3443), .A2(n3336), .ZN(\mult_20/ab[12][15] ) );
  NOR2_X1 U13131 ( .A1(n3437), .A2(n3336), .ZN(\mult_20/ab[12][13] ) );
  NOR2_X1 U13132 ( .A1(n3431), .A2(n3336), .ZN(\mult_20/ab[12][11] ) );
  NOR2_X1 U13133 ( .A1(n3299), .A2(n3151), .ZN(\mult_19/ab[12][29] ) );
  NOR2_X1 U13134 ( .A1(n3296), .A2(n3151), .ZN(\mult_19/ab[12][28] ) );
  NOR2_X1 U13135 ( .A1(n3293), .A2(n3151), .ZN(\mult_19/ab[12][27] ) );
  NOR2_X1 U13136 ( .A1(n3290), .A2(n3151), .ZN(\mult_19/ab[12][26] ) );
  NOR2_X1 U13137 ( .A1(n3287), .A2(n3151), .ZN(\mult_19/ab[12][25] ) );
  NOR2_X1 U13138 ( .A1(n3284), .A2(n3151), .ZN(\mult_19/ab[12][24] ) );
  NOR2_X1 U13139 ( .A1(n3281), .A2(n3151), .ZN(\mult_19/ab[12][23] ) );
  NOR2_X1 U13140 ( .A1(n3278), .A2(n3151), .ZN(\mult_19/ab[12][22] ) );
  NOR2_X1 U13141 ( .A1(n3275), .A2(n3151), .ZN(\mult_19/ab[12][21] ) );
  NOR2_X1 U13142 ( .A1(n3272), .A2(n3151), .ZN(\mult_19/ab[12][20] ) );
  NOR2_X1 U13143 ( .A1(n3266), .A2(n3150), .ZN(\mult_19/ab[12][18] ) );
  NOR2_X1 U13144 ( .A1(n3263), .A2(n3150), .ZN(\mult_19/ab[12][17] ) );
  NOR2_X1 U13145 ( .A1(n3260), .A2(n3150), .ZN(\mult_19/ab[12][16] ) );
  NOR2_X1 U13146 ( .A1(n3257), .A2(n3150), .ZN(\mult_19/ab[12][15] ) );
  NOR2_X1 U13147 ( .A1(n3254), .A2(n3150), .ZN(\mult_19/ab[12][14] ) );
  NOR2_X1 U13148 ( .A1(n3251), .A2(n3150), .ZN(\mult_19/ab[12][13] ) );
  NOR2_X1 U13149 ( .A1(n3482), .A2(n3340), .ZN(\mult_20/ab[13][28] ) );
  NOR2_X1 U13150 ( .A1(n3479), .A2(n3340), .ZN(\mult_20/ab[13][27] ) );
  NOR2_X1 U13151 ( .A1(n3476), .A2(n3340), .ZN(\mult_20/ab[13][26] ) );
  NOR2_X1 U13152 ( .A1(n3473), .A2(n3340), .ZN(\mult_20/ab[13][25] ) );
  NOR2_X1 U13153 ( .A1(n3470), .A2(n3340), .ZN(\mult_20/ab[13][24] ) );
  NOR2_X1 U13154 ( .A1(n3467), .A2(n3340), .ZN(\mult_20/ab[13][23] ) );
  NOR2_X1 U13155 ( .A1(n3464), .A2(n3340), .ZN(\mult_20/ab[13][22] ) );
  NOR2_X1 U13156 ( .A1(n3461), .A2(n3340), .ZN(\mult_20/ab[13][21] ) );
  NOR2_X1 U13157 ( .A1(n3458), .A2(n3340), .ZN(\mult_20/ab[13][20] ) );
  NOR2_X1 U13158 ( .A1(n3455), .A2(n3339), .ZN(\mult_20/ab[13][19] ) );
  NOR2_X1 U13159 ( .A1(n3449), .A2(n3339), .ZN(\mult_20/ab[13][17] ) );
  NOR2_X1 U13160 ( .A1(n3446), .A2(n3339), .ZN(\mult_20/ab[13][16] ) );
  NOR2_X1 U13161 ( .A1(n3443), .A2(n3339), .ZN(\mult_20/ab[13][15] ) );
  NOR2_X1 U13162 ( .A1(n3440), .A2(n3339), .ZN(\mult_20/ab[13][14] ) );
  NOR2_X1 U13163 ( .A1(n3437), .A2(n3339), .ZN(\mult_20/ab[13][13] ) );
  NOR2_X1 U13164 ( .A1(n3431), .A2(n3339), .ZN(\mult_20/ab[13][11] ) );
  NOR2_X1 U13165 ( .A1(n3296), .A2(n3154), .ZN(\mult_19/ab[13][28] ) );
  NOR2_X1 U13166 ( .A1(n3293), .A2(n3154), .ZN(\mult_19/ab[13][27] ) );
  NOR2_X1 U13167 ( .A1(n3290), .A2(n3154), .ZN(\mult_19/ab[13][26] ) );
  NOR2_X1 U13168 ( .A1(n3287), .A2(n3154), .ZN(\mult_19/ab[13][25] ) );
  NOR2_X1 U13169 ( .A1(n3284), .A2(n3154), .ZN(\mult_19/ab[13][24] ) );
  NOR2_X1 U13170 ( .A1(n3281), .A2(n3154), .ZN(\mult_19/ab[13][23] ) );
  NOR2_X1 U13171 ( .A1(n3278), .A2(n3154), .ZN(\mult_19/ab[13][22] ) );
  NOR2_X1 U13172 ( .A1(n3275), .A2(n3154), .ZN(\mult_19/ab[13][21] ) );
  NOR2_X1 U13173 ( .A1(n3272), .A2(n3154), .ZN(\mult_19/ab[13][20] ) );
  NOR2_X1 U13174 ( .A1(n3269), .A2(n3153), .ZN(\mult_19/ab[13][19] ) );
  NOR2_X1 U13175 ( .A1(n3266), .A2(n3153), .ZN(\mult_19/ab[13][18] ) );
  NOR2_X1 U13176 ( .A1(n3263), .A2(n3153), .ZN(\mult_19/ab[13][17] ) );
  NOR2_X1 U13177 ( .A1(n3260), .A2(n3153), .ZN(\mult_19/ab[13][16] ) );
  NOR2_X1 U13178 ( .A1(n3257), .A2(n3153), .ZN(\mult_19/ab[13][15] ) );
  NOR2_X1 U13179 ( .A1(n3245), .A2(n3153), .ZN(\mult_19/ab[13][11] ) );
  NOR2_X1 U13180 ( .A1(n3242), .A2(n3153), .ZN(\mult_19/ab[13][10] ) );
  NOR2_X1 U13181 ( .A1(n3479), .A2(n3343), .ZN(\mult_20/ab[14][27] ) );
  NOR2_X1 U13182 ( .A1(n3476), .A2(n3343), .ZN(\mult_20/ab[14][26] ) );
  NOR2_X1 U13183 ( .A1(n3473), .A2(n3343), .ZN(\mult_20/ab[14][25] ) );
  NOR2_X1 U13184 ( .A1(n3470), .A2(n3343), .ZN(\mult_20/ab[14][24] ) );
  NOR2_X1 U13185 ( .A1(n3467), .A2(n3343), .ZN(\mult_20/ab[14][23] ) );
  NOR2_X1 U13186 ( .A1(n3464), .A2(n3343), .ZN(\mult_20/ab[14][22] ) );
  NOR2_X1 U13187 ( .A1(n3461), .A2(n3343), .ZN(\mult_20/ab[14][21] ) );
  NOR2_X1 U13188 ( .A1(n3458), .A2(n3343), .ZN(\mult_20/ab[14][20] ) );
  NOR2_X1 U13189 ( .A1(n3455), .A2(n3342), .ZN(\mult_20/ab[14][19] ) );
  NOR2_X1 U13190 ( .A1(n3452), .A2(n3342), .ZN(\mult_20/ab[14][18] ) );
  NOR2_X1 U13191 ( .A1(n3449), .A2(n3342), .ZN(\mult_20/ab[14][17] ) );
  NOR2_X1 U13192 ( .A1(n3443), .A2(n3342), .ZN(\mult_20/ab[14][15] ) );
  NOR2_X1 U13193 ( .A1(n3437), .A2(n3342), .ZN(\mult_20/ab[14][13] ) );
  NOR2_X1 U13194 ( .A1(n3431), .A2(n3342), .ZN(\mult_20/ab[14][11] ) );
  NOR2_X1 U13195 ( .A1(n3293), .A2(n3157), .ZN(\mult_19/ab[14][27] ) );
  NOR2_X1 U13196 ( .A1(n3290), .A2(n3157), .ZN(\mult_19/ab[14][26] ) );
  NOR2_X1 U13197 ( .A1(n3287), .A2(n3157), .ZN(\mult_19/ab[14][25] ) );
  NOR2_X1 U13198 ( .A1(n3284), .A2(n3157), .ZN(\mult_19/ab[14][24] ) );
  NOR2_X1 U13199 ( .A1(n3281), .A2(n3157), .ZN(\mult_19/ab[14][23] ) );
  NOR2_X1 U13200 ( .A1(n3278), .A2(n3157), .ZN(\mult_19/ab[14][22] ) );
  NOR2_X1 U13201 ( .A1(n3275), .A2(n3157), .ZN(\mult_19/ab[14][21] ) );
  NOR2_X1 U13202 ( .A1(n3272), .A2(n3157), .ZN(\mult_19/ab[14][20] ) );
  NOR2_X1 U13203 ( .A1(n3269), .A2(n3156), .ZN(\mult_19/ab[14][19] ) );
  NOR2_X1 U13204 ( .A1(n3266), .A2(n3156), .ZN(\mult_19/ab[14][18] ) );
  NOR2_X1 U13205 ( .A1(n3260), .A2(n3156), .ZN(\mult_19/ab[14][16] ) );
  NOR2_X1 U13206 ( .A1(n3257), .A2(n3156), .ZN(\mult_19/ab[14][15] ) );
  NOR2_X1 U13207 ( .A1(n3254), .A2(n3156), .ZN(\mult_19/ab[14][14] ) );
  NOR2_X1 U13208 ( .A1(n3251), .A2(n3156), .ZN(\mult_19/ab[14][13] ) );
  NOR2_X1 U13209 ( .A1(n3248), .A2(n3156), .ZN(\mult_19/ab[14][12] ) );
  NOR2_X1 U13210 ( .A1(n3245), .A2(n3156), .ZN(\mult_19/ab[14][11] ) );
  NOR2_X1 U13211 ( .A1(n3476), .A2(n3346), .ZN(\mult_20/ab[15][26] ) );
  NOR2_X1 U13212 ( .A1(n3473), .A2(n3346), .ZN(\mult_20/ab[15][25] ) );
  NOR2_X1 U13213 ( .A1(n3470), .A2(n3346), .ZN(\mult_20/ab[15][24] ) );
  NOR2_X1 U13214 ( .A1(n3467), .A2(n3346), .ZN(\mult_20/ab[15][23] ) );
  NOR2_X1 U13215 ( .A1(n3464), .A2(n3346), .ZN(\mult_20/ab[15][22] ) );
  NOR2_X1 U13216 ( .A1(n3461), .A2(n3346), .ZN(\mult_20/ab[15][21] ) );
  NOR2_X1 U13217 ( .A1(n3458), .A2(n3346), .ZN(\mult_20/ab[15][20] ) );
  NOR2_X1 U13218 ( .A1(n3455), .A2(n3345), .ZN(\mult_20/ab[15][19] ) );
  NOR2_X1 U13219 ( .A1(n3452), .A2(n3345), .ZN(\mult_20/ab[15][18] ) );
  NOR2_X1 U13220 ( .A1(n3449), .A2(n3345), .ZN(\mult_20/ab[15][17] ) );
  NOR2_X1 U13221 ( .A1(n3443), .A2(n3345), .ZN(\mult_20/ab[15][15] ) );
  NOR2_X1 U13222 ( .A1(n3437), .A2(n3345), .ZN(\mult_20/ab[15][13] ) );
  NOR2_X1 U13223 ( .A1(n3431), .A2(n3345), .ZN(\mult_20/ab[15][11] ) );
  NOR2_X1 U13224 ( .A1(n3290), .A2(n3160), .ZN(\mult_19/ab[15][26] ) );
  NOR2_X1 U13225 ( .A1(n3287), .A2(n3160), .ZN(\mult_19/ab[15][25] ) );
  NOR2_X1 U13226 ( .A1(n3284), .A2(n3160), .ZN(\mult_19/ab[15][24] ) );
  NOR2_X1 U13227 ( .A1(n3281), .A2(n3160), .ZN(\mult_19/ab[15][23] ) );
  NOR2_X1 U13228 ( .A1(n3278), .A2(n3160), .ZN(\mult_19/ab[15][22] ) );
  NOR2_X1 U13229 ( .A1(n3275), .A2(n3160), .ZN(\mult_19/ab[15][21] ) );
  NOR2_X1 U13230 ( .A1(n3272), .A2(n3160), .ZN(\mult_19/ab[15][20] ) );
  NOR2_X1 U13231 ( .A1(n3269), .A2(n3159), .ZN(\mult_19/ab[15][19] ) );
  NOR2_X1 U13232 ( .A1(n3266), .A2(n3159), .ZN(\mult_19/ab[15][18] ) );
  NOR2_X1 U13233 ( .A1(n3260), .A2(n3159), .ZN(\mult_19/ab[15][16] ) );
  NOR2_X1 U13234 ( .A1(n3473), .A2(n3349), .ZN(\mult_20/ab[16][25] ) );
  NOR2_X1 U13235 ( .A1(n3470), .A2(n3349), .ZN(\mult_20/ab[16][24] ) );
  NOR2_X1 U13236 ( .A1(n3466), .A2(n3349), .ZN(\mult_20/ab[16][23] ) );
  NOR2_X1 U13237 ( .A1(n3464), .A2(n3349), .ZN(\mult_20/ab[16][22] ) );
  NOR2_X1 U13238 ( .A1(n3461), .A2(n3349), .ZN(\mult_20/ab[16][21] ) );
  NOR2_X1 U13239 ( .A1(n3458), .A2(n3349), .ZN(\mult_20/ab[16][20] ) );
  NOR2_X1 U13240 ( .A1(n3455), .A2(n3348), .ZN(\mult_20/ab[16][19] ) );
  NOR2_X1 U13241 ( .A1(n3452), .A2(n3348), .ZN(\mult_20/ab[16][18] ) );
  NOR2_X1 U13242 ( .A1(n3449), .A2(n3348), .ZN(\mult_20/ab[16][17] ) );
  NOR2_X1 U13243 ( .A1(n3446), .A2(n3348), .ZN(\mult_20/ab[16][16] ) );
  NOR2_X1 U13244 ( .A1(n3443), .A2(n3348), .ZN(\mult_20/ab[16][15] ) );
  NOR2_X1 U13245 ( .A1(n3437), .A2(n3348), .ZN(\mult_20/ab[16][13] ) );
  NOR2_X1 U13246 ( .A1(n3431), .A2(n3348), .ZN(\mult_20/ab[16][11] ) );
  NOR2_X1 U13247 ( .A1(n3287), .A2(n3163), .ZN(\mult_19/ab[16][25] ) );
  NOR2_X1 U13248 ( .A1(n3284), .A2(n3163), .ZN(\mult_19/ab[16][24] ) );
  NOR2_X1 U13249 ( .A1(n3280), .A2(n3163), .ZN(\mult_19/ab[16][23] ) );
  NOR2_X1 U13250 ( .A1(n3278), .A2(n3163), .ZN(\mult_19/ab[16][22] ) );
  NOR2_X1 U13251 ( .A1(n3275), .A2(n3163), .ZN(\mult_19/ab[16][21] ) );
  NOR2_X1 U13252 ( .A1(n3272), .A2(n3163), .ZN(\mult_19/ab[16][20] ) );
  NOR2_X1 U13253 ( .A1(n3269), .A2(n3162), .ZN(\mult_19/ab[16][19] ) );
  NOR2_X1 U13254 ( .A1(n3266), .A2(n3162), .ZN(\mult_19/ab[16][18] ) );
  NOR2_X1 U13255 ( .A1(n3263), .A2(n3162), .ZN(\mult_19/ab[16][17] ) );
  NOR2_X1 U13256 ( .A1(n3260), .A2(n3162), .ZN(\mult_19/ab[16][16] ) );
  NOR2_X1 U13257 ( .A1(n3254), .A2(n3162), .ZN(\mult_19/ab[16][14] ) );
  NOR2_X1 U13258 ( .A1(n3251), .A2(n3162), .ZN(\mult_19/ab[16][13] ) );
  NOR2_X1 U13259 ( .A1(n3248), .A2(n3162), .ZN(\mult_19/ab[16][12] ) );
  NOR2_X1 U13260 ( .A1(n3245), .A2(n3162), .ZN(\mult_19/ab[16][11] ) );
  NOR2_X1 U13261 ( .A1(n3242), .A2(n3162), .ZN(\mult_19/ab[16][10] ) );
  NOR2_X1 U13262 ( .A1(n3469), .A2(n3352), .ZN(\mult_20/ab[17][24] ) );
  NOR2_X1 U13263 ( .A1(n3466), .A2(n3352), .ZN(\mult_20/ab[17][23] ) );
  NOR2_X1 U13264 ( .A1(n3463), .A2(n3352), .ZN(\mult_20/ab[17][22] ) );
  NOR2_X1 U13265 ( .A1(n3460), .A2(n3352), .ZN(\mult_20/ab[17][21] ) );
  NOR2_X1 U13266 ( .A1(n3457), .A2(n3352), .ZN(\mult_20/ab[17][20] ) );
  NOR2_X1 U13267 ( .A1(n3454), .A2(n3351), .ZN(\mult_20/ab[17][19] ) );
  NOR2_X1 U13268 ( .A1(n3451), .A2(n3351), .ZN(\mult_20/ab[17][18] ) );
  NOR2_X1 U13269 ( .A1(n3448), .A2(n3351), .ZN(\mult_20/ab[17][17] ) );
  NOR2_X1 U13270 ( .A1(n3445), .A2(n3351), .ZN(\mult_20/ab[17][16] ) );
  NOR2_X1 U13271 ( .A1(n3442), .A2(n3351), .ZN(\mult_20/ab[17][15] ) );
  NOR2_X1 U13272 ( .A1(n3436), .A2(n3351), .ZN(\mult_20/ab[17][13] ) );
  NOR2_X1 U13273 ( .A1(n3430), .A2(n3351), .ZN(\mult_20/ab[17][11] ) );
  NOR2_X1 U13274 ( .A1(n3485), .A2(n3340), .ZN(\mult_20/ab[13][29] ) );
  NOR2_X1 U13275 ( .A1(n3283), .A2(n3166), .ZN(\mult_19/ab[17][24] ) );
  NOR2_X1 U13276 ( .A1(n3280), .A2(n3166), .ZN(\mult_19/ab[17][23] ) );
  NOR2_X1 U13277 ( .A1(n3277), .A2(n3166), .ZN(\mult_19/ab[17][22] ) );
  NOR2_X1 U13278 ( .A1(n3274), .A2(n3166), .ZN(\mult_19/ab[17][21] ) );
  NOR2_X1 U13279 ( .A1(n3271), .A2(n3166), .ZN(\mult_19/ab[17][20] ) );
  NOR2_X1 U13280 ( .A1(n3268), .A2(n3165), .ZN(\mult_19/ab[17][19] ) );
  NOR2_X1 U13281 ( .A1(n3265), .A2(n3165), .ZN(\mult_19/ab[17][18] ) );
  NOR2_X1 U13282 ( .A1(n3262), .A2(n3165), .ZN(\mult_19/ab[17][17] ) );
  NOR2_X1 U13283 ( .A1(n3259), .A2(n3165), .ZN(\mult_19/ab[17][16] ) );
  NOR2_X1 U13284 ( .A1(n3253), .A2(n3165), .ZN(\mult_19/ab[17][14] ) );
  NOR2_X1 U13285 ( .A1(n3299), .A2(n3154), .ZN(\mult_19/ab[13][29] ) );
  NOR2_X1 U13286 ( .A1(n3466), .A2(n3355), .ZN(\mult_20/ab[18][23] ) );
  NOR2_X1 U13287 ( .A1(n3463), .A2(n3355), .ZN(\mult_20/ab[18][22] ) );
  NOR2_X1 U13288 ( .A1(n3460), .A2(n3355), .ZN(\mult_20/ab[18][21] ) );
  NOR2_X1 U13289 ( .A1(n3457), .A2(n3355), .ZN(\mult_20/ab[18][20] ) );
  NOR2_X1 U13290 ( .A1(n3454), .A2(n3354), .ZN(\mult_20/ab[18][19] ) );
  NOR2_X1 U13291 ( .A1(n3451), .A2(n3354), .ZN(\mult_20/ab[18][18] ) );
  NOR2_X1 U13292 ( .A1(n3448), .A2(n3354), .ZN(\mult_20/ab[18][17] ) );
  NOR2_X1 U13293 ( .A1(n3445), .A2(n3354), .ZN(\mult_20/ab[18][16] ) );
  NOR2_X1 U13294 ( .A1(n3442), .A2(n3354), .ZN(\mult_20/ab[18][15] ) );
  NOR2_X1 U13295 ( .A1(n3439), .A2(n3354), .ZN(\mult_20/ab[18][14] ) );
  NOR2_X1 U13296 ( .A1(n3436), .A2(n3354), .ZN(\mult_20/ab[18][13] ) );
  NOR2_X1 U13297 ( .A1(n3430), .A2(n3354), .ZN(\mult_20/ab[18][11] ) );
  NOR2_X1 U13298 ( .A1(n3485), .A2(n3343), .ZN(\mult_20/ab[14][29] ) );
  NOR2_X1 U13299 ( .A1(n3482), .A2(n3343), .ZN(\mult_20/ab[14][28] ) );
  NOR2_X1 U13300 ( .A1(n3280), .A2(n3169), .ZN(\mult_19/ab[18][23] ) );
  NOR2_X1 U13301 ( .A1(n3277), .A2(n3169), .ZN(\mult_19/ab[18][22] ) );
  NOR2_X1 U13302 ( .A1(n3274), .A2(n3169), .ZN(\mult_19/ab[18][21] ) );
  NOR2_X1 U13303 ( .A1(n3271), .A2(n3169), .ZN(\mult_19/ab[18][20] ) );
  NOR2_X1 U13304 ( .A1(n3268), .A2(n3168), .ZN(\mult_19/ab[18][19] ) );
  NOR2_X1 U13305 ( .A1(n3265), .A2(n3168), .ZN(\mult_19/ab[18][18] ) );
  NOR2_X1 U13306 ( .A1(n3262), .A2(n3168), .ZN(\mult_19/ab[18][17] ) );
  NOR2_X1 U13307 ( .A1(n3259), .A2(n3168), .ZN(\mult_19/ab[18][16] ) );
  NOR2_X1 U13308 ( .A1(n3256), .A2(n3168), .ZN(\mult_19/ab[18][15] ) );
  NOR2_X1 U13309 ( .A1(n3253), .A2(n3168), .ZN(\mult_19/ab[18][14] ) );
  NOR2_X1 U13310 ( .A1(n3247), .A2(n3168), .ZN(\mult_19/ab[18][12] ) );
  NOR2_X1 U13311 ( .A1(n3244), .A2(n3168), .ZN(\mult_19/ab[18][11] ) );
  NOR2_X1 U13312 ( .A1(n3241), .A2(n3168), .ZN(\mult_19/ab[18][10] ) );
  NOR2_X1 U13313 ( .A1(n3299), .A2(n3157), .ZN(\mult_19/ab[14][29] ) );
  NOR2_X1 U13314 ( .A1(n3296), .A2(n3157), .ZN(\mult_19/ab[14][28] ) );
  NOR2_X1 U13315 ( .A1(n3463), .A2(n3358), .ZN(\mult_20/ab[19][22] ) );
  NOR2_X1 U13316 ( .A1(n3460), .A2(n3358), .ZN(\mult_20/ab[19][21] ) );
  NOR2_X1 U13317 ( .A1(n3457), .A2(n3358), .ZN(\mult_20/ab[19][20] ) );
  NOR2_X1 U13318 ( .A1(n3454), .A2(n3357), .ZN(\mult_20/ab[19][19] ) );
  NOR2_X1 U13319 ( .A1(n3451), .A2(n3357), .ZN(\mult_20/ab[19][18] ) );
  NOR2_X1 U13320 ( .A1(n3448), .A2(n3357), .ZN(\mult_20/ab[19][17] ) );
  NOR2_X1 U13321 ( .A1(n3445), .A2(n3357), .ZN(\mult_20/ab[19][16] ) );
  NOR2_X1 U13322 ( .A1(n3442), .A2(n3357), .ZN(\mult_20/ab[19][15] ) );
  NOR2_X1 U13323 ( .A1(n3439), .A2(n3357), .ZN(\mult_20/ab[19][14] ) );
  NOR2_X1 U13324 ( .A1(n3436), .A2(n3357), .ZN(\mult_20/ab[19][13] ) );
  NOR2_X1 U13325 ( .A1(n3430), .A2(n3357), .ZN(\mult_20/ab[19][11] ) );
  NOR2_X1 U13326 ( .A1(n3485), .A2(n3346), .ZN(\mult_20/ab[15][29] ) );
  NOR2_X1 U13327 ( .A1(n3482), .A2(n3346), .ZN(\mult_20/ab[15][28] ) );
  NOR2_X1 U13328 ( .A1(n3479), .A2(n3346), .ZN(\mult_20/ab[15][27] ) );
  NOR2_X1 U13329 ( .A1(n3277), .A2(n3172), .ZN(\mult_19/ab[19][22] ) );
  NOR2_X1 U13330 ( .A1(n3274), .A2(n3172), .ZN(\mult_19/ab[19][21] ) );
  NOR2_X1 U13331 ( .A1(n3271), .A2(n3172), .ZN(\mult_19/ab[19][20] ) );
  NOR2_X1 U13332 ( .A1(n3268), .A2(n3171), .ZN(\mult_19/ab[19][19] ) );
  NOR2_X1 U13333 ( .A1(n3265), .A2(n3171), .ZN(\mult_19/ab[19][18] ) );
  NOR2_X1 U13334 ( .A1(n3262), .A2(n3171), .ZN(\mult_19/ab[19][17] ) );
  NOR2_X1 U13335 ( .A1(n3259), .A2(n3171), .ZN(\mult_19/ab[19][16] ) );
  NOR2_X1 U13336 ( .A1(n3256), .A2(n3171), .ZN(\mult_19/ab[19][15] ) );
  NOR2_X1 U13337 ( .A1(n3253), .A2(n3171), .ZN(\mult_19/ab[19][14] ) );
  NOR2_X1 U13338 ( .A1(n3247), .A2(n3171), .ZN(\mult_19/ab[19][12] ) );
  NOR2_X1 U13339 ( .A1(n3299), .A2(n3160), .ZN(\mult_19/ab[15][29] ) );
  NOR2_X1 U13340 ( .A1(n3296), .A2(n3160), .ZN(\mult_19/ab[15][28] ) );
  NOR2_X1 U13341 ( .A1(n3293), .A2(n3160), .ZN(\mult_19/ab[15][27] ) );
  NOR2_X1 U13342 ( .A1(n3460), .A2(n3361), .ZN(\mult_20/ab[20][21] ) );
  NOR2_X1 U13343 ( .A1(n3457), .A2(n3361), .ZN(\mult_20/ab[20][20] ) );
  NOR2_X1 U13344 ( .A1(n3454), .A2(n3360), .ZN(\mult_20/ab[20][19] ) );
  NOR2_X1 U13345 ( .A1(n3451), .A2(n3360), .ZN(\mult_20/ab[20][18] ) );
  NOR2_X1 U13346 ( .A1(n3448), .A2(n3360), .ZN(\mult_20/ab[20][17] ) );
  NOR2_X1 U13347 ( .A1(n3445), .A2(n3360), .ZN(\mult_20/ab[20][16] ) );
  NOR2_X1 U13348 ( .A1(n3442), .A2(n3360), .ZN(\mult_20/ab[20][15] ) );
  NOR2_X1 U13349 ( .A1(n3439), .A2(n3360), .ZN(\mult_20/ab[20][14] ) );
  NOR2_X1 U13350 ( .A1(n3436), .A2(n3360), .ZN(\mult_20/ab[20][13] ) );
  NOR2_X1 U13351 ( .A1(n3433), .A2(n3360), .ZN(\mult_20/ab[20][12] ) );
  NOR2_X1 U13352 ( .A1(n3430), .A2(n3360), .ZN(\mult_20/ab[20][11] ) );
  NOR2_X1 U13353 ( .A1(n3482), .A2(n3349), .ZN(\mult_20/ab[16][28] ) );
  NOR2_X1 U13354 ( .A1(n3479), .A2(n3349), .ZN(\mult_20/ab[16][27] ) );
  NOR2_X1 U13355 ( .A1(n3476), .A2(n3349), .ZN(\mult_20/ab[16][26] ) );
  NOR2_X1 U13356 ( .A1(n3274), .A2(n3175), .ZN(\mult_19/ab[20][21] ) );
  NOR2_X1 U13357 ( .A1(n3271), .A2(n3175), .ZN(\mult_19/ab[20][20] ) );
  NOR2_X1 U13358 ( .A1(n3268), .A2(n3174), .ZN(\mult_19/ab[20][19] ) );
  NOR2_X1 U13359 ( .A1(n3265), .A2(n3174), .ZN(\mult_19/ab[20][18] ) );
  NOR2_X1 U13360 ( .A1(n3262), .A2(n3174), .ZN(\mult_19/ab[20][17] ) );
  NOR2_X1 U13361 ( .A1(n3259), .A2(n3174), .ZN(\mult_19/ab[20][16] ) );
  NOR2_X1 U13362 ( .A1(n3256), .A2(n3174), .ZN(\mult_19/ab[20][15] ) );
  NOR2_X1 U13363 ( .A1(n3253), .A2(n3174), .ZN(\mult_19/ab[20][14] ) );
  NOR2_X1 U13364 ( .A1(n3250), .A2(n3174), .ZN(\mult_19/ab[20][13] ) );
  NOR2_X1 U13365 ( .A1(n3247), .A2(n3174), .ZN(\mult_19/ab[20][12] ) );
  NOR2_X1 U13366 ( .A1(n3241), .A2(n3174), .ZN(\mult_19/ab[20][10] ) );
  NOR2_X1 U13367 ( .A1(n3296), .A2(n3163), .ZN(\mult_19/ab[16][28] ) );
  NOR2_X1 U13368 ( .A1(n3293), .A2(n3163), .ZN(\mult_19/ab[16][27] ) );
  NOR2_X1 U13369 ( .A1(n3290), .A2(n3163), .ZN(\mult_19/ab[16][26] ) );
  NOR2_X1 U13370 ( .A1(n3457), .A2(n3364), .ZN(\mult_20/ab[21][20] ) );
  NOR2_X1 U13371 ( .A1(n3454), .A2(n3363), .ZN(\mult_20/ab[21][19] ) );
  NOR2_X1 U13372 ( .A1(n3451), .A2(n3363), .ZN(\mult_20/ab[21][18] ) );
  NOR2_X1 U13373 ( .A1(n3448), .A2(n3363), .ZN(\mult_20/ab[21][17] ) );
  NOR2_X1 U13374 ( .A1(n3445), .A2(n3363), .ZN(\mult_20/ab[21][16] ) );
  NOR2_X1 U13375 ( .A1(n3442), .A2(n3363), .ZN(\mult_20/ab[21][15] ) );
  NOR2_X1 U13376 ( .A1(n3439), .A2(n3363), .ZN(\mult_20/ab[21][14] ) );
  NOR2_X1 U13377 ( .A1(n3436), .A2(n3363), .ZN(\mult_20/ab[21][13] ) );
  NOR2_X1 U13378 ( .A1(n3433), .A2(n3363), .ZN(\mult_20/ab[21][12] ) );
  NOR2_X1 U13379 ( .A1(n3430), .A2(n3363), .ZN(\mult_20/ab[21][11] ) );
  NOR2_X1 U13380 ( .A1(n3478), .A2(n3352), .ZN(\mult_20/ab[17][27] ) );
  NOR2_X1 U13381 ( .A1(n3475), .A2(n3352), .ZN(\mult_20/ab[17][26] ) );
  NOR2_X1 U13382 ( .A1(n3472), .A2(n3352), .ZN(\mult_20/ab[17][25] ) );
  NOR2_X1 U13383 ( .A1(n3271), .A2(n3178), .ZN(\mult_19/ab[21][20] ) );
  NOR2_X1 U13384 ( .A1(n3268), .A2(n3177), .ZN(\mult_19/ab[21][19] ) );
  NOR2_X1 U13385 ( .A1(n3265), .A2(n3177), .ZN(\mult_19/ab[21][18] ) );
  NOR2_X1 U13386 ( .A1(n3262), .A2(n3177), .ZN(\mult_19/ab[21][17] ) );
  NOR2_X1 U13387 ( .A1(n3259), .A2(n3177), .ZN(\mult_19/ab[21][16] ) );
  NOR2_X1 U13388 ( .A1(n3256), .A2(n3177), .ZN(\mult_19/ab[21][15] ) );
  NOR2_X1 U13389 ( .A1(n3253), .A2(n3177), .ZN(\mult_19/ab[21][14] ) );
  NOR2_X1 U13390 ( .A1(n3250), .A2(n3177), .ZN(\mult_19/ab[21][13] ) );
  NOR2_X1 U13391 ( .A1(n3247), .A2(n3177), .ZN(\mult_19/ab[21][12] ) );
  NOR2_X1 U13392 ( .A1(n3241), .A2(n3177), .ZN(\mult_19/ab[21][10] ) );
  NOR2_X1 U13393 ( .A1(n3292), .A2(n3166), .ZN(\mult_19/ab[17][27] ) );
  NOR2_X1 U13394 ( .A1(n3289), .A2(n3166), .ZN(\mult_19/ab[17][26] ) );
  NOR2_X1 U13395 ( .A1(n3286), .A2(n3166), .ZN(\mult_19/ab[17][25] ) );
  NOR2_X1 U13396 ( .A1(n3454), .A2(n3366), .ZN(\mult_20/ab[22][19] ) );
  NOR2_X1 U13397 ( .A1(n3451), .A2(n3366), .ZN(\mult_20/ab[22][18] ) );
  NOR2_X1 U13398 ( .A1(n3448), .A2(n3366), .ZN(\mult_20/ab[22][17] ) );
  NOR2_X1 U13399 ( .A1(n3445), .A2(n3366), .ZN(\mult_20/ab[22][16] ) );
  NOR2_X1 U13400 ( .A1(n3442), .A2(n3366), .ZN(\mult_20/ab[22][15] ) );
  NOR2_X1 U13401 ( .A1(n3439), .A2(n3366), .ZN(\mult_20/ab[22][14] ) );
  NOR2_X1 U13402 ( .A1(n3436), .A2(n3366), .ZN(\mult_20/ab[22][13] ) );
  NOR2_X1 U13403 ( .A1(n3433), .A2(n3366), .ZN(\mult_20/ab[22][12] ) );
  NOR2_X1 U13404 ( .A1(n3430), .A2(n3366), .ZN(\mult_20/ab[22][11] ) );
  NOR2_X1 U13405 ( .A1(n3427), .A2(n3366), .ZN(\mult_20/ab[22][10] ) );
  NOR2_X1 U13406 ( .A1(n3475), .A2(n3355), .ZN(\mult_20/ab[18][26] ) );
  NOR2_X1 U13407 ( .A1(n3472), .A2(n3355), .ZN(\mult_20/ab[18][25] ) );
  NOR2_X1 U13408 ( .A1(n3469), .A2(n3355), .ZN(\mult_20/ab[18][24] ) );
  NOR2_X1 U13409 ( .A1(n3268), .A2(n3180), .ZN(\mult_19/ab[22][19] ) );
  NOR2_X1 U13410 ( .A1(n3265), .A2(n3180), .ZN(\mult_19/ab[22][18] ) );
  NOR2_X1 U13411 ( .A1(n3262), .A2(n3180), .ZN(\mult_19/ab[22][17] ) );
  NOR2_X1 U13412 ( .A1(n3259), .A2(n3180), .ZN(\mult_19/ab[22][16] ) );
  NOR2_X1 U13413 ( .A1(n3256), .A2(n3180), .ZN(\mult_19/ab[22][15] ) );
  NOR2_X1 U13414 ( .A1(n3253), .A2(n3180), .ZN(\mult_19/ab[22][14] ) );
  NOR2_X1 U13415 ( .A1(n3250), .A2(n3180), .ZN(\mult_19/ab[22][13] ) );
  NOR2_X1 U13416 ( .A1(n3247), .A2(n3180), .ZN(\mult_19/ab[22][12] ) );
  NOR2_X1 U13417 ( .A1(n3244), .A2(n3180), .ZN(\mult_19/ab[22][11] ) );
  NOR2_X1 U13418 ( .A1(n3241), .A2(n3180), .ZN(\mult_19/ab[22][10] ) );
  NOR2_X1 U13419 ( .A1(n3289), .A2(n3169), .ZN(\mult_19/ab[18][26] ) );
  NOR2_X1 U13420 ( .A1(n3286), .A2(n3169), .ZN(\mult_19/ab[18][25] ) );
  NOR2_X1 U13421 ( .A1(n3283), .A2(n3169), .ZN(\mult_19/ab[18][24] ) );
  NOR2_X1 U13422 ( .A1(n3451), .A2(n3369), .ZN(\mult_20/ab[23][18] ) );
  NOR2_X1 U13423 ( .A1(n3448), .A2(n3369), .ZN(\mult_20/ab[23][17] ) );
  NOR2_X1 U13424 ( .A1(n3445), .A2(n3369), .ZN(\mult_20/ab[23][16] ) );
  NOR2_X1 U13425 ( .A1(n3442), .A2(n3369), .ZN(\mult_20/ab[23][15] ) );
  NOR2_X1 U13426 ( .A1(n3439), .A2(n3369), .ZN(\mult_20/ab[23][14] ) );
  NOR2_X1 U13427 ( .A1(n3436), .A2(n3369), .ZN(\mult_20/ab[23][13] ) );
  NOR2_X1 U13428 ( .A1(n3433), .A2(n3369), .ZN(\mult_20/ab[23][12] ) );
  NOR2_X1 U13429 ( .A1(n3430), .A2(n3369), .ZN(\mult_20/ab[23][11] ) );
  NOR2_X1 U13430 ( .A1(n3427), .A2(n3369), .ZN(\mult_20/ab[23][10] ) );
  NOR2_X1 U13431 ( .A1(n3472), .A2(n3358), .ZN(\mult_20/ab[19][25] ) );
  NOR2_X1 U13432 ( .A1(n3469), .A2(n3358), .ZN(\mult_20/ab[19][24] ) );
  NOR2_X1 U13433 ( .A1(n3466), .A2(n3358), .ZN(\mult_20/ab[19][23] ) );
  NOR2_X1 U13434 ( .A1(n3265), .A2(n3183), .ZN(\mult_19/ab[23][18] ) );
  NOR2_X1 U13435 ( .A1(n3262), .A2(n3183), .ZN(\mult_19/ab[23][17] ) );
  NOR2_X1 U13436 ( .A1(n3259), .A2(n3183), .ZN(\mult_19/ab[23][16] ) );
  NOR2_X1 U13437 ( .A1(n3256), .A2(n3183), .ZN(\mult_19/ab[23][15] ) );
  NOR2_X1 U13438 ( .A1(n3253), .A2(n3183), .ZN(\mult_19/ab[23][14] ) );
  NOR2_X1 U13439 ( .A1(n3250), .A2(n3183), .ZN(\mult_19/ab[23][13] ) );
  NOR2_X1 U13440 ( .A1(n3247), .A2(n3183), .ZN(\mult_19/ab[23][12] ) );
  NOR2_X1 U13441 ( .A1(n3244), .A2(n3183), .ZN(\mult_19/ab[23][11] ) );
  NOR2_X1 U13442 ( .A1(n3241), .A2(n3183), .ZN(\mult_19/ab[23][10] ) );
  NOR2_X1 U13443 ( .A1(n3286), .A2(n3172), .ZN(\mult_19/ab[19][25] ) );
  NOR2_X1 U13444 ( .A1(n3283), .A2(n3172), .ZN(\mult_19/ab[19][24] ) );
  NOR2_X1 U13445 ( .A1(n3280), .A2(n3172), .ZN(\mult_19/ab[19][23] ) );
  NOR2_X1 U13446 ( .A1(n3423), .A2(n3311), .ZN(\mult_20/ab[3][9] ) );
  NOR2_X1 U13447 ( .A1(n3417), .A2(n3311), .ZN(\mult_20/ab[3][7] ) );
  NOR2_X1 U13448 ( .A1(n3411), .A2(n3311), .ZN(\mult_20/ab[3][5] ) );
  NOR2_X1 U13449 ( .A1(n3448), .A2(n3372), .ZN(\mult_20/ab[24][17] ) );
  NOR2_X1 U13450 ( .A1(n3445), .A2(n3372), .ZN(\mult_20/ab[24][16] ) );
  NOR2_X1 U13451 ( .A1(n3442), .A2(n3372), .ZN(\mult_20/ab[24][15] ) );
  NOR2_X1 U13452 ( .A1(n3439), .A2(n3372), .ZN(\mult_20/ab[24][14] ) );
  NOR2_X1 U13453 ( .A1(n3436), .A2(n3372), .ZN(\mult_20/ab[24][13] ) );
  NOR2_X1 U13454 ( .A1(n3433), .A2(n3372), .ZN(\mult_20/ab[24][12] ) );
  NOR2_X1 U13455 ( .A1(n3430), .A2(n3372), .ZN(\mult_20/ab[24][11] ) );
  NOR2_X1 U13456 ( .A1(n3427), .A2(n3372), .ZN(\mult_20/ab[24][10] ) );
  NOR2_X1 U13457 ( .A1(n3469), .A2(n3361), .ZN(\mult_20/ab[20][24] ) );
  NOR2_X1 U13458 ( .A1(n3466), .A2(n3361), .ZN(\mult_20/ab[20][23] ) );
  NOR2_X1 U13459 ( .A1(n3463), .A2(n3361), .ZN(\mult_20/ab[20][22] ) );
  NOR2_X1 U13460 ( .A1(n3222), .A2(n3125), .ZN(\mult_19/ab[3][4] ) );
  NOR2_X1 U13461 ( .A1(n3219), .A2(n3125), .ZN(\mult_19/ab[3][3] ) );
  NOR2_X1 U13462 ( .A1(n3237), .A2(n3125), .ZN(\mult_19/ab[3][9] ) );
  NOR2_X1 U13463 ( .A1(n3234), .A2(n3125), .ZN(\mult_19/ab[3][8] ) );
  NOR2_X1 U13464 ( .A1(n3231), .A2(n3125), .ZN(\mult_19/ab[3][7] ) );
  NOR2_X1 U13465 ( .A1(n3228), .A2(n3125), .ZN(\mult_19/ab[3][6] ) );
  NOR2_X1 U13466 ( .A1(n3225), .A2(n3125), .ZN(\mult_19/ab[3][5] ) );
  NOR2_X1 U13467 ( .A1(n3262), .A2(n3186), .ZN(\mult_19/ab[24][17] ) );
  NOR2_X1 U13468 ( .A1(n3259), .A2(n3186), .ZN(\mult_19/ab[24][16] ) );
  NOR2_X1 U13469 ( .A1(n3256), .A2(n3186), .ZN(\mult_19/ab[24][15] ) );
  NOR2_X1 U13470 ( .A1(n3253), .A2(n3186), .ZN(\mult_19/ab[24][14] ) );
  NOR2_X1 U13471 ( .A1(n3250), .A2(n3186), .ZN(\mult_19/ab[24][13] ) );
  NOR2_X1 U13472 ( .A1(n3247), .A2(n3186), .ZN(\mult_19/ab[24][12] ) );
  NOR2_X1 U13473 ( .A1(n3244), .A2(n3186), .ZN(\mult_19/ab[24][11] ) );
  NOR2_X1 U13474 ( .A1(n3241), .A2(n3186), .ZN(\mult_19/ab[24][10] ) );
  NOR2_X1 U13475 ( .A1(n3283), .A2(n3175), .ZN(\mult_19/ab[20][24] ) );
  NOR2_X1 U13476 ( .A1(n3280), .A2(n3175), .ZN(\mult_19/ab[20][23] ) );
  NOR2_X1 U13477 ( .A1(n3277), .A2(n3175), .ZN(\mult_19/ab[20][22] ) );
  NOR2_X1 U13478 ( .A1(n3405), .A2(n3311), .ZN(\mult_20/ab[3][3] ) );
  NOR2_X1 U13479 ( .A1(n3423), .A2(n3314), .ZN(\mult_20/ab[4][9] ) );
  NOR2_X1 U13480 ( .A1(n3417), .A2(n3314), .ZN(\mult_20/ab[4][7] ) );
  NOR2_X1 U13481 ( .A1(n3411), .A2(n3314), .ZN(\mult_20/ab[4][5] ) );
  NOR2_X1 U13482 ( .A1(n3445), .A2(n3375), .ZN(\mult_20/ab[25][16] ) );
  NOR2_X1 U13483 ( .A1(n3442), .A2(n3375), .ZN(\mult_20/ab[25][15] ) );
  NOR2_X1 U13484 ( .A1(n3439), .A2(n3375), .ZN(\mult_20/ab[25][14] ) );
  NOR2_X1 U13485 ( .A1(n3436), .A2(n3375), .ZN(\mult_20/ab[25][13] ) );
  NOR2_X1 U13486 ( .A1(n3433), .A2(n3375), .ZN(\mult_20/ab[25][12] ) );
  NOR2_X1 U13487 ( .A1(n3430), .A2(n3375), .ZN(\mult_20/ab[25][11] ) );
  NOR2_X1 U13488 ( .A1(n3427), .A2(n3375), .ZN(\mult_20/ab[25][10] ) );
  NOR2_X1 U13489 ( .A1(n3466), .A2(n3364), .ZN(\mult_20/ab[21][23] ) );
  NOR2_X1 U13490 ( .A1(n3463), .A2(n3364), .ZN(\mult_20/ab[21][22] ) );
  NOR2_X1 U13491 ( .A1(n3460), .A2(n3364), .ZN(\mult_20/ab[21][21] ) );
  NOR2_X1 U13492 ( .A1(n3259), .A2(n3189), .ZN(\mult_19/ab[25][16] ) );
  NOR2_X1 U13493 ( .A1(n3256), .A2(n3189), .ZN(\mult_19/ab[25][15] ) );
  NOR2_X1 U13494 ( .A1(n3253), .A2(n3189), .ZN(\mult_19/ab[25][14] ) );
  NOR2_X1 U13495 ( .A1(n3250), .A2(n3189), .ZN(\mult_19/ab[25][13] ) );
  NOR2_X1 U13496 ( .A1(n3247), .A2(n3189), .ZN(\mult_19/ab[25][12] ) );
  NOR2_X1 U13497 ( .A1(n3244), .A2(n3189), .ZN(\mult_19/ab[25][11] ) );
  NOR2_X1 U13498 ( .A1(n3241), .A2(n3189), .ZN(\mult_19/ab[25][10] ) );
  NOR2_X1 U13499 ( .A1(n3280), .A2(n3178), .ZN(\mult_19/ab[21][23] ) );
  NOR2_X1 U13500 ( .A1(n3277), .A2(n3178), .ZN(\mult_19/ab[21][22] ) );
  NOR2_X1 U13501 ( .A1(n3274), .A2(n3178), .ZN(\mult_19/ab[21][21] ) );
  NOR2_X1 U13502 ( .A1(n3405), .A2(n3314), .ZN(\mult_20/ab[4][3] ) );
  NOR2_X1 U13503 ( .A1(n3423), .A2(n3317), .ZN(\mult_20/ab[5][9] ) );
  NOR2_X1 U13504 ( .A1(n3417), .A2(n3317), .ZN(\mult_20/ab[5][7] ) );
  NOR2_X1 U13505 ( .A1(n3411), .A2(n3317), .ZN(\mult_20/ab[5][5] ) );
  NOR2_X1 U13506 ( .A1(n3442), .A2(n3378), .ZN(\mult_20/ab[26][15] ) );
  NOR2_X1 U13507 ( .A1(n3439), .A2(n3378), .ZN(\mult_20/ab[26][14] ) );
  NOR2_X1 U13508 ( .A1(n3436), .A2(n3378), .ZN(\mult_20/ab[26][13] ) );
  NOR2_X1 U13509 ( .A1(n3433), .A2(n3378), .ZN(\mult_20/ab[26][12] ) );
  NOR2_X1 U13510 ( .A1(n3430), .A2(n3378), .ZN(\mult_20/ab[26][11] ) );
  NOR2_X1 U13511 ( .A1(n3427), .A2(n3378), .ZN(\mult_20/ab[26][10] ) );
  NOR2_X1 U13512 ( .A1(n3463), .A2(n3367), .ZN(\mult_20/ab[22][22] ) );
  NOR2_X1 U13513 ( .A1(n3460), .A2(n3367), .ZN(\mult_20/ab[22][21] ) );
  NOR2_X1 U13514 ( .A1(n3457), .A2(n3367), .ZN(\mult_20/ab[22][20] ) );
  NOR2_X1 U13515 ( .A1(n3222), .A2(n3131), .ZN(\mult_19/ab[5][4] ) );
  NOR2_X1 U13516 ( .A1(n3219), .A2(n3131), .ZN(\mult_19/ab[5][3] ) );
  NOR2_X1 U13517 ( .A1(n3237), .A2(n3131), .ZN(\mult_19/ab[5][9] ) );
  NOR2_X1 U13518 ( .A1(n3234), .A2(n3131), .ZN(\mult_19/ab[5][8] ) );
  NOR2_X1 U13519 ( .A1(n3231), .A2(n3131), .ZN(\mult_19/ab[5][7] ) );
  NOR2_X1 U13520 ( .A1(n3228), .A2(n3131), .ZN(\mult_19/ab[5][6] ) );
  NOR2_X1 U13521 ( .A1(n3225), .A2(n3131), .ZN(\mult_19/ab[5][5] ) );
  NOR2_X1 U13522 ( .A1(n3256), .A2(n3192), .ZN(\mult_19/ab[26][15] ) );
  NOR2_X1 U13523 ( .A1(n3253), .A2(n3192), .ZN(\mult_19/ab[26][14] ) );
  NOR2_X1 U13524 ( .A1(n3250), .A2(n3192), .ZN(\mult_19/ab[26][13] ) );
  NOR2_X1 U13525 ( .A1(n3247), .A2(n3192), .ZN(\mult_19/ab[26][12] ) );
  NOR2_X1 U13526 ( .A1(n3244), .A2(n3192), .ZN(\mult_19/ab[26][11] ) );
  NOR2_X1 U13527 ( .A1(n3241), .A2(n3192), .ZN(\mult_19/ab[26][10] ) );
  NOR2_X1 U13528 ( .A1(n3277), .A2(n3181), .ZN(\mult_19/ab[22][22] ) );
  NOR2_X1 U13529 ( .A1(n3274), .A2(n3181), .ZN(\mult_19/ab[22][21] ) );
  NOR2_X1 U13530 ( .A1(n3271), .A2(n3181), .ZN(\mult_19/ab[22][20] ) );
  NOR2_X1 U13531 ( .A1(n3405), .A2(n3317), .ZN(\mult_20/ab[5][3] ) );
  NOR2_X1 U13532 ( .A1(n3423), .A2(n3320), .ZN(\mult_20/ab[6][9] ) );
  NOR2_X1 U13533 ( .A1(n3417), .A2(n3320), .ZN(\mult_20/ab[6][7] ) );
  NOR2_X1 U13534 ( .A1(n3411), .A2(n3320), .ZN(\mult_20/ab[6][5] ) );
  NOR2_X1 U13535 ( .A1(n3439), .A2(n3381), .ZN(\mult_20/ab[27][14] ) );
  NOR2_X1 U13536 ( .A1(n3436), .A2(n3381), .ZN(\mult_20/ab[27][13] ) );
  NOR2_X1 U13537 ( .A1(n3433), .A2(n3381), .ZN(\mult_20/ab[27][12] ) );
  NOR2_X1 U13538 ( .A1(n3430), .A2(n3381), .ZN(\mult_20/ab[27][11] ) );
  NOR2_X1 U13539 ( .A1(n3427), .A2(n3381), .ZN(\mult_20/ab[27][10] ) );
  NOR2_X1 U13540 ( .A1(n3460), .A2(n3370), .ZN(\mult_20/ab[23][21] ) );
  NOR2_X1 U13541 ( .A1(n3457), .A2(n3370), .ZN(\mult_20/ab[23][20] ) );
  NOR2_X1 U13542 ( .A1(n3454), .A2(n3369), .ZN(\mult_20/ab[23][19] ) );
  NOR2_X1 U13543 ( .A1(n3253), .A2(n3195), .ZN(\mult_19/ab[27][14] ) );
  NOR2_X1 U13544 ( .A1(n3250), .A2(n3195), .ZN(\mult_19/ab[27][13] ) );
  NOR2_X1 U13545 ( .A1(n3247), .A2(n3195), .ZN(\mult_19/ab[27][12] ) );
  NOR2_X1 U13546 ( .A1(n3244), .A2(n3195), .ZN(\mult_19/ab[27][11] ) );
  NOR2_X1 U13547 ( .A1(n3241), .A2(n3195), .ZN(\mult_19/ab[27][10] ) );
  NOR2_X1 U13548 ( .A1(n3274), .A2(n3184), .ZN(\mult_19/ab[23][21] ) );
  NOR2_X1 U13549 ( .A1(n3271), .A2(n3184), .ZN(\mult_19/ab[23][20] ) );
  NOR2_X1 U13550 ( .A1(n3268), .A2(n3183), .ZN(\mult_19/ab[23][19] ) );
  NOR2_X1 U13551 ( .A1(n3405), .A2(n3320), .ZN(\mult_20/ab[6][3] ) );
  NOR2_X1 U13552 ( .A1(n3423), .A2(n3323), .ZN(\mult_20/ab[7][9] ) );
  NOR2_X1 U13553 ( .A1(n3417), .A2(n3323), .ZN(\mult_20/ab[7][7] ) );
  NOR2_X1 U13554 ( .A1(n3411), .A2(n3323), .ZN(\mult_20/ab[7][5] ) );
  NOR2_X1 U13555 ( .A1(n3436), .A2(n3384), .ZN(\mult_20/ab[28][13] ) );
  NOR2_X1 U13556 ( .A1(n3433), .A2(n3384), .ZN(\mult_20/ab[28][12] ) );
  NOR2_X1 U13557 ( .A1(n3430), .A2(n3384), .ZN(\mult_20/ab[28][11] ) );
  NOR2_X1 U13558 ( .A1(n3427), .A2(n3384), .ZN(\mult_20/ab[28][10] ) );
  NOR2_X1 U13559 ( .A1(n3457), .A2(n3373), .ZN(\mult_20/ab[24][20] ) );
  NOR2_X1 U13560 ( .A1(n3454), .A2(n3372), .ZN(\mult_20/ab[24][19] ) );
  NOR2_X1 U13561 ( .A1(n3451), .A2(n3372), .ZN(\mult_20/ab[24][18] ) );
  NOR2_X1 U13562 ( .A1(n3222), .A2(n3137), .ZN(\mult_19/ab[7][4] ) );
  NOR2_X1 U13563 ( .A1(n3219), .A2(n3137), .ZN(\mult_19/ab[7][3] ) );
  NOR2_X1 U13564 ( .A1(n3237), .A2(n3137), .ZN(\mult_19/ab[7][9] ) );
  NOR2_X1 U13565 ( .A1(n3234), .A2(n3137), .ZN(\mult_19/ab[7][8] ) );
  NOR2_X1 U13566 ( .A1(n3231), .A2(n3137), .ZN(\mult_19/ab[7][7] ) );
  NOR2_X1 U13567 ( .A1(n3228), .A2(n3137), .ZN(\mult_19/ab[7][6] ) );
  NOR2_X1 U13568 ( .A1(n3225), .A2(n3137), .ZN(\mult_19/ab[7][5] ) );
  NOR2_X1 U13569 ( .A1(n3250), .A2(n3198), .ZN(\mult_19/ab[28][13] ) );
  NOR2_X1 U13570 ( .A1(n3247), .A2(n3198), .ZN(\mult_19/ab[28][12] ) );
  NOR2_X1 U13571 ( .A1(n3244), .A2(n3198), .ZN(\mult_19/ab[28][11] ) );
  NOR2_X1 U13572 ( .A1(n3241), .A2(n3198), .ZN(\mult_19/ab[28][10] ) );
  NOR2_X1 U13573 ( .A1(n3271), .A2(n3187), .ZN(\mult_19/ab[24][20] ) );
  NOR2_X1 U13574 ( .A1(n3268), .A2(n3186), .ZN(\mult_19/ab[24][19] ) );
  NOR2_X1 U13575 ( .A1(n3265), .A2(n3186), .ZN(\mult_19/ab[24][18] ) );
  NOR2_X1 U13576 ( .A1(n3405), .A2(n3323), .ZN(\mult_20/ab[7][3] ) );
  NOR2_X1 U13577 ( .A1(n3423), .A2(n3326), .ZN(\mult_20/ab[8][9] ) );
  NOR2_X1 U13578 ( .A1(n3417), .A2(n3326), .ZN(\mult_20/ab[8][7] ) );
  NOR2_X1 U13579 ( .A1(n3411), .A2(n3326), .ZN(\mult_20/ab[8][5] ) );
  NOR2_X1 U13580 ( .A1(n3432), .A2(n3387), .ZN(\mult_20/ab[29][12] ) );
  NOR2_X1 U13581 ( .A1(n3429), .A2(n3387), .ZN(\mult_20/ab[29][11] ) );
  NOR2_X1 U13582 ( .A1(n3426), .A2(n3387), .ZN(\mult_20/ab[29][10] ) );
  NOR2_X1 U13583 ( .A1(n3454), .A2(n3375), .ZN(\mult_20/ab[25][19] ) );
  NOR2_X1 U13584 ( .A1(n3451), .A2(n3375), .ZN(\mult_20/ab[25][18] ) );
  NOR2_X1 U13585 ( .A1(n3448), .A2(n3375), .ZN(\mult_20/ab[25][17] ) );
  NOR2_X1 U13586 ( .A1(n3246), .A2(n3201), .ZN(\mult_19/ab[29][12] ) );
  NOR2_X1 U13587 ( .A1(n3243), .A2(n3201), .ZN(\mult_19/ab[29][11] ) );
  NOR2_X1 U13588 ( .A1(n3240), .A2(n3201), .ZN(\mult_19/ab[29][10] ) );
  NOR2_X1 U13589 ( .A1(n3268), .A2(n3189), .ZN(\mult_19/ab[25][19] ) );
  NOR2_X1 U13590 ( .A1(n3265), .A2(n3189), .ZN(\mult_19/ab[25][18] ) );
  NOR2_X1 U13591 ( .A1(n3262), .A2(n3189), .ZN(\mult_19/ab[25][17] ) );
  NOR2_X1 U13592 ( .A1(n3405), .A2(n3326), .ZN(\mult_20/ab[8][3] ) );
  NOR2_X1 U13593 ( .A1(n3423), .A2(n3329), .ZN(\mult_20/ab[9][9] ) );
  NOR2_X1 U13594 ( .A1(n3417), .A2(n3329), .ZN(\mult_20/ab[9][7] ) );
  NOR2_X1 U13595 ( .A1(n3411), .A2(n3329), .ZN(\mult_20/ab[9][5] ) );
  NOR2_X1 U13596 ( .A1(n3429), .A2(n3390), .ZN(\mult_20/ab[30][11] ) );
  NOR2_X1 U13597 ( .A1(n3426), .A2(n3390), .ZN(\mult_20/ab[30][10] ) );
  NOR2_X1 U13598 ( .A1(n3451), .A2(n3378), .ZN(\mult_20/ab[26][18] ) );
  NOR2_X1 U13599 ( .A1(n3448), .A2(n3378), .ZN(\mult_20/ab[26][17] ) );
  NOR2_X1 U13600 ( .A1(n3445), .A2(n3378), .ZN(\mult_20/ab[26][16] ) );
  NOR2_X1 U13601 ( .A1(n3222), .A2(n3143), .ZN(\mult_19/ab[9][4] ) );
  NOR2_X1 U13602 ( .A1(n3219), .A2(n3143), .ZN(\mult_19/ab[9][3] ) );
  NOR2_X1 U13603 ( .A1(n3237), .A2(n3143), .ZN(\mult_19/ab[9][9] ) );
  NOR2_X1 U13604 ( .A1(n3234), .A2(n3143), .ZN(\mult_19/ab[9][8] ) );
  NOR2_X1 U13605 ( .A1(n3231), .A2(n3143), .ZN(\mult_19/ab[9][7] ) );
  NOR2_X1 U13606 ( .A1(n3228), .A2(n3143), .ZN(\mult_19/ab[9][6] ) );
  NOR2_X1 U13607 ( .A1(n3225), .A2(n3143), .ZN(\mult_19/ab[9][5] ) );
  NOR2_X1 U13608 ( .A1(n3243), .A2(n3204), .ZN(\mult_19/ab[30][11] ) );
  NOR2_X1 U13609 ( .A1(n3240), .A2(n3204), .ZN(\mult_19/ab[30][10] ) );
  NOR2_X1 U13610 ( .A1(n3265), .A2(n3192), .ZN(\mult_19/ab[26][18] ) );
  NOR2_X1 U13611 ( .A1(n3262), .A2(n3192), .ZN(\mult_19/ab[26][17] ) );
  NOR2_X1 U13612 ( .A1(n3259), .A2(n3192), .ZN(\mult_19/ab[26][16] ) );
  NOR2_X1 U13613 ( .A1(n3405), .A2(n3329), .ZN(\mult_20/ab[9][3] ) );
  NOR2_X1 U13614 ( .A1(n3425), .A2(n3332), .ZN(\mult_20/ab[10][9] ) );
  NOR2_X1 U13615 ( .A1(n3419), .A2(n3332), .ZN(\mult_20/ab[10][7] ) );
  NOR2_X1 U13616 ( .A1(n3413), .A2(n3332), .ZN(\mult_20/ab[10][5] ) );
  NOR2_X1 U13617 ( .A1(n3448), .A2(n3381), .ZN(\mult_20/ab[27][17] ) );
  NOR2_X1 U13618 ( .A1(n3445), .A2(n3381), .ZN(\mult_20/ab[27][16] ) );
  NOR2_X1 U13619 ( .A1(n3442), .A2(n3381), .ZN(\mult_20/ab[27][15] ) );
  NOR2_X1 U13620 ( .A1(n3262), .A2(n3195), .ZN(\mult_19/ab[27][17] ) );
  NOR2_X1 U13621 ( .A1(n3259), .A2(n3195), .ZN(\mult_19/ab[27][16] ) );
  NOR2_X1 U13622 ( .A1(n3256), .A2(n3195), .ZN(\mult_19/ab[27][15] ) );
  NOR2_X1 U13623 ( .A1(n3407), .A2(n3332), .ZN(\mult_20/ab[10][3] ) );
  NOR2_X1 U13624 ( .A1(n3425), .A2(n3335), .ZN(\mult_20/ab[11][9] ) );
  NOR2_X1 U13625 ( .A1(n3419), .A2(n3335), .ZN(\mult_20/ab[11][7] ) );
  NOR2_X1 U13626 ( .A1(n3413), .A2(n3335), .ZN(\mult_20/ab[11][5] ) );
  NOR2_X1 U13627 ( .A1(n3445), .A2(n3384), .ZN(\mult_20/ab[28][16] ) );
  NOR2_X1 U13628 ( .A1(n3439), .A2(n3384), .ZN(\mult_20/ab[28][14] ) );
  NOR2_X1 U13629 ( .A1(n3442), .A2(n3384), .ZN(\mult_20/ab[28][15] ) );
  NOR2_X1 U13630 ( .A1(n3224), .A2(n3149), .ZN(\mult_19/ab[11][4] ) );
  NOR2_X1 U13631 ( .A1(n3221), .A2(n3149), .ZN(\mult_19/ab[11][3] ) );
  NOR2_X1 U13632 ( .A1(n3239), .A2(n3149), .ZN(\mult_19/ab[11][9] ) );
  NOR2_X1 U13633 ( .A1(n3236), .A2(n3149), .ZN(\mult_19/ab[11][8] ) );
  NOR2_X1 U13634 ( .A1(n3233), .A2(n3149), .ZN(\mult_19/ab[11][7] ) );
  NOR2_X1 U13635 ( .A1(n3230), .A2(n3149), .ZN(\mult_19/ab[11][6] ) );
  NOR2_X1 U13636 ( .A1(n3227), .A2(n3149), .ZN(\mult_19/ab[11][5] ) );
  NOR2_X1 U13637 ( .A1(n3259), .A2(n3198), .ZN(\mult_19/ab[28][16] ) );
  NOR2_X1 U13638 ( .A1(n3253), .A2(n3198), .ZN(\mult_19/ab[28][14] ) );
  NOR2_X1 U13639 ( .A1(n3256), .A2(n3198), .ZN(\mult_19/ab[28][15] ) );
  NOR2_X1 U13640 ( .A1(n3407), .A2(n3335), .ZN(\mult_20/ab[11][3] ) );
  NOR2_X1 U13641 ( .A1(n3425), .A2(n3338), .ZN(\mult_20/ab[12][9] ) );
  NOR2_X1 U13642 ( .A1(n3419), .A2(n3338), .ZN(\mult_20/ab[12][7] ) );
  NOR2_X1 U13643 ( .A1(n3413), .A2(n3338), .ZN(\mult_20/ab[12][5] ) );
  NOR2_X1 U13644 ( .A1(n3435), .A2(n3387), .ZN(\mult_20/ab[29][13] ) );
  NOR2_X1 U13645 ( .A1(n3441), .A2(n3387), .ZN(\mult_20/ab[29][15] ) );
  NOR2_X1 U13646 ( .A1(n3438), .A2(n3387), .ZN(\mult_20/ab[29][14] ) );
  NOR2_X1 U13647 ( .A1(n3249), .A2(n3201), .ZN(\mult_19/ab[29][13] ) );
  NOR2_X1 U13648 ( .A1(n3255), .A2(n3201), .ZN(\mult_19/ab[29][15] ) );
  NOR2_X1 U13649 ( .A1(n3252), .A2(n3201), .ZN(\mult_19/ab[29][14] ) );
  NOR2_X1 U13650 ( .A1(n3407), .A2(n3338), .ZN(\mult_20/ab[12][3] ) );
  NOR2_X1 U13651 ( .A1(n3425), .A2(n3341), .ZN(\mult_20/ab[13][9] ) );
  NOR2_X1 U13652 ( .A1(n3419), .A2(n3341), .ZN(\mult_20/ab[13][7] ) );
  NOR2_X1 U13653 ( .A1(n3413), .A2(n3341), .ZN(\mult_20/ab[13][5] ) );
  NOR2_X1 U13654 ( .A1(n3435), .A2(n3390), .ZN(\mult_20/ab[30][13] ) );
  NOR2_X1 U13655 ( .A1(n3438), .A2(n3390), .ZN(\mult_20/ab[30][14] ) );
  NOR2_X1 U13656 ( .A1(n3224), .A2(n3155), .ZN(\mult_19/ab[13][4] ) );
  NOR2_X1 U13657 ( .A1(n3221), .A2(n3155), .ZN(\mult_19/ab[13][3] ) );
  NOR2_X1 U13658 ( .A1(n3239), .A2(n3155), .ZN(\mult_19/ab[13][9] ) );
  NOR2_X1 U13659 ( .A1(n3236), .A2(n3155), .ZN(\mult_19/ab[13][8] ) );
  NOR2_X1 U13660 ( .A1(n3233), .A2(n3155), .ZN(\mult_19/ab[13][7] ) );
  NOR2_X1 U13661 ( .A1(n3230), .A2(n3155), .ZN(\mult_19/ab[13][6] ) );
  NOR2_X1 U13662 ( .A1(n3227), .A2(n3155), .ZN(\mult_19/ab[13][5] ) );
  NOR2_X1 U13663 ( .A1(n3249), .A2(n3204), .ZN(\mult_19/ab[30][13] ) );
  NOR2_X1 U13664 ( .A1(n3252), .A2(n3204), .ZN(\mult_19/ab[30][14] ) );
  NOR2_X1 U13665 ( .A1(n3407), .A2(n3341), .ZN(\mult_20/ab[13][3] ) );
  NOR2_X1 U13666 ( .A1(n3425), .A2(n3344), .ZN(\mult_20/ab[14][9] ) );
  NOR2_X1 U13667 ( .A1(n3419), .A2(n3344), .ZN(\mult_20/ab[14][7] ) );
  NOR2_X1 U13668 ( .A1(n3413), .A2(n3344), .ZN(\mult_20/ab[14][5] ) );
  NOR2_X1 U13669 ( .A1(n3407), .A2(n3344), .ZN(\mult_20/ab[14][3] ) );
  NOR2_X1 U13670 ( .A1(n3425), .A2(n3347), .ZN(\mult_20/ab[15][9] ) );
  NOR2_X1 U13671 ( .A1(n3419), .A2(n3347), .ZN(\mult_20/ab[15][7] ) );
  NOR2_X1 U13672 ( .A1(n3413), .A2(n3347), .ZN(\mult_20/ab[15][5] ) );
  NOR2_X1 U13673 ( .A1(n3224), .A2(n3161), .ZN(\mult_19/ab[15][4] ) );
  NOR2_X1 U13674 ( .A1(n3221), .A2(n3161), .ZN(\mult_19/ab[15][3] ) );
  NOR2_X1 U13675 ( .A1(n3239), .A2(n3161), .ZN(\mult_19/ab[15][9] ) );
  NOR2_X1 U13676 ( .A1(n3236), .A2(n3161), .ZN(\mult_19/ab[15][8] ) );
  NOR2_X1 U13677 ( .A1(n3233), .A2(n3161), .ZN(\mult_19/ab[15][7] ) );
  NOR2_X1 U13678 ( .A1(n3230), .A2(n3161), .ZN(\mult_19/ab[15][6] ) );
  NOR2_X1 U13679 ( .A1(n3227), .A2(n3161), .ZN(\mult_19/ab[15][5] ) );
  NOR2_X1 U13680 ( .A1(n3407), .A2(n3347), .ZN(\mult_20/ab[15][3] ) );
  NOR2_X1 U13681 ( .A1(n3425), .A2(n3350), .ZN(\mult_20/ab[16][9] ) );
  NOR2_X1 U13682 ( .A1(n3419), .A2(n3350), .ZN(\mult_20/ab[16][7] ) );
  NOR2_X1 U13683 ( .A1(n3413), .A2(n3350), .ZN(\mult_20/ab[16][5] ) );
  NOR2_X1 U13684 ( .A1(n3239), .A2(n3164), .ZN(\mult_19/ab[16][9] ) );
  NOR2_X1 U13685 ( .A1(n3407), .A2(n3350), .ZN(\mult_20/ab[16][3] ) );
  NOR2_X1 U13686 ( .A1(n3424), .A2(n3353), .ZN(\mult_20/ab[17][9] ) );
  NOR2_X1 U13687 ( .A1(n3418), .A2(n3353), .ZN(\mult_20/ab[17][7] ) );
  NOR2_X1 U13688 ( .A1(n3412), .A2(n3353), .ZN(\mult_20/ab[17][5] ) );
  NOR2_X1 U13689 ( .A1(n3223), .A2(n3167), .ZN(\mult_19/ab[17][4] ) );
  NOR2_X1 U13690 ( .A1(n3220), .A2(n3167), .ZN(\mult_19/ab[17][3] ) );
  NOR2_X1 U13691 ( .A1(n3232), .A2(n3167), .ZN(\mult_19/ab[17][7] ) );
  NOR2_X1 U13692 ( .A1(n3229), .A2(n3167), .ZN(\mult_19/ab[17][6] ) );
  NOR2_X1 U13693 ( .A1(n3226), .A2(n3167), .ZN(\mult_19/ab[17][5] ) );
  NOR2_X1 U13694 ( .A1(n3406), .A2(n3353), .ZN(\mult_20/ab[17][3] ) );
  NOR2_X1 U13695 ( .A1(n3424), .A2(n3356), .ZN(\mult_20/ab[18][9] ) );
  NOR2_X1 U13696 ( .A1(n3418), .A2(n3356), .ZN(\mult_20/ab[18][7] ) );
  NOR2_X1 U13697 ( .A1(n3412), .A2(n3356), .ZN(\mult_20/ab[18][5] ) );
  NOR2_X1 U13698 ( .A1(n3238), .A2(n3170), .ZN(\mult_19/ab[18][9] ) );
  NOR2_X1 U13699 ( .A1(n3235), .A2(n3170), .ZN(\mult_19/ab[18][8] ) );
  NOR2_X1 U13700 ( .A1(n3232), .A2(n3170), .ZN(\mult_19/ab[18][7] ) );
  NOR2_X1 U13701 ( .A1(n3406), .A2(n3356), .ZN(\mult_20/ab[18][3] ) );
  NOR2_X1 U13702 ( .A1(n3424), .A2(n3359), .ZN(\mult_20/ab[19][9] ) );
  NOR2_X1 U13703 ( .A1(n3418), .A2(n3359), .ZN(\mult_20/ab[19][7] ) );
  NOR2_X1 U13704 ( .A1(n3412), .A2(n3359), .ZN(\mult_20/ab[19][5] ) );
  NOR2_X1 U13705 ( .A1(n3223), .A2(n3173), .ZN(\mult_19/ab[19][4] ) );
  NOR2_X1 U13706 ( .A1(n3220), .A2(n3173), .ZN(\mult_19/ab[19][3] ) );
  NOR2_X1 U13707 ( .A1(n3226), .A2(n3173), .ZN(\mult_19/ab[19][5] ) );
  NOR2_X1 U13708 ( .A1(n3406), .A2(n3359), .ZN(\mult_20/ab[19][3] ) );
  NOR2_X1 U13709 ( .A1(n3424), .A2(n3362), .ZN(\mult_20/ab[20][9] ) );
  NOR2_X1 U13710 ( .A1(n3418), .A2(n3362), .ZN(\mult_20/ab[20][7] ) );
  NOR2_X1 U13711 ( .A1(n3412), .A2(n3362), .ZN(\mult_20/ab[20][5] ) );
  NOR2_X1 U13712 ( .A1(n3238), .A2(n3176), .ZN(\mult_19/ab[20][9] ) );
  NOR2_X1 U13713 ( .A1(n3235), .A2(n3176), .ZN(\mult_19/ab[20][8] ) );
  NOR2_X1 U13714 ( .A1(n3232), .A2(n3176), .ZN(\mult_19/ab[20][7] ) );
  NOR2_X1 U13715 ( .A1(n3229), .A2(n3176), .ZN(\mult_19/ab[20][6] ) );
  NOR2_X1 U13716 ( .A1(n3226), .A2(n3176), .ZN(\mult_19/ab[20][5] ) );
  NOR2_X1 U13717 ( .A1(n3406), .A2(n3362), .ZN(\mult_20/ab[20][3] ) );
  NOR2_X1 U13718 ( .A1(n3424), .A2(n3365), .ZN(\mult_20/ab[21][9] ) );
  NOR2_X1 U13719 ( .A1(n3418), .A2(n3365), .ZN(\mult_20/ab[21][7] ) );
  NOR2_X1 U13720 ( .A1(n3412), .A2(n3365), .ZN(\mult_20/ab[21][5] ) );
  NOR2_X1 U13721 ( .A1(n3220), .A2(n3179), .ZN(\mult_19/ab[21][3] ) );
  NOR2_X1 U13722 ( .A1(n3406), .A2(n3365), .ZN(\mult_20/ab[21][3] ) );
  NOR2_X1 U13723 ( .A1(n3424), .A2(n3368), .ZN(\mult_20/ab[22][9] ) );
  NOR2_X1 U13724 ( .A1(n3418), .A2(n3368), .ZN(\mult_20/ab[22][7] ) );
  NOR2_X1 U13725 ( .A1(n3412), .A2(n3368), .ZN(\mult_20/ab[22][5] ) );
  NOR2_X1 U13726 ( .A1(n3223), .A2(n3182), .ZN(\mult_19/ab[22][4] ) );
  NOR2_X1 U13727 ( .A1(n3220), .A2(n3182), .ZN(\mult_19/ab[22][3] ) );
  NOR2_X1 U13728 ( .A1(n3235), .A2(n3182), .ZN(\mult_19/ab[22][8] ) );
  NOR2_X1 U13729 ( .A1(n3232), .A2(n3182), .ZN(\mult_19/ab[22][7] ) );
  NOR2_X1 U13730 ( .A1(n3229), .A2(n3182), .ZN(\mult_19/ab[22][6] ) );
  NOR2_X1 U13731 ( .A1(n3226), .A2(n3182), .ZN(\mult_19/ab[22][5] ) );
  NOR2_X1 U13732 ( .A1(n3406), .A2(n3368), .ZN(\mult_20/ab[22][3] ) );
  NOR2_X1 U13733 ( .A1(n3424), .A2(n3371), .ZN(\mult_20/ab[23][9] ) );
  NOR2_X1 U13734 ( .A1(n3418), .A2(n3371), .ZN(\mult_20/ab[23][7] ) );
  NOR2_X1 U13735 ( .A1(n3412), .A2(n3371), .ZN(\mult_20/ab[23][5] ) );
  NOR2_X1 U13736 ( .A1(n3235), .A2(n3185), .ZN(\mult_19/ab[23][8] ) );
  NOR2_X1 U13737 ( .A1(n3406), .A2(n3371), .ZN(\mult_20/ab[23][3] ) );
  NOR2_X1 U13738 ( .A1(n3424), .A2(n3374), .ZN(\mult_20/ab[24][9] ) );
  NOR2_X1 U13739 ( .A1(n3421), .A2(n3374), .ZN(\mult_20/ab[24][8] ) );
  NOR2_X1 U13740 ( .A1(n3418), .A2(n3374), .ZN(\mult_20/ab[24][7] ) );
  NOR2_X1 U13741 ( .A1(n3412), .A2(n3374), .ZN(\mult_20/ab[24][5] ) );
  NOR2_X1 U13742 ( .A1(n3223), .A2(n3188), .ZN(\mult_19/ab[24][4] ) );
  NOR2_X1 U13743 ( .A1(n3220), .A2(n3188), .ZN(\mult_19/ab[24][3] ) );
  NOR2_X1 U13744 ( .A1(n3238), .A2(n3188), .ZN(\mult_19/ab[24][9] ) );
  NOR2_X1 U13745 ( .A1(n3235), .A2(n3188), .ZN(\mult_19/ab[24][8] ) );
  NOR2_X1 U13746 ( .A1(n3229), .A2(n3188), .ZN(\mult_19/ab[24][6] ) );
  NOR2_X1 U13747 ( .A1(n3226), .A2(n3188), .ZN(\mult_19/ab[24][5] ) );
  NOR2_X1 U13748 ( .A1(n3406), .A2(n3374), .ZN(\mult_20/ab[24][3] ) );
  NOR2_X1 U13749 ( .A1(n3424), .A2(n3377), .ZN(\mult_20/ab[25][9] ) );
  NOR2_X1 U13750 ( .A1(n3421), .A2(n3377), .ZN(\mult_20/ab[25][8] ) );
  NOR2_X1 U13751 ( .A1(n3418), .A2(n3377), .ZN(\mult_20/ab[25][7] ) );
  NOR2_X1 U13752 ( .A1(n3412), .A2(n3377), .ZN(\mult_20/ab[25][5] ) );
  NOR2_X1 U13753 ( .A1(n3238), .A2(n3191), .ZN(\mult_19/ab[25][9] ) );
  NOR2_X1 U13754 ( .A1(n3235), .A2(n3191), .ZN(\mult_19/ab[25][8] ) );
  NOR2_X1 U13755 ( .A1(n3229), .A2(n3191), .ZN(\mult_19/ab[25][6] ) );
  NOR2_X1 U13756 ( .A1(n3406), .A2(n3377), .ZN(\mult_20/ab[25][3] ) );
  NOR2_X1 U13757 ( .A1(n3424), .A2(n3380), .ZN(\mult_20/ab[26][9] ) );
  NOR2_X1 U13758 ( .A1(n3421), .A2(n3380), .ZN(\mult_20/ab[26][8] ) );
  NOR2_X1 U13759 ( .A1(n3418), .A2(n3380), .ZN(\mult_20/ab[26][7] ) );
  NOR2_X1 U13760 ( .A1(n3415), .A2(n3380), .ZN(\mult_20/ab[26][6] ) );
  NOR2_X1 U13761 ( .A1(n3412), .A2(n3380), .ZN(\mult_20/ab[26][5] ) );
  NOR2_X1 U13762 ( .A1(n3223), .A2(n3194), .ZN(\mult_19/ab[26][4] ) );
  NOR2_X1 U13763 ( .A1(n3220), .A2(n3194), .ZN(\mult_19/ab[26][3] ) );
  NOR2_X1 U13764 ( .A1(n3238), .A2(n3194), .ZN(\mult_19/ab[26][9] ) );
  NOR2_X1 U13765 ( .A1(n3235), .A2(n3194), .ZN(\mult_19/ab[26][8] ) );
  NOR2_X1 U13766 ( .A1(n3232), .A2(n3194), .ZN(\mult_19/ab[26][7] ) );
  NOR2_X1 U13767 ( .A1(n3229), .A2(n3194), .ZN(\mult_19/ab[26][6] ) );
  NOR2_X1 U13768 ( .A1(n3406), .A2(n3380), .ZN(\mult_20/ab[26][3] ) );
  NOR2_X1 U13769 ( .A1(n3424), .A2(n3383), .ZN(\mult_20/ab[27][9] ) );
  NOR2_X1 U13770 ( .A1(n3421), .A2(n3383), .ZN(\mult_20/ab[27][8] ) );
  NOR2_X1 U13771 ( .A1(n3418), .A2(n3383), .ZN(\mult_20/ab[27][7] ) );
  NOR2_X1 U13772 ( .A1(n3415), .A2(n3383), .ZN(\mult_20/ab[27][6] ) );
  NOR2_X1 U13773 ( .A1(n3412), .A2(n3383), .ZN(\mult_20/ab[27][5] ) );
  NOR2_X1 U13774 ( .A1(n3223), .A2(n3197), .ZN(\mult_19/ab[27][4] ) );
  NOR2_X1 U13775 ( .A1(n3238), .A2(n3197), .ZN(\mult_19/ab[27][9] ) );
  NOR2_X1 U13776 ( .A1(n3235), .A2(n3197), .ZN(\mult_19/ab[27][8] ) );
  NOR2_X1 U13777 ( .A1(n3232), .A2(n3197), .ZN(\mult_19/ab[27][7] ) );
  NOR2_X1 U13778 ( .A1(n3229), .A2(n3197), .ZN(\mult_19/ab[27][6] ) );
  NOR2_X1 U13779 ( .A1(n3406), .A2(n3383), .ZN(\mult_20/ab[27][3] ) );
  NOR2_X1 U13780 ( .A1(n3424), .A2(n3386), .ZN(\mult_20/ab[28][9] ) );
  NOR2_X1 U13781 ( .A1(n3421), .A2(n3386), .ZN(\mult_20/ab[28][8] ) );
  NOR2_X1 U13782 ( .A1(n3418), .A2(n3386), .ZN(\mult_20/ab[28][7] ) );
  NOR2_X1 U13783 ( .A1(n3415), .A2(n3386), .ZN(\mult_20/ab[28][6] ) );
  NOR2_X1 U13784 ( .A1(n3412), .A2(n3386), .ZN(\mult_20/ab[28][5] ) );
  NOR2_X1 U13785 ( .A1(n3223), .A2(n3200), .ZN(\mult_19/ab[28][4] ) );
  NOR2_X1 U13786 ( .A1(n3238), .A2(n3200), .ZN(\mult_19/ab[28][9] ) );
  NOR2_X1 U13787 ( .A1(n3235), .A2(n3200), .ZN(\mult_19/ab[28][8] ) );
  NOR2_X1 U13788 ( .A1(n3232), .A2(n3200), .ZN(\mult_19/ab[28][7] ) );
  NOR2_X1 U13789 ( .A1(n3229), .A2(n3200), .ZN(\mult_19/ab[28][6] ) );
  NOR2_X1 U13790 ( .A1(n3226), .A2(n3200), .ZN(\mult_19/ab[28][5] ) );
  NOR2_X1 U13791 ( .A1(n3409), .A2(n3386), .ZN(\mult_20/ab[28][4] ) );
  NOR2_X1 U13792 ( .A1(n3406), .A2(n3386), .ZN(\mult_20/ab[28][3] ) );
  NOR2_X1 U13793 ( .A1(n3420), .A2(n3389), .ZN(\mult_20/ab[29][8] ) );
  NOR2_X1 U13794 ( .A1(n3417), .A2(n3389), .ZN(\mult_20/ab[29][7] ) );
  NOR2_X1 U13795 ( .A1(n3414), .A2(n3389), .ZN(\mult_20/ab[29][6] ) );
  NOR2_X1 U13796 ( .A1(n3411), .A2(n3389), .ZN(\mult_20/ab[29][5] ) );
  NOR2_X1 U13797 ( .A1(n3222), .A2(n3203), .ZN(\mult_19/ab[29][4] ) );
  NOR2_X1 U13798 ( .A1(n3234), .A2(n3203), .ZN(\mult_19/ab[29][8] ) );
  NOR2_X1 U13799 ( .A1(n3231), .A2(n3203), .ZN(\mult_19/ab[29][7] ) );
  NOR2_X1 U13800 ( .A1(n3228), .A2(n3203), .ZN(\mult_19/ab[29][6] ) );
  NOR2_X1 U13801 ( .A1(n3225), .A2(n3203), .ZN(\mult_19/ab[29][5] ) );
  NOR2_X1 U13802 ( .A1(n3405), .A2(n3389), .ZN(\mult_20/ab[29][3] ) );
  NOR2_X1 U13803 ( .A1(n3417), .A2(n3392), .ZN(\mult_20/ab[30][7] ) );
  NOR2_X1 U13804 ( .A1(n3414), .A2(n3392), .ZN(\mult_20/ab[30][6] ) );
  NOR2_X1 U13805 ( .A1(n3231), .A2(n3206), .ZN(\mult_19/ab[30][7] ) );
  NOR2_X1 U13806 ( .A1(n3228), .A2(n3206), .ZN(\mult_19/ab[30][6] ) );
  NOR2_X1 U13807 ( .A1(n3225), .A2(n3206), .ZN(\mult_19/ab[30][5] ) );
  NOR2_X1 U13808 ( .A1(n3408), .A2(n3389), .ZN(\mult_20/ab[29][4] ) );
  NOR2_X1 U13809 ( .A1(n3423), .A2(n3389), .ZN(\mult_20/ab[29][9] ) );
  NOR2_X1 U13810 ( .A1(n3237), .A2(n3203), .ZN(\mult_19/ab[29][9] ) );
  NOR2_X1 U13811 ( .A1(n3405), .A2(n3392), .ZN(\mult_20/ab[30][3] ) );
  NOR2_X1 U13812 ( .A1(n3420), .A2(n3392), .ZN(\mult_20/ab[30][8] ) );
  NOR2_X1 U13813 ( .A1(n3423), .A2(n3392), .ZN(\mult_20/ab[30][9] ) );
  NOR2_X1 U13814 ( .A1(n3234), .A2(n3206), .ZN(\mult_19/ab[30][8] ) );
  NOR2_X1 U13815 ( .A1(n3237), .A2(n3206), .ZN(\mult_19/ab[30][9] ) );
  NOR2_X1 U13816 ( .A1(n3222), .A2(n3206), .ZN(\mult_19/ab[30][4] ) );
  NOR2_X1 U13817 ( .A1(n3408), .A2(n3392), .ZN(\mult_20/ab[30][4] ) );
  NOR2_X1 U13818 ( .A1(n3456), .A2(n3310), .ZN(\mult_20/ab[3][20] ) );
  NOR2_X1 U13819 ( .A1(n3450), .A2(n3309), .ZN(\mult_20/ab[3][18] ) );
  NOR2_X1 U13820 ( .A1(n3444), .A2(n3309), .ZN(\mult_20/ab[3][16] ) );
  NOR2_X1 U13821 ( .A1(n3438), .A2(n3309), .ZN(\mult_20/ab[3][14] ) );
  NOR2_X1 U13822 ( .A1(n3432), .A2(n3309), .ZN(\mult_20/ab[3][12] ) );
  NOR2_X1 U13823 ( .A1(n3426), .A2(n3309), .ZN(\mult_20/ab[3][10] ) );
  NOR2_X1 U13824 ( .A1(n3276), .A2(n3124), .ZN(\mult_19/ab[3][22] ) );
  NOR2_X1 U13825 ( .A1(n3450), .A2(n3312), .ZN(\mult_20/ab[4][18] ) );
  NOR2_X1 U13826 ( .A1(n3444), .A2(n3312), .ZN(\mult_20/ab[4][16] ) );
  NOR2_X1 U13827 ( .A1(n3438), .A2(n3312), .ZN(\mult_20/ab[4][14] ) );
  NOR2_X1 U13828 ( .A1(n3432), .A2(n3312), .ZN(\mult_20/ab[4][12] ) );
  NOR2_X1 U13829 ( .A1(n3426), .A2(n3312), .ZN(\mult_20/ab[4][10] ) );
  NOR2_X1 U13830 ( .A1(n3270), .A2(n3127), .ZN(\mult_19/ab[4][20] ) );
  NOR2_X1 U13831 ( .A1(n3267), .A2(n3126), .ZN(\mult_19/ab[4][19] ) );
  NOR2_X1 U13832 ( .A1(n3264), .A2(n3126), .ZN(\mult_19/ab[4][18] ) );
  NOR2_X1 U13833 ( .A1(n3261), .A2(n3126), .ZN(\mult_19/ab[4][17] ) );
  NOR2_X1 U13834 ( .A1(n3258), .A2(n3126), .ZN(\mult_19/ab[4][16] ) );
  NOR2_X1 U13835 ( .A1(n3255), .A2(n3126), .ZN(\mult_19/ab[4][15] ) );
  NOR2_X1 U13836 ( .A1(n3252), .A2(n3126), .ZN(\mult_19/ab[4][14] ) );
  NOR2_X1 U13837 ( .A1(n3249), .A2(n3126), .ZN(\mult_19/ab[4][13] ) );
  NOR2_X1 U13838 ( .A1(n3246), .A2(n3126), .ZN(\mult_19/ab[4][12] ) );
  NOR2_X1 U13839 ( .A1(n3243), .A2(n3126), .ZN(\mult_19/ab[4][11] ) );
  NOR2_X1 U13840 ( .A1(n3240), .A2(n3126), .ZN(\mult_19/ab[4][10] ) );
  NOR2_X1 U13841 ( .A1(n3456), .A2(n3316), .ZN(\mult_20/ab[5][20] ) );
  NOR2_X1 U13842 ( .A1(n3450), .A2(n3315), .ZN(\mult_20/ab[5][18] ) );
  NOR2_X1 U13843 ( .A1(n3444), .A2(n3315), .ZN(\mult_20/ab[5][16] ) );
  NOR2_X1 U13844 ( .A1(n3438), .A2(n3315), .ZN(\mult_20/ab[5][14] ) );
  NOR2_X1 U13845 ( .A1(n3432), .A2(n3315), .ZN(\mult_20/ab[5][12] ) );
  NOR2_X1 U13846 ( .A1(n3426), .A2(n3315), .ZN(\mult_20/ab[5][10] ) );
  NOR2_X1 U13847 ( .A1(n3273), .A2(n3130), .ZN(\mult_19/ab[5][21] ) );
  NOR2_X1 U13848 ( .A1(n3270), .A2(n3130), .ZN(\mult_19/ab[5][20] ) );
  NOR2_X1 U13849 ( .A1(n3450), .A2(n3318), .ZN(\mult_20/ab[6][18] ) );
  NOR2_X1 U13850 ( .A1(n3444), .A2(n3318), .ZN(\mult_20/ab[6][16] ) );
  NOR2_X1 U13851 ( .A1(n3438), .A2(n3318), .ZN(\mult_20/ab[6][14] ) );
  NOR2_X1 U13852 ( .A1(n3432), .A2(n3318), .ZN(\mult_20/ab[6][12] ) );
  NOR2_X1 U13853 ( .A1(n3426), .A2(n3318), .ZN(\mult_20/ab[6][10] ) );
  NOR2_X1 U13854 ( .A1(n3264), .A2(n3132), .ZN(\mult_19/ab[6][18] ) );
  NOR2_X1 U13855 ( .A1(n3261), .A2(n3132), .ZN(\mult_19/ab[6][17] ) );
  NOR2_X1 U13856 ( .A1(n3258), .A2(n3132), .ZN(\mult_19/ab[6][16] ) );
  NOR2_X1 U13857 ( .A1(n3255), .A2(n3132), .ZN(\mult_19/ab[6][15] ) );
  NOR2_X1 U13858 ( .A1(n3252), .A2(n3132), .ZN(\mult_19/ab[6][14] ) );
  NOR2_X1 U13859 ( .A1(n3249), .A2(n3132), .ZN(\mult_19/ab[6][13] ) );
  NOR2_X1 U13860 ( .A1(n3246), .A2(n3132), .ZN(\mult_19/ab[6][12] ) );
  NOR2_X1 U13861 ( .A1(n3243), .A2(n3132), .ZN(\mult_19/ab[6][11] ) );
  NOR2_X1 U13862 ( .A1(n3240), .A2(n3132), .ZN(\mult_19/ab[6][10] ) );
  NOR2_X1 U13863 ( .A1(n3444), .A2(n3321), .ZN(\mult_20/ab[7][16] ) );
  NOR2_X1 U13864 ( .A1(n3438), .A2(n3321), .ZN(\mult_20/ab[7][14] ) );
  NOR2_X1 U13865 ( .A1(n3432), .A2(n3321), .ZN(\mult_20/ab[7][12] ) );
  NOR2_X1 U13866 ( .A1(n3426), .A2(n3321), .ZN(\mult_20/ab[7][10] ) );
  NOR2_X1 U13867 ( .A1(n3264), .A2(n3135), .ZN(\mult_19/ab[7][18] ) );
  NOR2_X1 U13868 ( .A1(n3444), .A2(n3324), .ZN(\mult_20/ab[8][16] ) );
  NOR2_X1 U13869 ( .A1(n3438), .A2(n3324), .ZN(\mult_20/ab[8][14] ) );
  NOR2_X1 U13870 ( .A1(n3432), .A2(n3324), .ZN(\mult_20/ab[8][12] ) );
  NOR2_X1 U13871 ( .A1(n3426), .A2(n3324), .ZN(\mult_20/ab[8][10] ) );
  NOR2_X1 U13872 ( .A1(n3258), .A2(n3138), .ZN(\mult_19/ab[8][16] ) );
  NOR2_X1 U13873 ( .A1(n3255), .A2(n3138), .ZN(\mult_19/ab[8][15] ) );
  NOR2_X1 U13874 ( .A1(n3252), .A2(n3138), .ZN(\mult_19/ab[8][14] ) );
  NOR2_X1 U13875 ( .A1(n3249), .A2(n3138), .ZN(\mult_19/ab[8][13] ) );
  NOR2_X1 U13876 ( .A1(n3246), .A2(n3138), .ZN(\mult_19/ab[8][12] ) );
  NOR2_X1 U13877 ( .A1(n3243), .A2(n3138), .ZN(\mult_19/ab[8][11] ) );
  NOR2_X1 U13878 ( .A1(n3240), .A2(n3138), .ZN(\mult_19/ab[8][10] ) );
  NOR2_X1 U13879 ( .A1(n3444), .A2(n3327), .ZN(\mult_20/ab[9][16] ) );
  NOR2_X1 U13880 ( .A1(n3438), .A2(n3327), .ZN(\mult_20/ab[9][14] ) );
  NOR2_X1 U13881 ( .A1(n3432), .A2(n3327), .ZN(\mult_20/ab[9][12] ) );
  NOR2_X1 U13882 ( .A1(n3426), .A2(n3327), .ZN(\mult_20/ab[9][10] ) );
  NOR2_X1 U13883 ( .A1(n3261), .A2(n3141), .ZN(\mult_19/ab[9][17] ) );
  NOR2_X1 U13884 ( .A1(n3258), .A2(n3141), .ZN(\mult_19/ab[9][16] ) );
  NOR2_X1 U13885 ( .A1(n3452), .A2(n3330), .ZN(\mult_20/ab[10][18] ) );
  NOR2_X1 U13886 ( .A1(n3446), .A2(n3330), .ZN(\mult_20/ab[10][16] ) );
  NOR2_X1 U13887 ( .A1(n3440), .A2(n3330), .ZN(\mult_20/ab[10][14] ) );
  NOR2_X1 U13888 ( .A1(n3434), .A2(n3330), .ZN(\mult_20/ab[10][12] ) );
  NOR2_X1 U13889 ( .A1(n3428), .A2(n3330), .ZN(\mult_20/ab[10][10] ) );
  NOR2_X1 U13890 ( .A1(n3254), .A2(n3144), .ZN(\mult_19/ab[10][14] ) );
  NOR2_X1 U13891 ( .A1(n3251), .A2(n3144), .ZN(\mult_19/ab[10][13] ) );
  NOR2_X1 U13892 ( .A1(n3248), .A2(n3144), .ZN(\mult_19/ab[10][12] ) );
  NOR2_X1 U13893 ( .A1(n3245), .A2(n3144), .ZN(\mult_19/ab[10][11] ) );
  NOR2_X1 U13894 ( .A1(n3242), .A2(n3144), .ZN(\mult_19/ab[10][10] ) );
  NOR2_X1 U13895 ( .A1(n3458), .A2(n3334), .ZN(\mult_20/ab[11][20] ) );
  NOR2_X1 U13896 ( .A1(n3452), .A2(n3333), .ZN(\mult_20/ab[11][18] ) );
  NOR2_X1 U13897 ( .A1(n3446), .A2(n3333), .ZN(\mult_20/ab[11][16] ) );
  NOR2_X1 U13898 ( .A1(n3440), .A2(n3333), .ZN(\mult_20/ab[11][14] ) );
  NOR2_X1 U13899 ( .A1(n3434), .A2(n3333), .ZN(\mult_20/ab[11][12] ) );
  NOR2_X1 U13900 ( .A1(n3428), .A2(n3333), .ZN(\mult_20/ab[11][10] ) );
  NOR2_X1 U13901 ( .A1(n3275), .A2(n3148), .ZN(\mult_19/ab[11][21] ) );
  NOR2_X1 U13902 ( .A1(n3269), .A2(n3147), .ZN(\mult_19/ab[11][19] ) );
  NOR2_X1 U13903 ( .A1(n3266), .A2(n3147), .ZN(\mult_19/ab[11][18] ) );
  NOR2_X1 U13904 ( .A1(n3263), .A2(n3147), .ZN(\mult_19/ab[11][17] ) );
  NOR2_X1 U13905 ( .A1(n3260), .A2(n3147), .ZN(\mult_19/ab[11][16] ) );
  NOR2_X1 U13906 ( .A1(n3257), .A2(n3147), .ZN(\mult_19/ab[11][15] ) );
  NOR2_X1 U13907 ( .A1(n3254), .A2(n3147), .ZN(\mult_19/ab[11][14] ) );
  NOR2_X1 U13908 ( .A1(n3452), .A2(n3336), .ZN(\mult_20/ab[12][18] ) );
  NOR2_X1 U13909 ( .A1(n3446), .A2(n3336), .ZN(\mult_20/ab[12][16] ) );
  NOR2_X1 U13910 ( .A1(n3440), .A2(n3336), .ZN(\mult_20/ab[12][14] ) );
  NOR2_X1 U13911 ( .A1(n3434), .A2(n3336), .ZN(\mult_20/ab[12][12] ) );
  NOR2_X1 U13912 ( .A1(n3428), .A2(n3336), .ZN(\mult_20/ab[12][10] ) );
  NOR2_X1 U13913 ( .A1(n3269), .A2(n3150), .ZN(\mult_19/ab[12][19] ) );
  NOR2_X1 U13914 ( .A1(n3248), .A2(n3150), .ZN(\mult_19/ab[12][12] ) );
  NOR2_X1 U13915 ( .A1(n3245), .A2(n3150), .ZN(\mult_19/ab[12][11] ) );
  NOR2_X1 U13916 ( .A1(n3242), .A2(n3150), .ZN(\mult_19/ab[12][10] ) );
  NOR2_X1 U13917 ( .A1(n3452), .A2(n3339), .ZN(\mult_20/ab[13][18] ) );
  NOR2_X1 U13918 ( .A1(n3434), .A2(n3339), .ZN(\mult_20/ab[13][12] ) );
  NOR2_X1 U13919 ( .A1(n3428), .A2(n3339), .ZN(\mult_20/ab[13][10] ) );
  NOR2_X1 U13920 ( .A1(n3254), .A2(n3153), .ZN(\mult_19/ab[13][14] ) );
  NOR2_X1 U13921 ( .A1(n3251), .A2(n3153), .ZN(\mult_19/ab[13][13] ) );
  NOR2_X1 U13922 ( .A1(n3248), .A2(n3153), .ZN(\mult_19/ab[13][12] ) );
  NOR2_X1 U13923 ( .A1(n3446), .A2(n3342), .ZN(\mult_20/ab[14][16] ) );
  NOR2_X1 U13924 ( .A1(n3440), .A2(n3342), .ZN(\mult_20/ab[14][14] ) );
  NOR2_X1 U13925 ( .A1(n3434), .A2(n3342), .ZN(\mult_20/ab[14][12] ) );
  NOR2_X1 U13926 ( .A1(n3428), .A2(n3342), .ZN(\mult_20/ab[14][10] ) );
  NOR2_X1 U13927 ( .A1(n3263), .A2(n3156), .ZN(\mult_19/ab[14][17] ) );
  NOR2_X1 U13928 ( .A1(n3242), .A2(n3156), .ZN(\mult_19/ab[14][10] ) );
  NOR2_X1 U13929 ( .A1(n3446), .A2(n3345), .ZN(\mult_20/ab[15][16] ) );
  NOR2_X1 U13930 ( .A1(n3440), .A2(n3345), .ZN(\mult_20/ab[15][14] ) );
  NOR2_X1 U13931 ( .A1(n3434), .A2(n3345), .ZN(\mult_20/ab[15][12] ) );
  NOR2_X1 U13932 ( .A1(n3428), .A2(n3345), .ZN(\mult_20/ab[15][10] ) );
  NOR2_X1 U13933 ( .A1(n3263), .A2(n3159), .ZN(\mult_19/ab[15][17] ) );
  NOR2_X1 U13934 ( .A1(n3257), .A2(n3159), .ZN(\mult_19/ab[15][15] ) );
  NOR2_X1 U13935 ( .A1(n3254), .A2(n3159), .ZN(\mult_19/ab[15][14] ) );
  NOR2_X1 U13936 ( .A1(n3251), .A2(n3159), .ZN(\mult_19/ab[15][13] ) );
  NOR2_X1 U13937 ( .A1(n3248), .A2(n3159), .ZN(\mult_19/ab[15][12] ) );
  NOR2_X1 U13938 ( .A1(n3245), .A2(n3159), .ZN(\mult_19/ab[15][11] ) );
  NOR2_X1 U13939 ( .A1(n3242), .A2(n3159), .ZN(\mult_19/ab[15][10] ) );
  NOR2_X1 U13940 ( .A1(n3440), .A2(n3348), .ZN(\mult_20/ab[16][14] ) );
  NOR2_X1 U13941 ( .A1(n3434), .A2(n3348), .ZN(\mult_20/ab[16][12] ) );
  NOR2_X1 U13942 ( .A1(n3428), .A2(n3348), .ZN(\mult_20/ab[16][10] ) );
  NOR2_X1 U13943 ( .A1(n3257), .A2(n3162), .ZN(\mult_19/ab[16][15] ) );
  NOR2_X1 U13944 ( .A1(n3439), .A2(n3351), .ZN(\mult_20/ab[17][14] ) );
  NOR2_X1 U13945 ( .A1(n3433), .A2(n3351), .ZN(\mult_20/ab[17][12] ) );
  NOR2_X1 U13946 ( .A1(n3427), .A2(n3351), .ZN(\mult_20/ab[17][10] ) );
  NOR2_X1 U13947 ( .A1(n3256), .A2(n3165), .ZN(\mult_19/ab[17][15] ) );
  NOR2_X1 U13948 ( .A1(n3250), .A2(n3165), .ZN(\mult_19/ab[17][13] ) );
  NOR2_X1 U13949 ( .A1(n3247), .A2(n3165), .ZN(\mult_19/ab[17][12] ) );
  NOR2_X1 U13950 ( .A1(n3244), .A2(n3165), .ZN(\mult_19/ab[17][11] ) );
  NOR2_X1 U13951 ( .A1(n3241), .A2(n3165), .ZN(\mult_19/ab[17][10] ) );
  NOR2_X1 U13952 ( .A1(n3433), .A2(n3354), .ZN(\mult_20/ab[18][12] ) );
  NOR2_X1 U13953 ( .A1(n3427), .A2(n3354), .ZN(\mult_20/ab[18][10] ) );
  NOR2_X1 U13954 ( .A1(n3250), .A2(n3168), .ZN(\mult_19/ab[18][13] ) );
  NOR2_X1 U13955 ( .A1(n3433), .A2(n3357), .ZN(\mult_20/ab[19][12] ) );
  NOR2_X1 U13956 ( .A1(n3427), .A2(n3357), .ZN(\mult_20/ab[19][10] ) );
  NOR2_X1 U13957 ( .A1(n3250), .A2(n3171), .ZN(\mult_19/ab[19][13] ) );
  NOR2_X1 U13958 ( .A1(n3244), .A2(n3171), .ZN(\mult_19/ab[19][11] ) );
  NOR2_X1 U13959 ( .A1(n3241), .A2(n3171), .ZN(\mult_19/ab[19][10] ) );
  NOR2_X1 U13960 ( .A1(n3427), .A2(n3360), .ZN(\mult_20/ab[20][10] ) );
  NOR2_X1 U13961 ( .A1(n3244), .A2(n3174), .ZN(\mult_19/ab[20][11] ) );
  NOR2_X1 U13962 ( .A1(n3427), .A2(n3363), .ZN(\mult_20/ab[21][10] ) );
  NOR2_X1 U13963 ( .A1(n3244), .A2(n3177), .ZN(\mult_19/ab[21][11] ) );
  NOR2_X1 U13964 ( .A1(n3420), .A2(n3311), .ZN(\mult_20/ab[3][8] ) );
  NOR2_X1 U13965 ( .A1(n3414), .A2(n3311), .ZN(\mult_20/ab[3][6] ) );
  NOR2_X1 U13966 ( .A1(n3216), .A2(n3124), .ZN(\mult_19/ab[3][2] ) );
  NOR2_X1 U13967 ( .A1(n3213), .A2(n3123), .ZN(\mult_19/ab[3][1] ) );
  NOR2_X1 U13968 ( .A1(n3408), .A2(n3311), .ZN(\mult_20/ab[3][4] ) );
  NOR2_X1 U13969 ( .A1(n3402), .A2(n3310), .ZN(\mult_20/ab[3][2] ) );
  NOR2_X1 U13970 ( .A1(n3399), .A2(n3309), .ZN(\mult_20/ab[3][1] ) );
  NOR2_X1 U13971 ( .A1(n3420), .A2(n3314), .ZN(\mult_20/ab[4][8] ) );
  NOR2_X1 U13972 ( .A1(n3414), .A2(n3314), .ZN(\mult_20/ab[4][6] ) );
  NOR2_X1 U13973 ( .A1(n3222), .A2(n3128), .ZN(\mult_19/ab[4][4] ) );
  NOR2_X1 U13974 ( .A1(n3219), .A2(n3128), .ZN(\mult_19/ab[4][3] ) );
  NOR2_X1 U13975 ( .A1(n3216), .A2(n3127), .ZN(\mult_19/ab[4][2] ) );
  NOR2_X1 U13976 ( .A1(n3213), .A2(n3126), .ZN(\mult_19/ab[4][1] ) );
  NOR2_X1 U13977 ( .A1(n3237), .A2(n3128), .ZN(\mult_19/ab[4][9] ) );
  NOR2_X1 U13978 ( .A1(n3234), .A2(n3128), .ZN(\mult_19/ab[4][8] ) );
  NOR2_X1 U13979 ( .A1(n3231), .A2(n3128), .ZN(\mult_19/ab[4][7] ) );
  NOR2_X1 U13980 ( .A1(n3228), .A2(n3128), .ZN(\mult_19/ab[4][6] ) );
  NOR2_X1 U13981 ( .A1(n3225), .A2(n3128), .ZN(\mult_19/ab[4][5] ) );
  NOR2_X1 U13982 ( .A1(n3408), .A2(n3314), .ZN(\mult_20/ab[4][4] ) );
  NOR2_X1 U13983 ( .A1(n3402), .A2(n3313), .ZN(\mult_20/ab[4][2] ) );
  NOR2_X1 U13984 ( .A1(n3399), .A2(n3312), .ZN(\mult_20/ab[4][1] ) );
  NOR2_X1 U13985 ( .A1(n3420), .A2(n3317), .ZN(\mult_20/ab[5][8] ) );
  NOR2_X1 U13986 ( .A1(n3414), .A2(n3317), .ZN(\mult_20/ab[5][6] ) );
  NOR2_X1 U13987 ( .A1(n3216), .A2(n3130), .ZN(\mult_19/ab[5][2] ) );
  NOR2_X1 U13988 ( .A1(n3213), .A2(n3129), .ZN(\mult_19/ab[5][1] ) );
  NOR2_X1 U13989 ( .A1(n3408), .A2(n3317), .ZN(\mult_20/ab[5][4] ) );
  NOR2_X1 U13990 ( .A1(n3402), .A2(n3316), .ZN(\mult_20/ab[5][2] ) );
  NOR2_X1 U13991 ( .A1(n3399), .A2(n3315), .ZN(\mult_20/ab[5][1] ) );
  NOR2_X1 U13992 ( .A1(n3420), .A2(n3320), .ZN(\mult_20/ab[6][8] ) );
  NOR2_X1 U13993 ( .A1(n3414), .A2(n3320), .ZN(\mult_20/ab[6][6] ) );
  NOR2_X1 U13994 ( .A1(n3222), .A2(n3134), .ZN(\mult_19/ab[6][4] ) );
  NOR2_X1 U13995 ( .A1(n3219), .A2(n3134), .ZN(\mult_19/ab[6][3] ) );
  NOR2_X1 U13996 ( .A1(n3216), .A2(n3133), .ZN(\mult_19/ab[6][2] ) );
  NOR2_X1 U13997 ( .A1(n3213), .A2(n3132), .ZN(\mult_19/ab[6][1] ) );
  NOR2_X1 U13998 ( .A1(n3237), .A2(n3134), .ZN(\mult_19/ab[6][9] ) );
  NOR2_X1 U13999 ( .A1(n3234), .A2(n3134), .ZN(\mult_19/ab[6][8] ) );
  NOR2_X1 U14000 ( .A1(n3231), .A2(n3134), .ZN(\mult_19/ab[6][7] ) );
  NOR2_X1 U14001 ( .A1(n3228), .A2(n3134), .ZN(\mult_19/ab[6][6] ) );
  NOR2_X1 U14002 ( .A1(n3225), .A2(n3134), .ZN(\mult_19/ab[6][5] ) );
  NOR2_X1 U14003 ( .A1(n3408), .A2(n3320), .ZN(\mult_20/ab[6][4] ) );
  NOR2_X1 U14004 ( .A1(n3402), .A2(n3319), .ZN(\mult_20/ab[6][2] ) );
  NOR2_X1 U14005 ( .A1(n3399), .A2(n3318), .ZN(\mult_20/ab[6][1] ) );
  NOR2_X1 U14006 ( .A1(n3420), .A2(n3323), .ZN(\mult_20/ab[7][8] ) );
  NOR2_X1 U14007 ( .A1(n3414), .A2(n3323), .ZN(\mult_20/ab[7][6] ) );
  NOR2_X1 U14008 ( .A1(n3216), .A2(n3136), .ZN(\mult_19/ab[7][2] ) );
  NOR2_X1 U14009 ( .A1(n3213), .A2(n3135), .ZN(\mult_19/ab[7][1] ) );
  NOR2_X1 U14010 ( .A1(n3408), .A2(n3323), .ZN(\mult_20/ab[7][4] ) );
  NOR2_X1 U14011 ( .A1(n3402), .A2(n3322), .ZN(\mult_20/ab[7][2] ) );
  NOR2_X1 U14012 ( .A1(n3399), .A2(n3321), .ZN(\mult_20/ab[7][1] ) );
  NOR2_X1 U14013 ( .A1(n3420), .A2(n3326), .ZN(\mult_20/ab[8][8] ) );
  NOR2_X1 U14014 ( .A1(n3414), .A2(n3326), .ZN(\mult_20/ab[8][6] ) );
  NOR2_X1 U14015 ( .A1(n3222), .A2(n3140), .ZN(\mult_19/ab[8][4] ) );
  NOR2_X1 U14016 ( .A1(n3219), .A2(n3140), .ZN(\mult_19/ab[8][3] ) );
  NOR2_X1 U14017 ( .A1(n3216), .A2(n3139), .ZN(\mult_19/ab[8][2] ) );
  NOR2_X1 U14018 ( .A1(n3213), .A2(n3138), .ZN(\mult_19/ab[8][1] ) );
  NOR2_X1 U14019 ( .A1(n3237), .A2(n3140), .ZN(\mult_19/ab[8][9] ) );
  NOR2_X1 U14020 ( .A1(n3234), .A2(n3140), .ZN(\mult_19/ab[8][8] ) );
  NOR2_X1 U14021 ( .A1(n3231), .A2(n3140), .ZN(\mult_19/ab[8][7] ) );
  NOR2_X1 U14022 ( .A1(n3228), .A2(n3140), .ZN(\mult_19/ab[8][6] ) );
  NOR2_X1 U14023 ( .A1(n3225), .A2(n3140), .ZN(\mult_19/ab[8][5] ) );
  NOR2_X1 U14024 ( .A1(n3408), .A2(n3326), .ZN(\mult_20/ab[8][4] ) );
  NOR2_X1 U14025 ( .A1(n3402), .A2(n3325), .ZN(\mult_20/ab[8][2] ) );
  NOR2_X1 U14026 ( .A1(n3399), .A2(n3324), .ZN(\mult_20/ab[8][1] ) );
  NOR2_X1 U14027 ( .A1(n3420), .A2(n3329), .ZN(\mult_20/ab[9][8] ) );
  NOR2_X1 U14028 ( .A1(n3414), .A2(n3329), .ZN(\mult_20/ab[9][6] ) );
  NOR2_X1 U14029 ( .A1(n3216), .A2(n3142), .ZN(\mult_19/ab[9][2] ) );
  NOR2_X1 U14030 ( .A1(n3213), .A2(n3141), .ZN(\mult_19/ab[9][1] ) );
  NOR2_X1 U14031 ( .A1(n3408), .A2(n3329), .ZN(\mult_20/ab[9][4] ) );
  NOR2_X1 U14032 ( .A1(n3402), .A2(n3328), .ZN(\mult_20/ab[9][2] ) );
  NOR2_X1 U14033 ( .A1(n3399), .A2(n3327), .ZN(\mult_20/ab[9][1] ) );
  NOR2_X1 U14034 ( .A1(n3422), .A2(n3332), .ZN(\mult_20/ab[10][8] ) );
  NOR2_X1 U14035 ( .A1(n3416), .A2(n3332), .ZN(\mult_20/ab[10][6] ) );
  NOR2_X1 U14036 ( .A1(n3224), .A2(n3146), .ZN(\mult_19/ab[10][4] ) );
  NOR2_X1 U14037 ( .A1(n3221), .A2(n3146), .ZN(\mult_19/ab[10][3] ) );
  NOR2_X1 U14038 ( .A1(n3218), .A2(n3145), .ZN(\mult_19/ab[10][2] ) );
  NOR2_X1 U14039 ( .A1(n3215), .A2(n3144), .ZN(\mult_19/ab[10][1] ) );
  NOR2_X1 U14040 ( .A1(n3239), .A2(n3146), .ZN(\mult_19/ab[10][9] ) );
  NOR2_X1 U14041 ( .A1(n3236), .A2(n3146), .ZN(\mult_19/ab[10][8] ) );
  NOR2_X1 U14042 ( .A1(n3233), .A2(n3146), .ZN(\mult_19/ab[10][7] ) );
  NOR2_X1 U14043 ( .A1(n3230), .A2(n3146), .ZN(\mult_19/ab[10][6] ) );
  NOR2_X1 U14044 ( .A1(n3227), .A2(n3146), .ZN(\mult_19/ab[10][5] ) );
  NOR2_X1 U14045 ( .A1(n3410), .A2(n3332), .ZN(\mult_20/ab[10][4] ) );
  NOR2_X1 U14046 ( .A1(n3404), .A2(n3331), .ZN(\mult_20/ab[10][2] ) );
  NOR2_X1 U14047 ( .A1(n3401), .A2(n3330), .ZN(\mult_20/ab[10][1] ) );
  NOR2_X1 U14048 ( .A1(n3422), .A2(n3335), .ZN(\mult_20/ab[11][8] ) );
  NOR2_X1 U14049 ( .A1(n3416), .A2(n3335), .ZN(\mult_20/ab[11][6] ) );
  NOR2_X1 U14050 ( .A1(n3218), .A2(n3148), .ZN(\mult_19/ab[11][2] ) );
  NOR2_X1 U14051 ( .A1(n3215), .A2(n3147), .ZN(\mult_19/ab[11][1] ) );
  NOR2_X1 U14052 ( .A1(n3410), .A2(n3335), .ZN(\mult_20/ab[11][4] ) );
  NOR2_X1 U14053 ( .A1(n3404), .A2(n3334), .ZN(\mult_20/ab[11][2] ) );
  NOR2_X1 U14054 ( .A1(n3401), .A2(n3333), .ZN(\mult_20/ab[11][1] ) );
  NOR2_X1 U14055 ( .A1(n3422), .A2(n3338), .ZN(\mult_20/ab[12][8] ) );
  NOR2_X1 U14056 ( .A1(n3416), .A2(n3338), .ZN(\mult_20/ab[12][6] ) );
  NOR2_X1 U14057 ( .A1(n3224), .A2(n3152), .ZN(\mult_19/ab[12][4] ) );
  NOR2_X1 U14058 ( .A1(n3221), .A2(n3152), .ZN(\mult_19/ab[12][3] ) );
  NOR2_X1 U14059 ( .A1(n3218), .A2(n3151), .ZN(\mult_19/ab[12][2] ) );
  NOR2_X1 U14060 ( .A1(n3215), .A2(n3150), .ZN(\mult_19/ab[12][1] ) );
  NOR2_X1 U14061 ( .A1(n3239), .A2(n3152), .ZN(\mult_19/ab[12][9] ) );
  NOR2_X1 U14062 ( .A1(n3236), .A2(n3152), .ZN(\mult_19/ab[12][8] ) );
  NOR2_X1 U14063 ( .A1(n3233), .A2(n3152), .ZN(\mult_19/ab[12][7] ) );
  NOR2_X1 U14064 ( .A1(n3230), .A2(n3152), .ZN(\mult_19/ab[12][6] ) );
  NOR2_X1 U14065 ( .A1(n3227), .A2(n3152), .ZN(\mult_19/ab[12][5] ) );
  NOR2_X1 U14066 ( .A1(n3410), .A2(n3338), .ZN(\mult_20/ab[12][4] ) );
  NOR2_X1 U14067 ( .A1(n3404), .A2(n3337), .ZN(\mult_20/ab[12][2] ) );
  NOR2_X1 U14068 ( .A1(n3401), .A2(n3336), .ZN(\mult_20/ab[12][1] ) );
  NOR2_X1 U14069 ( .A1(n3422), .A2(n3341), .ZN(\mult_20/ab[13][8] ) );
  NOR2_X1 U14070 ( .A1(n3416), .A2(n3341), .ZN(\mult_20/ab[13][6] ) );
  NOR2_X1 U14071 ( .A1(n3218), .A2(n3154), .ZN(\mult_19/ab[13][2] ) );
  NOR2_X1 U14072 ( .A1(n3215), .A2(n3153), .ZN(\mult_19/ab[13][1] ) );
  NOR2_X1 U14073 ( .A1(n3410), .A2(n3341), .ZN(\mult_20/ab[13][4] ) );
  NOR2_X1 U14074 ( .A1(n3404), .A2(n3340), .ZN(\mult_20/ab[13][2] ) );
  NOR2_X1 U14075 ( .A1(n3401), .A2(n3339), .ZN(\mult_20/ab[13][1] ) );
  NOR2_X1 U14076 ( .A1(n3422), .A2(n3344), .ZN(\mult_20/ab[14][8] ) );
  NOR2_X1 U14077 ( .A1(n3416), .A2(n3344), .ZN(\mult_20/ab[14][6] ) );
  NOR2_X1 U14078 ( .A1(n3224), .A2(n3158), .ZN(\mult_19/ab[14][4] ) );
  NOR2_X1 U14079 ( .A1(n3221), .A2(n3158), .ZN(\mult_19/ab[14][3] ) );
  NOR2_X1 U14080 ( .A1(n3218), .A2(n3157), .ZN(\mult_19/ab[14][2] ) );
  NOR2_X1 U14081 ( .A1(n3215), .A2(n3156), .ZN(\mult_19/ab[14][1] ) );
  NOR2_X1 U14082 ( .A1(n3239), .A2(n3158), .ZN(\mult_19/ab[14][9] ) );
  NOR2_X1 U14083 ( .A1(n3236), .A2(n3158), .ZN(\mult_19/ab[14][8] ) );
  NOR2_X1 U14084 ( .A1(n3233), .A2(n3158), .ZN(\mult_19/ab[14][7] ) );
  NOR2_X1 U14085 ( .A1(n3230), .A2(n3158), .ZN(\mult_19/ab[14][6] ) );
  NOR2_X1 U14086 ( .A1(n3227), .A2(n3158), .ZN(\mult_19/ab[14][5] ) );
  NOR2_X1 U14087 ( .A1(n3410), .A2(n3344), .ZN(\mult_20/ab[14][4] ) );
  NOR2_X1 U14088 ( .A1(n3404), .A2(n3343), .ZN(\mult_20/ab[14][2] ) );
  NOR2_X1 U14089 ( .A1(n3401), .A2(n3342), .ZN(\mult_20/ab[14][1] ) );
  NOR2_X1 U14090 ( .A1(n3422), .A2(n3347), .ZN(\mult_20/ab[15][8] ) );
  NOR2_X1 U14091 ( .A1(n3416), .A2(n3347), .ZN(\mult_20/ab[15][6] ) );
  NOR2_X1 U14092 ( .A1(n3218), .A2(n3160), .ZN(\mult_19/ab[15][2] ) );
  NOR2_X1 U14093 ( .A1(n3215), .A2(n3159), .ZN(\mult_19/ab[15][1] ) );
  NOR2_X1 U14094 ( .A1(n3410), .A2(n3347), .ZN(\mult_20/ab[15][4] ) );
  NOR2_X1 U14095 ( .A1(n3404), .A2(n3346), .ZN(\mult_20/ab[15][2] ) );
  NOR2_X1 U14096 ( .A1(n3401), .A2(n3345), .ZN(\mult_20/ab[15][1] ) );
  NOR2_X1 U14097 ( .A1(n3422), .A2(n3350), .ZN(\mult_20/ab[16][8] ) );
  NOR2_X1 U14098 ( .A1(n3416), .A2(n3350), .ZN(\mult_20/ab[16][6] ) );
  NOR2_X1 U14099 ( .A1(n3224), .A2(n3164), .ZN(\mult_19/ab[16][4] ) );
  NOR2_X1 U14100 ( .A1(n3221), .A2(n3164), .ZN(\mult_19/ab[16][3] ) );
  NOR2_X1 U14101 ( .A1(n3218), .A2(n3163), .ZN(\mult_19/ab[16][2] ) );
  NOR2_X1 U14102 ( .A1(n3215), .A2(n3162), .ZN(\mult_19/ab[16][1] ) );
  NOR2_X1 U14103 ( .A1(n3236), .A2(n3164), .ZN(\mult_19/ab[16][8] ) );
  NOR2_X1 U14104 ( .A1(n3233), .A2(n3164), .ZN(\mult_19/ab[16][7] ) );
  NOR2_X1 U14105 ( .A1(n3230), .A2(n3164), .ZN(\mult_19/ab[16][6] ) );
  NOR2_X1 U14106 ( .A1(n3227), .A2(n3164), .ZN(\mult_19/ab[16][5] ) );
  NOR2_X1 U14107 ( .A1(n3410), .A2(n3350), .ZN(\mult_20/ab[16][4] ) );
  NOR2_X1 U14108 ( .A1(n3404), .A2(n3349), .ZN(\mult_20/ab[16][2] ) );
  NOR2_X1 U14109 ( .A1(n3401), .A2(n3348), .ZN(\mult_20/ab[16][1] ) );
  NOR2_X1 U14110 ( .A1(n3421), .A2(n3353), .ZN(\mult_20/ab[17][8] ) );
  NOR2_X1 U14111 ( .A1(n3415), .A2(n3353), .ZN(\mult_20/ab[17][6] ) );
  NOR2_X1 U14112 ( .A1(n3217), .A2(n3166), .ZN(\mult_19/ab[17][2] ) );
  NOR2_X1 U14113 ( .A1(n3215), .A2(n3165), .ZN(\mult_19/ab[17][1] ) );
  NOR2_X1 U14114 ( .A1(n3238), .A2(n3167), .ZN(\mult_19/ab[17][9] ) );
  NOR2_X1 U14115 ( .A1(n3235), .A2(n3167), .ZN(\mult_19/ab[17][8] ) );
  NOR2_X1 U14116 ( .A1(n3409), .A2(n3353), .ZN(\mult_20/ab[17][4] ) );
  NOR2_X1 U14117 ( .A1(n3403), .A2(n3352), .ZN(\mult_20/ab[17][2] ) );
  NOR2_X1 U14118 ( .A1(n3401), .A2(n3351), .ZN(\mult_20/ab[17][1] ) );
  NOR2_X1 U14119 ( .A1(n3421), .A2(n3356), .ZN(\mult_20/ab[18][8] ) );
  NOR2_X1 U14120 ( .A1(n3415), .A2(n3356), .ZN(\mult_20/ab[18][6] ) );
  NOR2_X1 U14121 ( .A1(n3223), .A2(n3170), .ZN(\mult_19/ab[18][4] ) );
  NOR2_X1 U14122 ( .A1(n3220), .A2(n3170), .ZN(\mult_19/ab[18][3] ) );
  NOR2_X1 U14123 ( .A1(n3217), .A2(n3169), .ZN(\mult_19/ab[18][2] ) );
  NOR2_X1 U14124 ( .A1(n3214), .A2(n3168), .ZN(\mult_19/ab[18][1] ) );
  NOR2_X1 U14125 ( .A1(n3229), .A2(n3170), .ZN(\mult_19/ab[18][6] ) );
  NOR2_X1 U14126 ( .A1(n3226), .A2(n3170), .ZN(\mult_19/ab[18][5] ) );
  NOR2_X1 U14127 ( .A1(n3409), .A2(n3356), .ZN(\mult_20/ab[18][4] ) );
  NOR2_X1 U14128 ( .A1(n3403), .A2(n3355), .ZN(\mult_20/ab[18][2] ) );
  NOR2_X1 U14129 ( .A1(n3400), .A2(n3354), .ZN(\mult_20/ab[18][1] ) );
  NOR2_X1 U14130 ( .A1(n3421), .A2(n3359), .ZN(\mult_20/ab[19][8] ) );
  NOR2_X1 U14131 ( .A1(n3415), .A2(n3359), .ZN(\mult_20/ab[19][6] ) );
  NOR2_X1 U14132 ( .A1(n3217), .A2(n3172), .ZN(\mult_19/ab[19][2] ) );
  NOR2_X1 U14133 ( .A1(n3214), .A2(n3171), .ZN(\mult_19/ab[19][1] ) );
  NOR2_X1 U14134 ( .A1(n3238), .A2(n3173), .ZN(\mult_19/ab[19][9] ) );
  NOR2_X1 U14135 ( .A1(n3235), .A2(n3173), .ZN(\mult_19/ab[19][8] ) );
  NOR2_X1 U14136 ( .A1(n3232), .A2(n3173), .ZN(\mult_19/ab[19][7] ) );
  NOR2_X1 U14137 ( .A1(n3229), .A2(n3173), .ZN(\mult_19/ab[19][6] ) );
  NOR2_X1 U14138 ( .A1(n3409), .A2(n3359), .ZN(\mult_20/ab[19][4] ) );
  NOR2_X1 U14139 ( .A1(n3403), .A2(n3358), .ZN(\mult_20/ab[19][2] ) );
  NOR2_X1 U14140 ( .A1(n3400), .A2(n3357), .ZN(\mult_20/ab[19][1] ) );
  NOR2_X1 U14141 ( .A1(n3421), .A2(n3362), .ZN(\mult_20/ab[20][8] ) );
  NOR2_X1 U14142 ( .A1(n3415), .A2(n3362), .ZN(\mult_20/ab[20][6] ) );
  NOR2_X1 U14143 ( .A1(n3223), .A2(n3176), .ZN(\mult_19/ab[20][4] ) );
  NOR2_X1 U14144 ( .A1(n3220), .A2(n3176), .ZN(\mult_19/ab[20][3] ) );
  NOR2_X1 U14145 ( .A1(n3217), .A2(n3175), .ZN(\mult_19/ab[20][2] ) );
  NOR2_X1 U14146 ( .A1(n3214), .A2(n3174), .ZN(\mult_19/ab[20][1] ) );
  NOR2_X1 U14147 ( .A1(n3409), .A2(n3362), .ZN(\mult_20/ab[20][4] ) );
  NOR2_X1 U14148 ( .A1(n3403), .A2(n3361), .ZN(\mult_20/ab[20][2] ) );
  NOR2_X1 U14149 ( .A1(n3400), .A2(n3360), .ZN(\mult_20/ab[20][1] ) );
  NOR2_X1 U14150 ( .A1(n3421), .A2(n3365), .ZN(\mult_20/ab[21][8] ) );
  NOR2_X1 U14151 ( .A1(n3415), .A2(n3365), .ZN(\mult_20/ab[21][6] ) );
  NOR2_X1 U14152 ( .A1(n3223), .A2(n3179), .ZN(\mult_19/ab[21][4] ) );
  NOR2_X1 U14153 ( .A1(n3217), .A2(n3178), .ZN(\mult_19/ab[21][2] ) );
  NOR2_X1 U14154 ( .A1(n3214), .A2(n3177), .ZN(\mult_19/ab[21][1] ) );
  NOR2_X1 U14155 ( .A1(n3238), .A2(n3179), .ZN(\mult_19/ab[21][9] ) );
  NOR2_X1 U14156 ( .A1(n3235), .A2(n3179), .ZN(\mult_19/ab[21][8] ) );
  NOR2_X1 U14157 ( .A1(n3232), .A2(n3179), .ZN(\mult_19/ab[21][7] ) );
  NOR2_X1 U14158 ( .A1(n3229), .A2(n3179), .ZN(\mult_19/ab[21][6] ) );
  NOR2_X1 U14159 ( .A1(n3226), .A2(n3179), .ZN(\mult_19/ab[21][5] ) );
  NOR2_X1 U14160 ( .A1(n3409), .A2(n3365), .ZN(\mult_20/ab[21][4] ) );
  NOR2_X1 U14161 ( .A1(n3403), .A2(n3364), .ZN(\mult_20/ab[21][2] ) );
  NOR2_X1 U14162 ( .A1(n3400), .A2(n3363), .ZN(\mult_20/ab[21][1] ) );
  NOR2_X1 U14163 ( .A1(n3421), .A2(n3368), .ZN(\mult_20/ab[22][8] ) );
  NOR2_X1 U14164 ( .A1(n3415), .A2(n3368), .ZN(\mult_20/ab[22][6] ) );
  NOR2_X1 U14165 ( .A1(n3217), .A2(n3181), .ZN(\mult_19/ab[22][2] ) );
  NOR2_X1 U14166 ( .A1(n3214), .A2(n3180), .ZN(\mult_19/ab[22][1] ) );
  NOR2_X1 U14167 ( .A1(n3238), .A2(n3182), .ZN(\mult_19/ab[22][9] ) );
  NOR2_X1 U14168 ( .A1(n3409), .A2(n3368), .ZN(\mult_20/ab[22][4] ) );
  NOR2_X1 U14169 ( .A1(n3403), .A2(n3367), .ZN(\mult_20/ab[22][2] ) );
  NOR2_X1 U14170 ( .A1(n3400), .A2(n3366), .ZN(\mult_20/ab[22][1] ) );
  NOR2_X1 U14171 ( .A1(n3421), .A2(n3371), .ZN(\mult_20/ab[23][8] ) );
  NOR2_X1 U14172 ( .A1(n3415), .A2(n3371), .ZN(\mult_20/ab[23][6] ) );
  NOR2_X1 U14173 ( .A1(n3223), .A2(n3185), .ZN(\mult_19/ab[23][4] ) );
  NOR2_X1 U14174 ( .A1(n3220), .A2(n3185), .ZN(\mult_19/ab[23][3] ) );
  NOR2_X1 U14175 ( .A1(n3217), .A2(n3184), .ZN(\mult_19/ab[23][2] ) );
  NOR2_X1 U14176 ( .A1(n3214), .A2(n3183), .ZN(\mult_19/ab[23][1] ) );
  NOR2_X1 U14177 ( .A1(n3238), .A2(n3185), .ZN(\mult_19/ab[23][9] ) );
  NOR2_X1 U14178 ( .A1(n3232), .A2(n3185), .ZN(\mult_19/ab[23][7] ) );
  NOR2_X1 U14179 ( .A1(n3229), .A2(n3185), .ZN(\mult_19/ab[23][6] ) );
  NOR2_X1 U14180 ( .A1(n3226), .A2(n3185), .ZN(\mult_19/ab[23][5] ) );
  NOR2_X1 U14181 ( .A1(n3409), .A2(n3371), .ZN(\mult_20/ab[23][4] ) );
  NOR2_X1 U14182 ( .A1(n3403), .A2(n3370), .ZN(\mult_20/ab[23][2] ) );
  NOR2_X1 U14183 ( .A1(n3400), .A2(n3369), .ZN(\mult_20/ab[23][1] ) );
  NOR2_X1 U14184 ( .A1(n3415), .A2(n3374), .ZN(\mult_20/ab[24][6] ) );
  NOR2_X1 U14185 ( .A1(n3217), .A2(n3187), .ZN(\mult_19/ab[24][2] ) );
  NOR2_X1 U14186 ( .A1(n3214), .A2(n3186), .ZN(\mult_19/ab[24][1] ) );
  NOR2_X1 U14187 ( .A1(n3232), .A2(n3188), .ZN(\mult_19/ab[24][7] ) );
  NOR2_X1 U14188 ( .A1(n3409), .A2(n3374), .ZN(\mult_20/ab[24][4] ) );
  NOR2_X1 U14189 ( .A1(n3403), .A2(n3373), .ZN(\mult_20/ab[24][2] ) );
  NOR2_X1 U14190 ( .A1(n3400), .A2(n3372), .ZN(\mult_20/ab[24][1] ) );
  NOR2_X1 U14191 ( .A1(n3415), .A2(n3377), .ZN(\mult_20/ab[25][6] ) );
  NOR2_X1 U14192 ( .A1(n3223), .A2(n3191), .ZN(\mult_19/ab[25][4] ) );
  NOR2_X1 U14193 ( .A1(n3220), .A2(n3191), .ZN(\mult_19/ab[25][3] ) );
  NOR2_X1 U14194 ( .A1(n3217), .A2(n3190), .ZN(\mult_19/ab[25][2] ) );
  NOR2_X1 U14195 ( .A1(n3214), .A2(n3189), .ZN(\mult_19/ab[25][1] ) );
  NOR2_X1 U14196 ( .A1(n3232), .A2(n3191), .ZN(\mult_19/ab[25][7] ) );
  NOR2_X1 U14197 ( .A1(n3226), .A2(n3191), .ZN(\mult_19/ab[25][5] ) );
  NOR2_X1 U14198 ( .A1(n3409), .A2(n3377), .ZN(\mult_20/ab[25][4] ) );
  NOR2_X1 U14199 ( .A1(n3403), .A2(n3376), .ZN(\mult_20/ab[25][2] ) );
  NOR2_X1 U14200 ( .A1(n3400), .A2(n3375), .ZN(\mult_20/ab[25][1] ) );
  NOR2_X1 U14201 ( .A1(n3217), .A2(n3193), .ZN(\mult_19/ab[26][2] ) );
  NOR2_X1 U14202 ( .A1(n3214), .A2(n3192), .ZN(\mult_19/ab[26][1] ) );
  NOR2_X1 U14203 ( .A1(n3226), .A2(n3194), .ZN(\mult_19/ab[26][5] ) );
  NOR2_X1 U14204 ( .A1(n3409), .A2(n3380), .ZN(\mult_20/ab[26][4] ) );
  NOR2_X1 U14205 ( .A1(n3403), .A2(n3379), .ZN(\mult_20/ab[26][2] ) );
  NOR2_X1 U14206 ( .A1(n3400), .A2(n3378), .ZN(\mult_20/ab[26][1] ) );
  NOR2_X1 U14207 ( .A1(n3220), .A2(n3197), .ZN(\mult_19/ab[27][3] ) );
  NOR2_X1 U14208 ( .A1(n3217), .A2(n3196), .ZN(\mult_19/ab[27][2] ) );
  NOR2_X1 U14209 ( .A1(n3214), .A2(n3195), .ZN(\mult_19/ab[27][1] ) );
  NOR2_X1 U14210 ( .A1(n3226), .A2(n3197), .ZN(\mult_19/ab[27][5] ) );
  NOR2_X1 U14211 ( .A1(n3409), .A2(n3383), .ZN(\mult_20/ab[27][4] ) );
  NOR2_X1 U14212 ( .A1(n3403), .A2(n3382), .ZN(\mult_20/ab[27][2] ) );
  NOR2_X1 U14213 ( .A1(n3400), .A2(n3381), .ZN(\mult_20/ab[27][1] ) );
  NOR2_X1 U14214 ( .A1(n3220), .A2(n3200), .ZN(\mult_19/ab[28][3] ) );
  NOR2_X1 U14215 ( .A1(n3217), .A2(n3199), .ZN(\mult_19/ab[28][2] ) );
  NOR2_X1 U14216 ( .A1(n3214), .A2(n3198), .ZN(\mult_19/ab[28][1] ) );
  NOR2_X1 U14217 ( .A1(n3403), .A2(n3385), .ZN(\mult_20/ab[28][2] ) );
  NOR2_X1 U14218 ( .A1(n3400), .A2(n3384), .ZN(\mult_20/ab[28][1] ) );
  NOR2_X1 U14219 ( .A1(n3219), .A2(n3203), .ZN(\mult_19/ab[29][3] ) );
  NOR2_X1 U14220 ( .A1(n3216), .A2(n3202), .ZN(\mult_19/ab[29][2] ) );
  NOR2_X1 U14221 ( .A1(n3214), .A2(n3201), .ZN(\mult_19/ab[29][1] ) );
  NOR2_X1 U14222 ( .A1(n3402), .A2(n3388), .ZN(\mult_20/ab[29][2] ) );
  NOR2_X1 U14223 ( .A1(n3400), .A2(n3387), .ZN(\mult_20/ab[29][1] ) );
  NOR2_X1 U14224 ( .A1(n3411), .A2(n3392), .ZN(\mult_20/ab[30][5] ) );
  NOR2_X1 U14225 ( .A1(n3219), .A2(n3206), .ZN(\mult_19/ab[30][3] ) );
  NOR2_X1 U14226 ( .A1(n3216), .A2(n3205), .ZN(\mult_19/ab[30][2] ) );
  NOR2_X1 U14227 ( .A1(n3213), .A2(n3204), .ZN(\mult_19/ab[30][1] ) );
  NOR2_X1 U14228 ( .A1(n3402), .A2(n3391), .ZN(\mult_20/ab[30][2] ) );
  NOR2_X1 U14229 ( .A1(n3399), .A2(n3390), .ZN(\mult_20/ab[30][1] ) );
  NOR2_X1 U14230 ( .A1(n3432), .A2(n3390), .ZN(\mult_20/ab[30][12] ) );
  NOR2_X1 U14231 ( .A1(n3246), .A2(n3204), .ZN(\mult_19/ab[30][12] ) );
  NOR2_X1 U14232 ( .A1(n3398), .A2(n3318), .ZN(\mult_20/ab[6][0] ) );
  NOR2_X1 U14233 ( .A1(n3398), .A2(n3321), .ZN(\mult_20/ab[7][0] ) );
  NOR2_X1 U14234 ( .A1(n3398), .A2(n3324), .ZN(\mult_20/ab[8][0] ) );
  NOR2_X1 U14235 ( .A1(n3398), .A2(n3327), .ZN(\mult_20/ab[9][0] ) );
  NOR2_X1 U14236 ( .A1(n3396), .A2(n3330), .ZN(\mult_20/ab[10][0] ) );
  NOR2_X1 U14237 ( .A1(n3396), .A2(n3333), .ZN(\mult_20/ab[11][0] ) );
  NOR2_X1 U14238 ( .A1(n3396), .A2(n3336), .ZN(\mult_20/ab[12][0] ) );
  NOR2_X1 U14239 ( .A1(n3396), .A2(n3339), .ZN(\mult_20/ab[13][0] ) );
  NOR2_X1 U14240 ( .A1(n3396), .A2(n3342), .ZN(\mult_20/ab[14][0] ) );
  NOR2_X1 U14241 ( .A1(n3396), .A2(n3345), .ZN(\mult_20/ab[15][0] ) );
  NOR2_X1 U14242 ( .A1(n3396), .A2(n3348), .ZN(\mult_20/ab[16][0] ) );
  NOR2_X1 U14243 ( .A1(n3396), .A2(n3351), .ZN(\mult_20/ab[17][0] ) );
  NOR2_X1 U14244 ( .A1(n3396), .A2(n3354), .ZN(\mult_20/ab[18][0] ) );
  NOR2_X1 U14245 ( .A1(n3396), .A2(n3357), .ZN(\mult_20/ab[19][0] ) );
  NOR2_X1 U14246 ( .A1(n3396), .A2(n3360), .ZN(\mult_20/ab[20][0] ) );
  NOR2_X1 U14247 ( .A1(n3397), .A2(n3363), .ZN(\mult_20/ab[21][0] ) );
  NOR2_X1 U14248 ( .A1(n3397), .A2(n3366), .ZN(\mult_20/ab[22][0] ) );
  NOR2_X1 U14249 ( .A1(n3397), .A2(n3369), .ZN(\mult_20/ab[23][0] ) );
  NOR2_X1 U14250 ( .A1(n3397), .A2(n3372), .ZN(\mult_20/ab[24][0] ) );
  NOR2_X1 U14251 ( .A1(n3397), .A2(n3375), .ZN(\mult_20/ab[25][0] ) );
  NOR2_X1 U14252 ( .A1(n3397), .A2(n3378), .ZN(\mult_20/ab[26][0] ) );
  NOR2_X1 U14253 ( .A1(n3397), .A2(n3381), .ZN(\mult_20/ab[27][0] ) );
  NOR2_X1 U14254 ( .A1(n3397), .A2(n3384), .ZN(\mult_20/ab[28][0] ) );
  NOR2_X1 U14255 ( .A1(n3397), .A2(n3387), .ZN(\mult_20/ab[29][0] ) );
  NOR2_X1 U14256 ( .A1(n3397), .A2(n3390), .ZN(\mult_20/ab[30][0] ) );
  NOR2_X1 U14257 ( .A1(n3212), .A2(n3132), .ZN(\mult_19/ab[6][0] ) );
  NOR2_X1 U14258 ( .A1(n3212), .A2(n3135), .ZN(\mult_19/ab[7][0] ) );
  NOR2_X1 U14259 ( .A1(n3212), .A2(n3138), .ZN(\mult_19/ab[8][0] ) );
  NOR2_X1 U14260 ( .A1(n3212), .A2(n3141), .ZN(\mult_19/ab[9][0] ) );
  NOR2_X1 U14261 ( .A1(n3210), .A2(n3144), .ZN(\mult_19/ab[10][0] ) );
  NOR2_X1 U14262 ( .A1(n3210), .A2(n3147), .ZN(\mult_19/ab[11][0] ) );
  NOR2_X1 U14263 ( .A1(n3210), .A2(n3150), .ZN(\mult_19/ab[12][0] ) );
  NOR2_X1 U14264 ( .A1(n3210), .A2(n3153), .ZN(\mult_19/ab[13][0] ) );
  NOR2_X1 U14265 ( .A1(n3210), .A2(n3156), .ZN(\mult_19/ab[14][0] ) );
  NOR2_X1 U14266 ( .A1(n3210), .A2(n3159), .ZN(\mult_19/ab[15][0] ) );
  NOR2_X1 U14267 ( .A1(n3210), .A2(n3162), .ZN(\mult_19/ab[16][0] ) );
  NOR2_X1 U14268 ( .A1(n3210), .A2(n3165), .ZN(\mult_19/ab[17][0] ) );
  NOR2_X1 U14269 ( .A1(n3210), .A2(n3168), .ZN(\mult_19/ab[18][0] ) );
  NOR2_X1 U14270 ( .A1(n3210), .A2(n3171), .ZN(\mult_19/ab[19][0] ) );
  NOR2_X1 U14271 ( .A1(n3210), .A2(n3174), .ZN(\mult_19/ab[20][0] ) );
  NOR2_X1 U14272 ( .A1(n3211), .A2(n3177), .ZN(\mult_19/ab[21][0] ) );
  NOR2_X1 U14273 ( .A1(n3211), .A2(n3180), .ZN(\mult_19/ab[22][0] ) );
  NOR2_X1 U14274 ( .A1(n3211), .A2(n3183), .ZN(\mult_19/ab[23][0] ) );
  NOR2_X1 U14275 ( .A1(n3211), .A2(n3186), .ZN(\mult_19/ab[24][0] ) );
  NOR2_X1 U14276 ( .A1(n3211), .A2(n3189), .ZN(\mult_19/ab[25][0] ) );
  NOR2_X1 U14277 ( .A1(n3211), .A2(n3192), .ZN(\mult_19/ab[26][0] ) );
  NOR2_X1 U14278 ( .A1(n3211), .A2(n3195), .ZN(\mult_19/ab[27][0] ) );
  NOR2_X1 U14279 ( .A1(n3211), .A2(n3198), .ZN(\mult_19/ab[28][0] ) );
  NOR2_X1 U14280 ( .A1(n3211), .A2(n3201), .ZN(\mult_19/ab[29][0] ) );
  NOR2_X1 U14281 ( .A1(n3211), .A2(n3204), .ZN(\mult_19/ab[30][0] ) );
  NOR2_X1 U14282 ( .A1(n3468), .A2(n3394), .ZN(\mult_20/ab[31][24] ) );
  NOR2_X1 U14283 ( .A1(n3282), .A2(n3208), .ZN(\mult_19/ab[31][24] ) );
  NOR2_X1 U14284 ( .A1(n3462), .A2(n3394), .ZN(\mult_20/ab[31][22] ) );
  NOR2_X1 U14285 ( .A1(n3276), .A2(n3208), .ZN(\mult_19/ab[31][22] ) );
  NOR2_X1 U14286 ( .A1(n3438), .A2(n3393), .ZN(\mult_20/ab[31][14] ) );
  NOR2_X1 U14287 ( .A1(n3252), .A2(n3207), .ZN(\mult_19/ab[31][14] ) );
  NOR2_X1 U14288 ( .A1(n3444), .A2(n3393), .ZN(\mult_20/ab[31][16] ) );
  NOR2_X1 U14289 ( .A1(n3258), .A2(n3207), .ZN(\mult_19/ab[31][16] ) );
  NOR2_X1 U14290 ( .A1(n3450), .A2(n3393), .ZN(\mult_20/ab[31][18] ) );
  NOR2_X1 U14291 ( .A1(n3264), .A2(n3207), .ZN(\mult_19/ab[31][18] ) );
  NOR2_X1 U14292 ( .A1(n3456), .A2(n3394), .ZN(\mult_20/ab[31][20] ) );
  NOR2_X1 U14293 ( .A1(n3270), .A2(n3208), .ZN(\mult_19/ab[31][20] ) );
  NOR2_X1 U14294 ( .A1(n3447), .A2(n3393), .ZN(\mult_20/ab[31][17] ) );
  NOR2_X1 U14295 ( .A1(n3261), .A2(n3207), .ZN(\mult_19/ab[31][17] ) );
  NOR2_X1 U14296 ( .A1(n3459), .A2(n3394), .ZN(\mult_20/ab[31][21] ) );
  NOR2_X1 U14297 ( .A1(n3273), .A2(n3208), .ZN(\mult_19/ab[31][21] ) );
  NOR2_X1 U14298 ( .A1(n3465), .A2(n3394), .ZN(\mult_20/ab[31][23] ) );
  NOR2_X1 U14299 ( .A1(n3279), .A2(n3208), .ZN(\mult_19/ab[31][23] ) );
  NOR2_X1 U14300 ( .A1(n3471), .A2(n3394), .ZN(\mult_20/ab[31][25] ) );
  NOR2_X1 U14301 ( .A1(n3285), .A2(n3208), .ZN(\mult_19/ab[31][25] ) );
  NOR2_X1 U14302 ( .A1(n3441), .A2(n3393), .ZN(\mult_20/ab[31][15] ) );
  NOR2_X1 U14303 ( .A1(n3255), .A2(n3207), .ZN(\mult_19/ab[31][15] ) );
  NOR2_X1 U14304 ( .A1(n3453), .A2(n3393), .ZN(\mult_20/ab[31][19] ) );
  NOR2_X1 U14305 ( .A1(n3267), .A2(n3207), .ZN(\mult_19/ab[31][19] ) );
  NOR2_X1 U14306 ( .A1(n3489), .A2(n3341), .ZN(\mult_20/ab[13][31] ) );
  NOR2_X1 U14307 ( .A1(n3488), .A2(n3343), .ZN(\mult_20/ab[14][30] ) );
  NOR2_X1 U14308 ( .A1(n3303), .A2(n3155), .ZN(\mult_19/ab[13][31] ) );
  NOR2_X1 U14309 ( .A1(n3302), .A2(n3157), .ZN(\mult_19/ab[14][30] ) );
  NOR2_X1 U14310 ( .A1(n3488), .A2(n3346), .ZN(\mult_20/ab[15][30] ) );
  NOR2_X1 U14311 ( .A1(n3489), .A2(n3344), .ZN(\mult_20/ab[14][31] ) );
  NOR2_X1 U14312 ( .A1(n3302), .A2(n3160), .ZN(\mult_19/ab[15][30] ) );
  NOR2_X1 U14313 ( .A1(n3303), .A2(n3158), .ZN(\mult_19/ab[14][31] ) );
  NOR2_X1 U14314 ( .A1(n3489), .A2(n3347), .ZN(\mult_20/ab[15][31] ) );
  NOR2_X1 U14315 ( .A1(n3488), .A2(n3349), .ZN(\mult_20/ab[16][30] ) );
  NOR2_X1 U14316 ( .A1(n3303), .A2(n3161), .ZN(\mult_19/ab[15][31] ) );
  NOR2_X1 U14317 ( .A1(n3302), .A2(n3163), .ZN(\mult_19/ab[16][30] ) );
  NOR2_X1 U14318 ( .A1(n3489), .A2(n3350), .ZN(\mult_20/ab[16][31] ) );
  NOR2_X1 U14319 ( .A1(n3487), .A2(n3352), .ZN(\mult_20/ab[17][30] ) );
  NOR2_X1 U14320 ( .A1(n3303), .A2(n3164), .ZN(\mult_19/ab[16][31] ) );
  NOR2_X1 U14321 ( .A1(n3301), .A2(n3166), .ZN(\mult_19/ab[17][30] ) );
  NOR2_X1 U14322 ( .A1(n3489), .A2(n3353), .ZN(\mult_20/ab[17][31] ) );
  NOR2_X1 U14323 ( .A1(n3487), .A2(n3355), .ZN(\mult_20/ab[18][30] ) );
  NOR2_X1 U14324 ( .A1(n3303), .A2(n3167), .ZN(\mult_19/ab[17][31] ) );
  NOR2_X1 U14325 ( .A1(n3301), .A2(n3169), .ZN(\mult_19/ab[18][30] ) );
  NOR2_X1 U14326 ( .A1(n3489), .A2(n3356), .ZN(\mult_20/ab[18][31] ) );
  NOR2_X1 U14327 ( .A1(n3487), .A2(n3358), .ZN(\mult_20/ab[19][30] ) );
  NOR2_X1 U14328 ( .A1(n3303), .A2(n3170), .ZN(\mult_19/ab[18][31] ) );
  NOR2_X1 U14329 ( .A1(n3301), .A2(n3172), .ZN(\mult_19/ab[19][30] ) );
  NOR2_X1 U14330 ( .A1(n3489), .A2(n3359), .ZN(\mult_20/ab[19][31] ) );
  NOR2_X1 U14331 ( .A1(n3487), .A2(n3361), .ZN(\mult_20/ab[20][30] ) );
  NOR2_X1 U14332 ( .A1(n3303), .A2(n3173), .ZN(\mult_19/ab[19][31] ) );
  NOR2_X1 U14333 ( .A1(n3301), .A2(n3175), .ZN(\mult_19/ab[20][30] ) );
  NOR2_X1 U14334 ( .A1(n3489), .A2(n3362), .ZN(\mult_20/ab[20][31] ) );
  NOR2_X1 U14335 ( .A1(n3487), .A2(n3364), .ZN(\mult_20/ab[21][30] ) );
  NOR2_X1 U14336 ( .A1(n3303), .A2(n3176), .ZN(\mult_19/ab[20][31] ) );
  NOR2_X1 U14337 ( .A1(n3301), .A2(n3178), .ZN(\mult_19/ab[21][30] ) );
  NOR2_X1 U14338 ( .A1(n3490), .A2(n3365), .ZN(\mult_20/ab[21][31] ) );
  NOR2_X1 U14339 ( .A1(n3487), .A2(n3367), .ZN(\mult_20/ab[22][30] ) );
  NOR2_X1 U14340 ( .A1(n3304), .A2(n3179), .ZN(\mult_19/ab[21][31] ) );
  NOR2_X1 U14341 ( .A1(n3301), .A2(n3181), .ZN(\mult_19/ab[22][30] ) );
  NOR2_X1 U14342 ( .A1(n3490), .A2(n3368), .ZN(\mult_20/ab[22][31] ) );
  NOR2_X1 U14343 ( .A1(n3487), .A2(n3370), .ZN(\mult_20/ab[23][30] ) );
  NOR2_X1 U14344 ( .A1(n3304), .A2(n3182), .ZN(\mult_19/ab[22][31] ) );
  NOR2_X1 U14345 ( .A1(n3301), .A2(n3184), .ZN(\mult_19/ab[23][30] ) );
  NOR2_X1 U14346 ( .A1(n3490), .A2(n3371), .ZN(\mult_20/ab[23][31] ) );
  NOR2_X1 U14347 ( .A1(n3487), .A2(n3373), .ZN(\mult_20/ab[24][30] ) );
  NOR2_X1 U14348 ( .A1(n3304), .A2(n3185), .ZN(\mult_19/ab[23][31] ) );
  NOR2_X1 U14349 ( .A1(n3301), .A2(n3187), .ZN(\mult_19/ab[24][30] ) );
  NOR2_X1 U14350 ( .A1(n3490), .A2(n3374), .ZN(\mult_20/ab[24][31] ) );
  NOR2_X1 U14351 ( .A1(n3487), .A2(n3376), .ZN(\mult_20/ab[25][30] ) );
  NOR2_X1 U14352 ( .A1(n3304), .A2(n3188), .ZN(\mult_19/ab[24][31] ) );
  NOR2_X1 U14353 ( .A1(n3301), .A2(n3190), .ZN(\mult_19/ab[25][30] ) );
  NOR2_X1 U14354 ( .A1(n3490), .A2(n3377), .ZN(\mult_20/ab[25][31] ) );
  NOR2_X1 U14355 ( .A1(n3487), .A2(n3379), .ZN(\mult_20/ab[26][30] ) );
  NOR2_X1 U14356 ( .A1(n3304), .A2(n3191), .ZN(\mult_19/ab[25][31] ) );
  NOR2_X1 U14357 ( .A1(n3301), .A2(n3193), .ZN(\mult_19/ab[26][30] ) );
  NOR2_X1 U14358 ( .A1(n3485), .A2(n3349), .ZN(\mult_20/ab[16][29] ) );
  NOR2_X1 U14359 ( .A1(n3299), .A2(n3163), .ZN(\mult_19/ab[16][29] ) );
  NOR2_X1 U14360 ( .A1(n3481), .A2(n3352), .ZN(\mult_20/ab[17][28] ) );
  NOR2_X1 U14361 ( .A1(n3295), .A2(n3166), .ZN(\mult_19/ab[17][28] ) );
  NOR2_X1 U14362 ( .A1(n3478), .A2(n3355), .ZN(\mult_20/ab[18][27] ) );
  NOR2_X1 U14363 ( .A1(n3485), .A2(n3352), .ZN(\mult_20/ab[17][29] ) );
  NOR2_X1 U14364 ( .A1(n3292), .A2(n3169), .ZN(\mult_19/ab[18][27] ) );
  NOR2_X1 U14365 ( .A1(n3299), .A2(n3166), .ZN(\mult_19/ab[17][29] ) );
  NOR2_X1 U14366 ( .A1(n3475), .A2(n3358), .ZN(\mult_20/ab[19][26] ) );
  NOR2_X1 U14367 ( .A1(n3481), .A2(n3355), .ZN(\mult_20/ab[18][28] ) );
  NOR2_X1 U14368 ( .A1(n3289), .A2(n3172), .ZN(\mult_19/ab[19][26] ) );
  NOR2_X1 U14369 ( .A1(n3295), .A2(n3169), .ZN(\mult_19/ab[18][28] ) );
  NOR2_X1 U14370 ( .A1(n3472), .A2(n3361), .ZN(\mult_20/ab[20][25] ) );
  NOR2_X1 U14371 ( .A1(n3478), .A2(n3358), .ZN(\mult_20/ab[19][27] ) );
  NOR2_X1 U14372 ( .A1(n3286), .A2(n3175), .ZN(\mult_19/ab[20][25] ) );
  NOR2_X1 U14373 ( .A1(n3292), .A2(n3172), .ZN(\mult_19/ab[19][27] ) );
  NOR2_X1 U14374 ( .A1(n3469), .A2(n3364), .ZN(\mult_20/ab[21][24] ) );
  NOR2_X1 U14375 ( .A1(n3475), .A2(n3361), .ZN(\mult_20/ab[20][26] ) );
  NOR2_X1 U14376 ( .A1(n3485), .A2(n3355), .ZN(\mult_20/ab[18][29] ) );
  NOR2_X1 U14377 ( .A1(n3283), .A2(n3178), .ZN(\mult_19/ab[21][24] ) );
  NOR2_X1 U14378 ( .A1(n3289), .A2(n3175), .ZN(\mult_19/ab[20][26] ) );
  NOR2_X1 U14379 ( .A1(n3299), .A2(n3169), .ZN(\mult_19/ab[18][29] ) );
  NOR2_X1 U14380 ( .A1(n3466), .A2(n3367), .ZN(\mult_20/ab[22][23] ) );
  NOR2_X1 U14381 ( .A1(n3472), .A2(n3364), .ZN(\mult_20/ab[21][25] ) );
  NOR2_X1 U14382 ( .A1(n3484), .A2(n3358), .ZN(\mult_20/ab[19][29] ) );
  NOR2_X1 U14383 ( .A1(n3481), .A2(n3358), .ZN(\mult_20/ab[19][28] ) );
  NOR2_X1 U14384 ( .A1(n3280), .A2(n3181), .ZN(\mult_19/ab[22][23] ) );
  NOR2_X1 U14385 ( .A1(n3286), .A2(n3178), .ZN(\mult_19/ab[21][25] ) );
  NOR2_X1 U14386 ( .A1(n3298), .A2(n3172), .ZN(\mult_19/ab[19][29] ) );
  NOR2_X1 U14387 ( .A1(n3295), .A2(n3172), .ZN(\mult_19/ab[19][28] ) );
  NOR2_X1 U14388 ( .A1(n3463), .A2(n3370), .ZN(\mult_20/ab[23][22] ) );
  NOR2_X1 U14389 ( .A1(n3469), .A2(n3367), .ZN(\mult_20/ab[22][24] ) );
  NOR2_X1 U14390 ( .A1(n3481), .A2(n3361), .ZN(\mult_20/ab[20][28] ) );
  NOR2_X1 U14391 ( .A1(n3478), .A2(n3361), .ZN(\mult_20/ab[20][27] ) );
  NOR2_X1 U14392 ( .A1(n3277), .A2(n3184), .ZN(\mult_19/ab[23][22] ) );
  NOR2_X1 U14393 ( .A1(n3283), .A2(n3181), .ZN(\mult_19/ab[22][24] ) );
  NOR2_X1 U14394 ( .A1(n3295), .A2(n3175), .ZN(\mult_19/ab[20][28] ) );
  NOR2_X1 U14395 ( .A1(n3292), .A2(n3175), .ZN(\mult_19/ab[20][27] ) );
  NOR2_X1 U14396 ( .A1(n3460), .A2(n3373), .ZN(\mult_20/ab[24][21] ) );
  NOR2_X1 U14397 ( .A1(n3466), .A2(n3370), .ZN(\mult_20/ab[23][23] ) );
  NOR2_X1 U14398 ( .A1(n3478), .A2(n3364), .ZN(\mult_20/ab[21][27] ) );
  NOR2_X1 U14399 ( .A1(n3475), .A2(n3364), .ZN(\mult_20/ab[21][26] ) );
  NOR2_X1 U14400 ( .A1(n3484), .A2(n3361), .ZN(\mult_20/ab[20][29] ) );
  NOR2_X1 U14401 ( .A1(n3274), .A2(n3187), .ZN(\mult_19/ab[24][21] ) );
  NOR2_X1 U14402 ( .A1(n3280), .A2(n3184), .ZN(\mult_19/ab[23][23] ) );
  NOR2_X1 U14403 ( .A1(n3292), .A2(n3178), .ZN(\mult_19/ab[21][27] ) );
  NOR2_X1 U14404 ( .A1(n3289), .A2(n3178), .ZN(\mult_19/ab[21][26] ) );
  NOR2_X1 U14405 ( .A1(n3298), .A2(n3175), .ZN(\mult_19/ab[20][29] ) );
  NOR2_X1 U14406 ( .A1(n3457), .A2(n3376), .ZN(\mult_20/ab[25][20] ) );
  NOR2_X1 U14407 ( .A1(n3463), .A2(n3373), .ZN(\mult_20/ab[24][22] ) );
  NOR2_X1 U14408 ( .A1(n3475), .A2(n3367), .ZN(\mult_20/ab[22][26] ) );
  NOR2_X1 U14409 ( .A1(n3472), .A2(n3367), .ZN(\mult_20/ab[22][25] ) );
  NOR2_X1 U14410 ( .A1(n3481), .A2(n3364), .ZN(\mult_20/ab[21][28] ) );
  NOR2_X1 U14411 ( .A1(n3271), .A2(n3190), .ZN(\mult_19/ab[25][20] ) );
  NOR2_X1 U14412 ( .A1(n3277), .A2(n3187), .ZN(\mult_19/ab[24][22] ) );
  NOR2_X1 U14413 ( .A1(n3289), .A2(n3181), .ZN(\mult_19/ab[22][26] ) );
  NOR2_X1 U14414 ( .A1(n3286), .A2(n3181), .ZN(\mult_19/ab[22][25] ) );
  NOR2_X1 U14415 ( .A1(n3295), .A2(n3178), .ZN(\mult_19/ab[21][28] ) );
  NOR2_X1 U14416 ( .A1(n3454), .A2(n3378), .ZN(\mult_20/ab[26][19] ) );
  NOR2_X1 U14417 ( .A1(n3460), .A2(n3376), .ZN(\mult_20/ab[25][21] ) );
  NOR2_X1 U14418 ( .A1(n3472), .A2(n3370), .ZN(\mult_20/ab[23][25] ) );
  NOR2_X1 U14419 ( .A1(n3469), .A2(n3370), .ZN(\mult_20/ab[23][24] ) );
  NOR2_X1 U14420 ( .A1(n3478), .A2(n3367), .ZN(\mult_20/ab[22][27] ) );
  NOR2_X1 U14421 ( .A1(n3268), .A2(n3192), .ZN(\mult_19/ab[26][19] ) );
  NOR2_X1 U14422 ( .A1(n3274), .A2(n3190), .ZN(\mult_19/ab[25][21] ) );
  NOR2_X1 U14423 ( .A1(n3286), .A2(n3184), .ZN(\mult_19/ab[23][25] ) );
  NOR2_X1 U14424 ( .A1(n3283), .A2(n3184), .ZN(\mult_19/ab[23][24] ) );
  NOR2_X1 U14425 ( .A1(n3292), .A2(n3181), .ZN(\mult_19/ab[22][27] ) );
  NOR2_X1 U14426 ( .A1(n3451), .A2(n3381), .ZN(\mult_20/ab[27][18] ) );
  NOR2_X1 U14427 ( .A1(n3457), .A2(n3379), .ZN(\mult_20/ab[26][20] ) );
  NOR2_X1 U14428 ( .A1(n3469), .A2(n3373), .ZN(\mult_20/ab[24][24] ) );
  NOR2_X1 U14429 ( .A1(n3466), .A2(n3373), .ZN(\mult_20/ab[24][23] ) );
  NOR2_X1 U14430 ( .A1(n3475), .A2(n3370), .ZN(\mult_20/ab[23][26] ) );
  NOR2_X1 U14431 ( .A1(n3265), .A2(n3195), .ZN(\mult_19/ab[27][18] ) );
  NOR2_X1 U14432 ( .A1(n3271), .A2(n3193), .ZN(\mult_19/ab[26][20] ) );
  NOR2_X1 U14433 ( .A1(n3283), .A2(n3187), .ZN(\mult_19/ab[24][24] ) );
  NOR2_X1 U14434 ( .A1(n3280), .A2(n3187), .ZN(\mult_19/ab[24][23] ) );
  NOR2_X1 U14435 ( .A1(n3289), .A2(n3184), .ZN(\mult_19/ab[23][26] ) );
  NOR2_X1 U14436 ( .A1(n3448), .A2(n3384), .ZN(\mult_20/ab[28][17] ) );
  NOR2_X1 U14437 ( .A1(n3454), .A2(n3381), .ZN(\mult_20/ab[27][19] ) );
  NOR2_X1 U14438 ( .A1(n3466), .A2(n3376), .ZN(\mult_20/ab[25][23] ) );
  NOR2_X1 U14439 ( .A1(n3463), .A2(n3376), .ZN(\mult_20/ab[25][22] ) );
  NOR2_X1 U14440 ( .A1(n3472), .A2(n3373), .ZN(\mult_20/ab[24][25] ) );
  NOR2_X1 U14441 ( .A1(n3484), .A2(n3364), .ZN(\mult_20/ab[21][29] ) );
  NOR2_X1 U14442 ( .A1(n3262), .A2(n3198), .ZN(\mult_19/ab[28][17] ) );
  NOR2_X1 U14443 ( .A1(n3268), .A2(n3195), .ZN(\mult_19/ab[27][19] ) );
  NOR2_X1 U14444 ( .A1(n3280), .A2(n3190), .ZN(\mult_19/ab[25][23] ) );
  NOR2_X1 U14445 ( .A1(n3277), .A2(n3190), .ZN(\mult_19/ab[25][22] ) );
  NOR2_X1 U14446 ( .A1(n3286), .A2(n3187), .ZN(\mult_19/ab[24][25] ) );
  NOR2_X1 U14447 ( .A1(n3298), .A2(n3178), .ZN(\mult_19/ab[21][29] ) );
  NOR2_X1 U14448 ( .A1(n3444), .A2(n3387), .ZN(\mult_20/ab[29][16] ) );
  NOR2_X1 U14449 ( .A1(n3451), .A2(n3384), .ZN(\mult_20/ab[28][18] ) );
  NOR2_X1 U14450 ( .A1(n3463), .A2(n3379), .ZN(\mult_20/ab[26][22] ) );
  NOR2_X1 U14451 ( .A1(n3460), .A2(n3379), .ZN(\mult_20/ab[26][21] ) );
  NOR2_X1 U14452 ( .A1(n3469), .A2(n3376), .ZN(\mult_20/ab[25][24] ) );
  NOR2_X1 U14453 ( .A1(n3484), .A2(n3367), .ZN(\mult_20/ab[22][29] ) );
  NOR2_X1 U14454 ( .A1(n3481), .A2(n3367), .ZN(\mult_20/ab[22][28] ) );
  NOR2_X1 U14455 ( .A1(n3258), .A2(n3201), .ZN(\mult_19/ab[29][16] ) );
  NOR2_X1 U14456 ( .A1(n3265), .A2(n3198), .ZN(\mult_19/ab[28][18] ) );
  NOR2_X1 U14457 ( .A1(n3277), .A2(n3193), .ZN(\mult_19/ab[26][22] ) );
  NOR2_X1 U14458 ( .A1(n3274), .A2(n3193), .ZN(\mult_19/ab[26][21] ) );
  NOR2_X1 U14459 ( .A1(n3283), .A2(n3190), .ZN(\mult_19/ab[25][24] ) );
  NOR2_X1 U14460 ( .A1(n3298), .A2(n3181), .ZN(\mult_19/ab[22][29] ) );
  NOR2_X1 U14461 ( .A1(n3295), .A2(n3181), .ZN(\mult_19/ab[22][28] ) );
  NOR2_X1 U14462 ( .A1(n3441), .A2(n3390), .ZN(\mult_20/ab[30][15] ) );
  NOR2_X1 U14463 ( .A1(n3447), .A2(n3387), .ZN(\mult_20/ab[29][17] ) );
  NOR2_X1 U14464 ( .A1(n3460), .A2(n3382), .ZN(\mult_20/ab[27][21] ) );
  NOR2_X1 U14465 ( .A1(n3457), .A2(n3382), .ZN(\mult_20/ab[27][20] ) );
  NOR2_X1 U14466 ( .A1(n3466), .A2(n3379), .ZN(\mult_20/ab[26][23] ) );
  NOR2_X1 U14467 ( .A1(n3484), .A2(n3370), .ZN(\mult_20/ab[23][29] ) );
  NOR2_X1 U14468 ( .A1(n3481), .A2(n3370), .ZN(\mult_20/ab[23][28] ) );
  NOR2_X1 U14469 ( .A1(n3478), .A2(n3370), .ZN(\mult_20/ab[23][27] ) );
  NOR2_X1 U14470 ( .A1(n3255), .A2(n3204), .ZN(\mult_19/ab[30][15] ) );
  NOR2_X1 U14471 ( .A1(n3261), .A2(n3201), .ZN(\mult_19/ab[29][17] ) );
  NOR2_X1 U14472 ( .A1(n3274), .A2(n3196), .ZN(\mult_19/ab[27][21] ) );
  NOR2_X1 U14473 ( .A1(n3271), .A2(n3196), .ZN(\mult_19/ab[27][20] ) );
  NOR2_X1 U14474 ( .A1(n3280), .A2(n3193), .ZN(\mult_19/ab[26][23] ) );
  NOR2_X1 U14475 ( .A1(n3298), .A2(n3184), .ZN(\mult_19/ab[23][29] ) );
  NOR2_X1 U14476 ( .A1(n3295), .A2(n3184), .ZN(\mult_19/ab[23][28] ) );
  NOR2_X1 U14477 ( .A1(n3292), .A2(n3184), .ZN(\mult_19/ab[23][27] ) );
  NOR2_X1 U14478 ( .A1(n3444), .A2(n3390), .ZN(\mult_20/ab[30][16] ) );
  NOR2_X1 U14479 ( .A1(n3457), .A2(n3385), .ZN(\mult_20/ab[28][20] ) );
  NOR2_X1 U14480 ( .A1(n3454), .A2(n3384), .ZN(\mult_20/ab[28][19] ) );
  NOR2_X1 U14481 ( .A1(n3463), .A2(n3382), .ZN(\mult_20/ab[27][22] ) );
  NOR2_X1 U14482 ( .A1(n3481), .A2(n3373), .ZN(\mult_20/ab[24][28] ) );
  NOR2_X1 U14483 ( .A1(n3478), .A2(n3373), .ZN(\mult_20/ab[24][27] ) );
  NOR2_X1 U14484 ( .A1(n3475), .A2(n3373), .ZN(\mult_20/ab[24][26] ) );
  NOR2_X1 U14485 ( .A1(n3258), .A2(n3204), .ZN(\mult_19/ab[30][16] ) );
  NOR2_X1 U14486 ( .A1(n3271), .A2(n3199), .ZN(\mult_19/ab[28][20] ) );
  NOR2_X1 U14487 ( .A1(n3268), .A2(n3198), .ZN(\mult_19/ab[28][19] ) );
  NOR2_X1 U14488 ( .A1(n3277), .A2(n3196), .ZN(\mult_19/ab[27][22] ) );
  NOR2_X1 U14489 ( .A1(n3295), .A2(n3187), .ZN(\mult_19/ab[24][28] ) );
  NOR2_X1 U14490 ( .A1(n3292), .A2(n3187), .ZN(\mult_19/ab[24][27] ) );
  NOR2_X1 U14491 ( .A1(n3289), .A2(n3187), .ZN(\mult_19/ab[24][26] ) );
  NOR2_X1 U14492 ( .A1(n3453), .A2(n3387), .ZN(\mult_20/ab[29][19] ) );
  NOR2_X1 U14493 ( .A1(n3450), .A2(n3387), .ZN(\mult_20/ab[29][18] ) );
  NOR2_X1 U14494 ( .A1(n3460), .A2(n3385), .ZN(\mult_20/ab[28][21] ) );
  NOR2_X1 U14495 ( .A1(n3478), .A2(n3376), .ZN(\mult_20/ab[25][27] ) );
  NOR2_X1 U14496 ( .A1(n3475), .A2(n3376), .ZN(\mult_20/ab[25][26] ) );
  NOR2_X1 U14497 ( .A1(n3472), .A2(n3376), .ZN(\mult_20/ab[25][25] ) );
  NOR2_X1 U14498 ( .A1(n3267), .A2(n3201), .ZN(\mult_19/ab[29][19] ) );
  NOR2_X1 U14499 ( .A1(n3264), .A2(n3201), .ZN(\mult_19/ab[29][18] ) );
  NOR2_X1 U14500 ( .A1(n3274), .A2(n3199), .ZN(\mult_19/ab[28][21] ) );
  NOR2_X1 U14501 ( .A1(n3292), .A2(n3190), .ZN(\mult_19/ab[25][27] ) );
  NOR2_X1 U14502 ( .A1(n3289), .A2(n3190), .ZN(\mult_19/ab[25][26] ) );
  NOR2_X1 U14503 ( .A1(n3286), .A2(n3190), .ZN(\mult_19/ab[25][25] ) );
  NOR2_X1 U14504 ( .A1(n3447), .A2(n3390), .ZN(\mult_20/ab[30][17] ) );
  NOR2_X1 U14505 ( .A1(n3450), .A2(n3390), .ZN(\mult_20/ab[30][18] ) );
  NOR2_X1 U14506 ( .A1(n3456), .A2(n3388), .ZN(\mult_20/ab[29][20] ) );
  NOR2_X1 U14507 ( .A1(n3475), .A2(n3379), .ZN(\mult_20/ab[26][26] ) );
  NOR2_X1 U14508 ( .A1(n3472), .A2(n3379), .ZN(\mult_20/ab[26][25] ) );
  NOR2_X1 U14509 ( .A1(n3469), .A2(n3379), .ZN(\mult_20/ab[26][24] ) );
  NOR2_X1 U14510 ( .A1(n3484), .A2(n3373), .ZN(\mult_20/ab[24][29] ) );
  NOR2_X1 U14511 ( .A1(n3261), .A2(n3204), .ZN(\mult_19/ab[30][17] ) );
  NOR2_X1 U14512 ( .A1(n3264), .A2(n3204), .ZN(\mult_19/ab[30][18] ) );
  NOR2_X1 U14513 ( .A1(n3270), .A2(n3202), .ZN(\mult_19/ab[29][20] ) );
  NOR2_X1 U14514 ( .A1(n3289), .A2(n3193), .ZN(\mult_19/ab[26][26] ) );
  NOR2_X1 U14515 ( .A1(n3286), .A2(n3193), .ZN(\mult_19/ab[26][25] ) );
  NOR2_X1 U14516 ( .A1(n3283), .A2(n3193), .ZN(\mult_19/ab[26][24] ) );
  NOR2_X1 U14517 ( .A1(n3298), .A2(n3187), .ZN(\mult_19/ab[24][29] ) );
  NOR2_X1 U14518 ( .A1(n3453), .A2(n3390), .ZN(\mult_20/ab[30][19] ) );
  NOR2_X1 U14519 ( .A1(n3472), .A2(n3382), .ZN(\mult_20/ab[27][25] ) );
  NOR2_X1 U14520 ( .A1(n3469), .A2(n3382), .ZN(\mult_20/ab[27][24] ) );
  NOR2_X1 U14521 ( .A1(n3466), .A2(n3382), .ZN(\mult_20/ab[27][23] ) );
  NOR2_X1 U14522 ( .A1(n3484), .A2(n3376), .ZN(\mult_20/ab[25][29] ) );
  NOR2_X1 U14523 ( .A1(n3481), .A2(n3376), .ZN(\mult_20/ab[25][28] ) );
  NOR2_X1 U14524 ( .A1(n3267), .A2(n3204), .ZN(\mult_19/ab[30][19] ) );
  NOR2_X1 U14525 ( .A1(n3286), .A2(n3196), .ZN(\mult_19/ab[27][25] ) );
  NOR2_X1 U14526 ( .A1(n3283), .A2(n3196), .ZN(\mult_19/ab[27][24] ) );
  NOR2_X1 U14527 ( .A1(n3280), .A2(n3196), .ZN(\mult_19/ab[27][23] ) );
  NOR2_X1 U14528 ( .A1(n3298), .A2(n3190), .ZN(\mult_19/ab[25][29] ) );
  NOR2_X1 U14529 ( .A1(n3295), .A2(n3190), .ZN(\mult_19/ab[25][28] ) );
  NOR2_X1 U14530 ( .A1(n3469), .A2(n3385), .ZN(\mult_20/ab[28][24] ) );
  NOR2_X1 U14531 ( .A1(n3465), .A2(n3385), .ZN(\mult_20/ab[28][23] ) );
  NOR2_X1 U14532 ( .A1(n3463), .A2(n3385), .ZN(\mult_20/ab[28][22] ) );
  NOR2_X1 U14533 ( .A1(n3481), .A2(n3379), .ZN(\mult_20/ab[26][28] ) );
  NOR2_X1 U14534 ( .A1(n3478), .A2(n3379), .ZN(\mult_20/ab[26][27] ) );
  NOR2_X1 U14535 ( .A1(n3283), .A2(n3199), .ZN(\mult_19/ab[28][24] ) );
  NOR2_X1 U14536 ( .A1(n3279), .A2(n3199), .ZN(\mult_19/ab[28][23] ) );
  NOR2_X1 U14537 ( .A1(n3277), .A2(n3199), .ZN(\mult_19/ab[28][22] ) );
  NOR2_X1 U14538 ( .A1(n3295), .A2(n3193), .ZN(\mult_19/ab[26][28] ) );
  NOR2_X1 U14539 ( .A1(n3292), .A2(n3193), .ZN(\mult_19/ab[26][27] ) );
  NOR2_X1 U14540 ( .A1(n3459), .A2(n3388), .ZN(\mult_20/ab[29][21] ) );
  NOR2_X1 U14541 ( .A1(n3465), .A2(n3388), .ZN(\mult_20/ab[29][23] ) );
  NOR2_X1 U14542 ( .A1(n3462), .A2(n3388), .ZN(\mult_20/ab[29][22] ) );
  NOR2_X1 U14543 ( .A1(n3478), .A2(n3382), .ZN(\mult_20/ab[27][27] ) );
  NOR2_X1 U14544 ( .A1(n3475), .A2(n3382), .ZN(\mult_20/ab[27][26] ) );
  NOR2_X1 U14545 ( .A1(n3273), .A2(n3202), .ZN(\mult_19/ab[29][21] ) );
  NOR2_X1 U14546 ( .A1(n3279), .A2(n3202), .ZN(\mult_19/ab[29][23] ) );
  NOR2_X1 U14547 ( .A1(n3276), .A2(n3202), .ZN(\mult_19/ab[29][22] ) );
  NOR2_X1 U14548 ( .A1(n3292), .A2(n3196), .ZN(\mult_19/ab[27][27] ) );
  NOR2_X1 U14549 ( .A1(n3289), .A2(n3196), .ZN(\mult_19/ab[27][26] ) );
  NOR2_X1 U14550 ( .A1(n3456), .A2(n3391), .ZN(\mult_20/ab[30][20] ) );
  NOR2_X1 U14551 ( .A1(n3459), .A2(n3391), .ZN(\mult_20/ab[30][21] ) );
  NOR2_X1 U14552 ( .A1(n3462), .A2(n3391), .ZN(\mult_20/ab[30][22] ) );
  NOR2_X1 U14553 ( .A1(n3475), .A2(n3385), .ZN(\mult_20/ab[28][26] ) );
  NOR2_X1 U14554 ( .A1(n3472), .A2(n3385), .ZN(\mult_20/ab[28][25] ) );
  NOR2_X1 U14555 ( .A1(n3484), .A2(n3379), .ZN(\mult_20/ab[26][29] ) );
  NOR2_X1 U14556 ( .A1(n3270), .A2(n3205), .ZN(\mult_19/ab[30][20] ) );
  NOR2_X1 U14557 ( .A1(n3273), .A2(n3205), .ZN(\mult_19/ab[30][21] ) );
  NOR2_X1 U14558 ( .A1(n3276), .A2(n3205), .ZN(\mult_19/ab[30][22] ) );
  NOR2_X1 U14559 ( .A1(n3289), .A2(n3199), .ZN(\mult_19/ab[28][26] ) );
  NOR2_X1 U14560 ( .A1(n3286), .A2(n3199), .ZN(\mult_19/ab[28][25] ) );
  NOR2_X1 U14561 ( .A1(n3298), .A2(n3193), .ZN(\mult_19/ab[26][29] ) );
  NOR2_X1 U14562 ( .A1(n3471), .A2(n3388), .ZN(\mult_20/ab[29][25] ) );
  NOR2_X1 U14563 ( .A1(n3468), .A2(n3388), .ZN(\mult_20/ab[29][24] ) );
  NOR2_X1 U14564 ( .A1(n3481), .A2(n3382), .ZN(\mult_20/ab[27][28] ) );
  NOR2_X1 U14565 ( .A1(n3285), .A2(n3202), .ZN(\mult_19/ab[29][25] ) );
  NOR2_X1 U14566 ( .A1(n3282), .A2(n3202), .ZN(\mult_19/ab[29][24] ) );
  NOR2_X1 U14567 ( .A1(n3295), .A2(n3196), .ZN(\mult_19/ab[27][28] ) );
  NOR2_X1 U14568 ( .A1(n3465), .A2(n3391), .ZN(\mult_20/ab[30][23] ) );
  NOR2_X1 U14569 ( .A1(n3468), .A2(n3391), .ZN(\mult_20/ab[30][24] ) );
  NOR2_X1 U14570 ( .A1(n3478), .A2(n3385), .ZN(\mult_20/ab[28][27] ) );
  NOR2_X1 U14571 ( .A1(n3279), .A2(n3205), .ZN(\mult_19/ab[30][23] ) );
  NOR2_X1 U14572 ( .A1(n3282), .A2(n3205), .ZN(\mult_19/ab[30][24] ) );
  NOR2_X1 U14573 ( .A1(n3292), .A2(n3199), .ZN(\mult_19/ab[28][27] ) );
  NOR2_X1 U14574 ( .A1(n3474), .A2(n3388), .ZN(\mult_20/ab[29][26] ) );
  NOR2_X1 U14575 ( .A1(n3484), .A2(n3382), .ZN(\mult_20/ab[27][29] ) );
  NOR2_X1 U14576 ( .A1(n3288), .A2(n3202), .ZN(\mult_19/ab[29][26] ) );
  NOR2_X1 U14577 ( .A1(n3298), .A2(n3196), .ZN(\mult_19/ab[27][29] ) );
  NOR2_X1 U14578 ( .A1(n3471), .A2(n3391), .ZN(\mult_20/ab[30][25] ) );
  NOR2_X1 U14579 ( .A1(n3481), .A2(n3385), .ZN(\mult_20/ab[28][28] ) );
  NOR2_X1 U14580 ( .A1(n3285), .A2(n3205), .ZN(\mult_19/ab[30][25] ) );
  NOR2_X1 U14581 ( .A1(n3295), .A2(n3199), .ZN(\mult_19/ab[28][28] ) );
  NOR2_X1 U14582 ( .A1(n3477), .A2(n3388), .ZN(\mult_20/ab[29][27] ) );
  NOR2_X1 U14583 ( .A1(n3291), .A2(n3202), .ZN(\mult_19/ab[29][27] ) );
  NOR2_X1 U14584 ( .A1(n3474), .A2(n3391), .ZN(\mult_20/ab[30][26] ) );
  NOR2_X1 U14585 ( .A1(n3288), .A2(n3205), .ZN(\mult_19/ab[30][26] ) );
  NOR2_X1 U14586 ( .A1(n3398), .A2(n3309), .ZN(\mult_20/ab[3][0] ) );
  NOR2_X1 U14587 ( .A1(n3398), .A2(n3312), .ZN(\mult_20/ab[4][0] ) );
  NOR2_X1 U14588 ( .A1(n3398), .A2(n3315), .ZN(\mult_20/ab[5][0] ) );
  NOR2_X1 U14589 ( .A1(n3212), .A2(n3123), .ZN(\mult_19/ab[3][0] ) );
  NOR2_X1 U14590 ( .A1(n3212), .A2(n3126), .ZN(\mult_19/ab[4][0] ) );
  NOR2_X1 U14591 ( .A1(n3212), .A2(n3129), .ZN(\mult_19/ab[5][0] ) );
  NOR2_X1 U14592 ( .A1(n3474), .A2(n3394), .ZN(\mult_20/ab[31][26] ) );
  NOR2_X1 U14593 ( .A1(n3288), .A2(n3208), .ZN(\mult_19/ab[31][26] ) );
  NOR2_X1 U14594 ( .A1(n3480), .A2(n3394), .ZN(\mult_20/ab[31][28] ) );
  NOR2_X1 U14595 ( .A1(n3294), .A2(n3208), .ZN(\mult_19/ab[31][28] ) );
  NOR2_X1 U14596 ( .A1(n3490), .A2(n3392), .ZN(\mult_20/ab[30][31] ) );
  NOR2_X1 U14597 ( .A1(n3486), .A2(n3394), .ZN(\mult_20/ab[31][30] ) );
  NOR2_X1 U14598 ( .A1(n3304), .A2(n3206), .ZN(\mult_19/ab[30][31] ) );
  NOR2_X1 U14599 ( .A1(n3300), .A2(n3208), .ZN(\mult_19/ab[31][30] ) );
  NOR2_X1 U14600 ( .A1(n3477), .A2(n3394), .ZN(\mult_20/ab[31][27] ) );
  NOR2_X1 U14601 ( .A1(n3291), .A2(n3208), .ZN(\mult_19/ab[31][27] ) );
  NOR2_X1 U14602 ( .A1(n3483), .A2(n3394), .ZN(\mult_20/ab[31][29] ) );
  NOR2_X1 U14603 ( .A1(n3297), .A2(n3208), .ZN(\mult_19/ab[31][29] ) );
  NOR2_X1 U14604 ( .A1(n3490), .A2(n3380), .ZN(\mult_20/ab[26][31] ) );
  NOR2_X1 U14605 ( .A1(n3487), .A2(n3382), .ZN(\mult_20/ab[27][30] ) );
  NOR2_X1 U14606 ( .A1(n3304), .A2(n3194), .ZN(\mult_19/ab[26][31] ) );
  NOR2_X1 U14607 ( .A1(n3301), .A2(n3196), .ZN(\mult_19/ab[27][30] ) );
  NOR2_X1 U14608 ( .A1(n3490), .A2(n3383), .ZN(\mult_20/ab[27][31] ) );
  NOR2_X1 U14609 ( .A1(n3487), .A2(n3385), .ZN(\mult_20/ab[28][30] ) );
  NOR2_X1 U14610 ( .A1(n3304), .A2(n3197), .ZN(\mult_19/ab[27][31] ) );
  NOR2_X1 U14611 ( .A1(n3301), .A2(n3199), .ZN(\mult_19/ab[28][30] ) );
  NOR2_X1 U14612 ( .A1(n3490), .A2(n3386), .ZN(\mult_20/ab[28][31] ) );
  NOR2_X1 U14613 ( .A1(n3486), .A2(n3388), .ZN(\mult_20/ab[29][30] ) );
  NOR2_X1 U14614 ( .A1(n3304), .A2(n3200), .ZN(\mult_19/ab[28][31] ) );
  NOR2_X1 U14615 ( .A1(n3300), .A2(n3202), .ZN(\mult_19/ab[29][30] ) );
  NOR2_X1 U14616 ( .A1(n3490), .A2(n3389), .ZN(\mult_20/ab[29][31] ) );
  NOR2_X1 U14617 ( .A1(n3486), .A2(n3391), .ZN(\mult_20/ab[30][30] ) );
  NOR2_X1 U14618 ( .A1(n3304), .A2(n3203), .ZN(\mult_19/ab[29][31] ) );
  NOR2_X1 U14619 ( .A1(n3300), .A2(n3205), .ZN(\mult_19/ab[30][30] ) );
  NOR2_X1 U14620 ( .A1(n3484), .A2(n3385), .ZN(\mult_20/ab[28][29] ) );
  NOR2_X1 U14621 ( .A1(n3298), .A2(n3199), .ZN(\mult_19/ab[28][29] ) );
  NOR2_X1 U14622 ( .A1(n3480), .A2(n3388), .ZN(\mult_20/ab[29][28] ) );
  NOR2_X1 U14623 ( .A1(n3294), .A2(n3202), .ZN(\mult_19/ab[29][28] ) );
  NOR2_X1 U14624 ( .A1(n3477), .A2(n3391), .ZN(\mult_20/ab[30][27] ) );
  NOR2_X1 U14625 ( .A1(n3291), .A2(n3205), .ZN(\mult_19/ab[30][27] ) );
  NOR2_X1 U14626 ( .A1(n3484), .A2(n3388), .ZN(\mult_20/ab[29][29] ) );
  NOR2_X1 U14627 ( .A1(n3298), .A2(n3202), .ZN(\mult_19/ab[29][29] ) );
  NOR2_X1 U14628 ( .A1(n3480), .A2(n3391), .ZN(\mult_20/ab[30][28] ) );
  NOR2_X1 U14629 ( .A1(n3294), .A2(n3205), .ZN(\mult_19/ab[30][28] ) );
  NOR2_X1 U14630 ( .A1(n3483), .A2(n3391), .ZN(\mult_20/ab[30][29] ) );
  NOR2_X1 U14631 ( .A1(n3297), .A2(n3205), .ZN(\mult_19/ab[30][29] ) );
  INV_X1 U14632 ( .A(n1636), .ZN(n394) );
  INV_X1 U14633 ( .A(n1110), .ZN(n488) );
  BUF_X1 U14634 ( .A(n1827), .Z(n2763) );
  BUF_X1 U14635 ( .A(n1827), .Z(n2764) );
  BUF_X1 U14636 ( .A(n2363), .Z(n2654) );
  BUF_X1 U14637 ( .A(n2359), .Z(n2678) );
  BUF_X1 U14638 ( .A(n1821), .Z(n2686) );
  BUF_X1 U14639 ( .A(n1821), .Z(n2687) );
  BUF_X1 U14640 ( .A(n2359), .Z(n2681) );
  BUF_X1 U14641 ( .A(n754), .Z(n2702) );
  BUF_X1 U14642 ( .A(n2360), .Z(n2669) );
  BUF_X1 U14643 ( .A(n1826), .Z(n2673) );
  BUF_X1 U14644 ( .A(n753), .Z(n2708) );
  BUF_X1 U14645 ( .A(n2361), .Z(n2663) );
  BUF_X1 U14646 ( .A(n2359), .Z(n2680) );
  BUF_X1 U14647 ( .A(n2363), .Z(n2657) );
  BUF_X1 U14648 ( .A(n2362), .Z(n2649) );
  BUF_X1 U14649 ( .A(n2158), .Z(n2738) );
  BUF_X1 U14650 ( .A(n2360), .Z(n2668) );
  BUF_X1 U14651 ( .A(n1826), .Z(n2674) );
  BUF_X1 U14652 ( .A(n1813), .Z(n2645) );
  BUF_X1 U14653 ( .A(n1825), .Z(n2637) );
  BUF_X1 U14654 ( .A(n748), .Z(n2733) );
  BUF_X1 U14655 ( .A(n2361), .Z(n2662) );
  BUF_X1 U14656 ( .A(n1818), .Z(n2633) );
  BUF_X1 U14657 ( .A(n1824), .Z(n2625) );
  BUF_X1 U14658 ( .A(n2363), .Z(n2656) );
  BUF_X1 U14659 ( .A(n1812), .Z(n2621) );
  BUF_X1 U14660 ( .A(n1882), .Z(n2610) );
  BUF_X1 U14661 ( .A(n2362), .Z(n2650) );
  BUF_X1 U14662 ( .A(n1820), .Z(n2615) );
  CLKBUF_X1 U14663 ( .A(n1809), .Z(n2695) );
  NOR3_X1 U14664 ( .A1(n2133), .A2(n886), .A3(n2369), .ZN(\mult_22/n60 ) );
  NOR2_X1 U14665 ( .A1(n2599), .A2(n2882), .ZN(\mult_22/ab[24][36] ) );
  XNOR2_X1 U14666 ( .A(\mult_22/CARRYB[22][37] ), .B(n948), .ZN(n947) );
  BUF_X2 U14667 ( .A(n1809), .Z(n2699) );
  NOR2_X1 U14668 ( .A1(n2615), .A2(n2155), .ZN(\mult_22/ab[2][39] ) );
  NOR3_X1 U14669 ( .A1(n822), .A2(n3510), .A3(n2612), .ZN(\mult_22/n24 ) );
  NOR2_X1 U14670 ( .A1(n2592), .A2(n2157), .ZN(\mult_22/ab[2][35] ) );
  NOR3_X1 U14671 ( .A1(n814), .A2(n3511), .A3(n2589), .ZN(\mult_22/n28 ) );
  NOR2_X1 U14672 ( .A1(n2563), .A2(n2153), .ZN(\mult_22/ab[2][30] ) );
  NOR2_X1 U14673 ( .A1(n2625), .A2(n2153), .ZN(\mult_22/ab[2][41] ) );
  NOR2_X1 U14674 ( .A1(n2569), .A2(n2147), .ZN(\mult_22/ab[2][31] ) );
  NOR3_X1 U14675 ( .A1(n870), .A2(n3503), .A3(n2566), .ZN(\mult_22/n15 ) );
  NOR2_X1 U14676 ( .A1(n2610), .A2(n2147), .ZN(\mult_22/ab[2][38] ) );
  NOR3_X1 U14677 ( .A1(n820), .A2(n3503), .A3(n2607), .ZN(\mult_22/n25 ) );
  NOR2_X1 U14678 ( .A1(n2695), .A2(n2758), .ZN(\mult_22/ab[3][53] ) );
  NOR2_X1 U14679 ( .A1(n2616), .A2(n2858), .ZN(\mult_22/ab[20][39] ) );
  NOR2_X1 U14680 ( .A1(n2611), .A2(n2858), .ZN(\mult_22/ab[20][38] ) );
  NOR2_X1 U14681 ( .A1(n3504), .A2(n2748), .ZN(\mult_22/ab[1][63] ) );
  NOR3_X1 U14682 ( .A1(n2141), .A2(n2742), .A3(n2369), .ZN(\mult_22/n181 ) );
  NOR2_X1 U14683 ( .A1(n2687), .A2(n2154), .ZN(\mult_22/ab[2][51] ) );
  NOR3_X1 U14684 ( .A1(n880), .A2(n3512), .A3(n2684), .ZN(\mult_22/n10 ) );
  NOR2_X1 U14685 ( .A1(n2593), .A2(n2870), .ZN(\mult_22/ab[22][35] ) );
  OAI21_X1 U14686 ( .B1(\mult_22/CARRYB[20][36] ), .B2(n952), .A(n953), .ZN(
        n951) );
  NOR2_X1 U14687 ( .A1(n2637), .A2(n2151), .ZN(\mult_22/ab[2][43] ) );
  NOR3_X1 U14688 ( .A1(n889), .A2(n3497), .A3(n2642), .ZN(\mult_22/n57 ) );
  NOR2_X1 U14689 ( .A1(n2649), .A2(n2149), .ZN(\mult_22/ab[2][45] ) );
  NOR3_X1 U14690 ( .A1(n2654), .A2(n3497), .A3(n875), .ZN(\mult_22/n68 ) );
  NOR3_X1 U14691 ( .A1(n2684), .A2(n3499), .A3(n851), .ZN(\mult_22/n8 ) );
  NOR2_X1 U14692 ( .A1(n2681), .A2(n2155), .ZN(\mult_22/ab[2][50] ) );
  NOR2_X1 U14693 ( .A1(n2673), .A2(n2157), .ZN(\mult_22/ab[2][49] ) );
  NOR3_X1 U14694 ( .A1(n2678), .A2(n3497), .A3(n830), .ZN(\mult_22/n9 ) );
  NOR2_X1 U14695 ( .A1(n2622), .A2(n2852), .ZN(\mult_22/ab[19][40] ) );
  NOR2_X1 U14696 ( .A1(n2647), .A2(n2817), .ZN(\mult_22/ab[13][44] ) );
  NOR2_X1 U14697 ( .A1(n2648), .A2(n2817), .ZN(\mult_22/ab[13][45] ) );
  NOR2_X1 U14698 ( .A1(n2659), .A2(n2811), .ZN(\mult_22/ab[12][46] ) );
  NOR2_X1 U14699 ( .A1(n2599), .A2(n2876), .ZN(\mult_22/ab[23][36] ) );
  NOR2_X1 U14700 ( .A1(n2593), .A2(n2876), .ZN(\mult_22/ab[23][35] ) );
  NOR2_X1 U14701 ( .A1(n2545), .A2(n2947), .ZN(\mult_22/ab[35][27] ) );
  NOR2_X1 U14702 ( .A1(n2672), .A2(n2799), .ZN(\mult_22/ab[10][49] ) );
  NOR2_X1 U14703 ( .A1(n2671), .A2(n2799), .ZN(\mult_22/ab[10][48] ) );
  NOR2_X1 U14704 ( .A1(n2580), .A2(n2900), .ZN(\mult_22/ab[27][33] ) );
  NOR2_X1 U14705 ( .A1(n2678), .A2(n2793), .ZN(\mult_22/ab[9][50] ) );
  INV_X1 U14706 ( .A(\mult_22/SUMB[7][51] ), .ZN(n732) );
  OAI21_X1 U14707 ( .B1(n701), .B2(n700), .A(n967), .ZN(
        \mult_22/CARRYB[25][35] ) );
  INV_X1 U14708 ( .A(\mult_22/CARRYB[24][35] ), .ZN(n700) );
  NOR2_X1 U14709 ( .A1(n2605), .A2(n2882), .ZN(\mult_22/ab[24][37] ) );
  INV_X1 U14710 ( .A(\mult_22/CARRYB[22][37] ), .ZN(n706) );
  NOR2_X1 U14711 ( .A1(n2586), .A2(n2900), .ZN(\mult_22/ab[27][34] ) );
  NOR2_X1 U14712 ( .A1(n2702), .A2(n2758), .ZN(\mult_22/ab[3][54] ) );
  NOR2_X1 U14713 ( .A1(n2694), .A2(n2769), .ZN(\mult_22/ab[5][52] ) );
  INV_X1 U14714 ( .A(\mult_22/SUMB[3][53] ), .ZN(n738) );
  NOR2_X1 U14715 ( .A1(n2573), .A2(n2888), .ZN(\mult_22/ab[25][32] ) );
  OAI21_X1 U14716 ( .B1(n704), .B2(n703), .A(n968), .ZN(
        \mult_22/CARRYB[24][32] ) );
  INV_X1 U14717 ( .A(\mult_22/SUMB[23][33] ), .ZN(n704) );
  NOR2_X1 U14718 ( .A1(n2611), .A2(n2882), .ZN(\mult_22/ab[24][38] ) );
  NOR2_X1 U14719 ( .A1(n2708), .A2(n2758), .ZN(\mult_22/ab[3][55] ) );
  NOR2_X1 U14720 ( .A1(n2713), .A2(n2788), .ZN(\mult_22/ab[8][56] ) );
  NOR2_X1 U14721 ( .A1(n2714), .A2(n2794), .ZN(\mult_22/ab[9][56] ) );
  NOR2_X1 U14722 ( .A1(n2705), .A2(n2800), .ZN(\mult_22/ab[10][54] ) );
  NOR2_X1 U14723 ( .A1(n2714), .A2(n2776), .ZN(\mult_22/ab[6][56] ) );
  NOR2_X1 U14724 ( .A1(n1881), .A2(n2793), .ZN(\mult_22/ab[9][52] ) );
  NOR2_X1 U14725 ( .A1(n752), .A2(n2770), .ZN(\mult_22/ab[5][56] ) );
  NOR2_X1 U14726 ( .A1(n2691), .A2(n2153), .ZN(\mult_22/ab[2][52] ) );
  NOR2_X1 U14727 ( .A1(n2569), .A2(n2894), .ZN(\mult_22/ab[26][31] ) );
  NOR2_X1 U14728 ( .A1(n2563), .A2(n2894), .ZN(\mult_22/ab[26][30] ) );
  NOR2_X1 U14729 ( .A1(n2684), .A2(n2775), .ZN(\mult_22/ab[6][51] ) );
  NOR2_X1 U14730 ( .A1(n2678), .A2(n2775), .ZN(\mult_22/ab[6][50] ) );
  NOR2_X1 U14731 ( .A1(n2557), .A2(n2917), .ZN(\mult_22/ab[30][29] ) );
  NOR2_X1 U14732 ( .A1(n2539), .A2(n2947), .ZN(\mult_22/ab[35][26] ) );
  NOR2_X1 U14733 ( .A1(n2669), .A2(n2147), .ZN(\mult_22/ab[2][48] ) );
  NOR3_X1 U14734 ( .A1(n828), .A2(n3506), .A3(n2666), .ZN(\mult_22/n67 ) );
  NOR2_X1 U14735 ( .A1(n2551), .A2(n2941), .ZN(\mult_22/ab[34][28] ) );
  OAI21_X1 U14736 ( .B1(n687), .B2(n686), .A(n962), .ZN(
        \mult_22/CARRYB[33][28] ) );
  NOR2_X1 U14737 ( .A1(n2633), .A2(n2147), .ZN(\mult_22/ab[2][42] ) );
  NOR3_X1 U14738 ( .A1(n824), .A2(n3508), .A3(n2630), .ZN(\mult_22/n23 ) );
  NOR2_X1 U14739 ( .A1(n1882), .A2(n2798), .ZN(\mult_22/ab[10][38] ) );
  NOR2_X1 U14740 ( .A1(n2663), .A2(n2156), .ZN(\mult_22/ab[2][47] ) );
  NOR3_X1 U14741 ( .A1(n878), .A2(n3505), .A3(n2660), .ZN(\mult_22/n11 ) );
  NOR2_X1 U14742 ( .A1(n2657), .A2(n2148), .ZN(\mult_22/ab[2][46] ) );
  NOR3_X1 U14743 ( .A1(n892), .A2(n3497), .A3(n2660), .ZN(\mult_22/n5 ) );
  NOR2_X1 U14744 ( .A1(n2621), .A2(n2154), .ZN(\mult_22/ab[2][40] ) );
  NOR3_X1 U14745 ( .A1(n873), .A2(n3509), .A3(n2618), .ZN(\mult_22/n14 ) );
  NOR2_X1 U14746 ( .A1(n2645), .A2(n2150), .ZN(\mult_22/ab[2][44] ) );
  NOR3_X1 U14747 ( .A1(n826), .A2(n3507), .A3(n2642), .ZN(\mult_22/n22 ) );
  NOR2_X1 U14748 ( .A1(n2563), .A2(n2911), .ZN(\mult_22/ab[29][30] ) );
  OAI21_X1 U14749 ( .B1(n694), .B2(n693), .A(n963), .ZN(
        \mult_22/CARRYB[28][30] ) );
  INV_X1 U14750 ( .A(\mult_22/SUMB[27][31] ), .ZN(n694) );
  NOR2_X1 U14751 ( .A1(n2551), .A2(n2917), .ZN(\mult_22/ab[30][28] ) );
  NOR2_X1 U14752 ( .A1(n2713), .A2(n2782), .ZN(\mult_22/ab[7][56] ) );
  NOR2_X1 U14753 ( .A1(n2604), .A2(n2149), .ZN(\mult_22/ab[2][37] ) );
  NOR3_X1 U14754 ( .A1(n818), .A2(n3503), .A3(n2601), .ZN(\mult_22/n26 ) );
  NOR2_X1 U14755 ( .A1(n1883), .A2(n2792), .ZN(\mult_22/ab[9][32] ) );
  NOR2_X1 U14756 ( .A1(n2598), .A2(n2156), .ZN(\mult_22/ab[2][36] ) );
  NOR3_X1 U14757 ( .A1(n816), .A2(n3511), .A3(n2595), .ZN(\mult_22/n27 ) );
  NOR2_X1 U14758 ( .A1(n2586), .A2(n2148), .ZN(\mult_22/ab[2][34] ) );
  NOR3_X1 U14759 ( .A1(n812), .A2(n3511), .A3(n2583), .ZN(\mult_22/n29 ) );
  NOR2_X1 U14760 ( .A1(n2580), .A2(n2150), .ZN(\mult_22/ab[2][33] ) );
  NOR3_X1 U14761 ( .A1(n810), .A2(n3511), .A3(n2577), .ZN(\mult_22/n30 ) );
  NOR2_X1 U14762 ( .A1(n2573), .A2(n2151), .ZN(\mult_22/ab[2][32] ) );
  BUF_X4 U14763 ( .A(n752), .Z(n2712) );
  CLKBUF_X1 U14764 ( .A(n1809), .Z(n2700) );
  BUF_X1 U14765 ( .A(n1829), .Z(n2769) );
  BUF_X1 U14766 ( .A(n1871), .Z(n2805) );
  BUF_X1 U14767 ( .A(n1872), .Z(n2799) );
  BUF_X1 U14768 ( .A(n1828), .Z(n2775) );
  BUF_X1 U14769 ( .A(n1878), .Z(n2781) );
  BUF_X1 U14770 ( .A(n1866), .Z(n2793) );
  BUF_X1 U14771 ( .A(n1866), .Z(n2792) );
  BUF_X1 U14772 ( .A(n1872), .Z(n2798) );
  BUF_X1 U14773 ( .A(n1871), .Z(n2804) );
  BUF_X1 U14774 ( .A(n1861), .Z(n2446) );
  BUF_X1 U14775 ( .A(n1856), .Z(n2554) );
  BUF_X1 U14776 ( .A(n1862), .Z(n2536) );
  BUF_X1 U14777 ( .A(n1837), .Z(n2460) );
  BUF_X1 U14778 ( .A(n1835), .Z(n2472) );
  BUF_X1 U14779 ( .A(n1836), .Z(n2478) );
  BUF_X1 U14780 ( .A(n1843), .Z(n2466) );
  BUF_X1 U14781 ( .A(n1842), .Z(n2484) );
  BUF_X1 U14782 ( .A(n1841), .Z(n2490) );
  BUF_X1 U14783 ( .A(n1863), .Z(n2454) );
  BUF_X1 U14784 ( .A(n1840), .Z(n2496) );
  BUF_X1 U14785 ( .A(n1861), .Z(n2448) );
  BUF_X1 U14786 ( .A(n1839), .Z(n2502) );
  BUF_X1 U14787 ( .A(n1811), .Z(n2592) );
  BUF_X1 U14788 ( .A(n1819), .Z(n2586) );
  BUF_X1 U14789 ( .A(n1814), .Z(n2604) );
  BUF_X1 U14790 ( .A(n1813), .Z(n2644) );
  BUF_X1 U14791 ( .A(n1825), .Z(n2638) );
  BUF_X1 U14792 ( .A(n1815), .Z(n2598) );
  BUF_X1 U14793 ( .A(n1818), .Z(n2632) );
  BUF_X1 U14794 ( .A(n1883), .Z(n2573) );
  BUF_X1 U14795 ( .A(n1824), .Z(n2626) );
  BUF_X1 U14796 ( .A(n1812), .Z(n2620) );
  BUF_X1 U14797 ( .A(n1882), .Z(n2609) );
  BUF_X1 U14798 ( .A(n1838), .Z(n2508) );
  BUF_X1 U14799 ( .A(n1817), .Z(n2580) );
  BUF_X1 U14800 ( .A(n1820), .Z(n2614) );
  BUF_X1 U14801 ( .A(n1814), .Z(n2603) );
  BUF_X1 U14802 ( .A(n1816), .Z(n2569) );
  BUF_X1 U14803 ( .A(n1815), .Z(n2597) );
  BUF_X1 U14804 ( .A(n1823), .Z(n2563) );
  BUF_X1 U14805 ( .A(n1811), .Z(n2591) );
  BUF_X1 U14806 ( .A(n1819), .Z(n2585) );
  BUF_X1 U14807 ( .A(n1817), .Z(n2579) );
  BUF_X1 U14808 ( .A(n1883), .Z(n2574) );
  BUF_X1 U14809 ( .A(n1868), .Z(n2551) );
  BUF_X1 U14810 ( .A(n1816), .Z(n2568) );
  BUF_X1 U14811 ( .A(n1823), .Z(n2562) );
  BUF_X1 U14812 ( .A(n1834), .Z(n2514) );
  BUF_X1 U14813 ( .A(n1865), .Z(n2545) );
  BUF_X1 U14814 ( .A(n1862), .Z(n2539) );
  BUF_X1 U14815 ( .A(n1856), .Z(n2556) );
  BUF_X1 U14816 ( .A(n1864), .Z(n2533) );
  BUF_X1 U14817 ( .A(n1868), .Z(n2550) );
  BUF_X1 U14818 ( .A(n1873), .Z(n2525) );
  BUF_X1 U14819 ( .A(n1833), .Z(n2521) );
  BUF_X1 U14820 ( .A(n1844), .Z(n2436) );
  BUF_X1 U14821 ( .A(n1834), .Z(n2515) );
  BUF_X1 U14822 ( .A(n1838), .Z(n2509) );
  BUF_X1 U14823 ( .A(n1865), .Z(n2544) );
  BUF_X1 U14824 ( .A(n1839), .Z(n2503) );
  BUF_X1 U14825 ( .A(n1862), .Z(n2538) );
  BUF_X1 U14826 ( .A(n1833), .Z(n2520) );
  BUF_X1 U14827 ( .A(n1840), .Z(n2497) );
  BUF_X1 U14828 ( .A(n1864), .Z(n2532) );
  BUF_X1 U14829 ( .A(n1841), .Z(n2491) );
  BUF_X1 U14830 ( .A(n1873), .Z(n2526) );
  BUF_X1 U14831 ( .A(n1842), .Z(n2485) );
  BUF_X1 U14832 ( .A(n1836), .Z(n2479) );
  BUF_X1 U14833 ( .A(n1835), .Z(n2473) );
  BUF_X1 U14834 ( .A(n1843), .Z(n2467) );
  BUF_X1 U14835 ( .A(n1837), .Z(n2461) );
  BUF_X1 U14836 ( .A(n1863), .Z(n2455) );
  BUF_X1 U14837 ( .A(n1861), .Z(n2449) );
  BUF_X1 U14838 ( .A(n1874), .Z(n2441) );
  BUF_X1 U14839 ( .A(n1844), .Z(n2437) );
  BUF_X1 U14840 ( .A(n1845), .Z(n2431) );
  BUF_X1 U14841 ( .A(n1845), .Z(n2430) );
  BUF_X1 U14842 ( .A(n1832), .Z(n2425) );
  BUF_X1 U14843 ( .A(n1846), .Z(n2419) );
  BUF_X1 U14844 ( .A(n1874), .Z(n2442) );
  BUF_X1 U14845 ( .A(n1875), .Z(n2405) );
  BUF_X1 U14846 ( .A(n1853), .Z(n2401) );
  BUF_X1 U14847 ( .A(n1832), .Z(n2424) );
  BUF_X1 U14848 ( .A(n1854), .Z(n2395) );
  BUF_X1 U14849 ( .A(n1846), .Z(n2418) );
  BUF_X1 U14850 ( .A(n1847), .Z(n2412) );
  BUF_X1 U14851 ( .A(n1875), .Z(n2406) );
  BUF_X1 U14852 ( .A(n1853), .Z(n2400) );
  BUF_X1 U14853 ( .A(n1855), .Z(n2389) );
  BUF_X1 U14854 ( .A(n1854), .Z(n2394) );
  BUF_X1 U14855 ( .A(n1876), .Z(n2381) );
  BUF_X1 U14856 ( .A(n1877), .Z(n2787) );
  BUF_X1 U14857 ( .A(n1877), .Z(n2788) );
  BUF_X1 U14858 ( .A(n1866), .Z(n2794) );
  BUF_X1 U14859 ( .A(n1871), .Z(n2806) );
  BUF_X1 U14860 ( .A(n1851), .Z(n2812) );
  BUF_X1 U14861 ( .A(n1863), .Z(n2452) );
  BUF_X1 U14862 ( .A(n1868), .Z(n2548) );
  BUF_X1 U14863 ( .A(n1865), .Z(n2542) );
  BUF_X1 U14864 ( .A(n1823), .Z(n2560) );
  BUF_X1 U14865 ( .A(n1864), .Z(n2530) );
  BUF_X1 U14866 ( .A(n1847), .Z(n2413) );
  BUF_X1 U14867 ( .A(n1829), .Z(n2770) );
  BUF_X1 U14868 ( .A(n1828), .Z(n2776) );
  BUF_X1 U14869 ( .A(n1878), .Z(n2782) );
  BUF_X1 U14870 ( .A(n1872), .Z(n2800) );
  NOR2_X1 U14871 ( .A1(n2425), .A2(n2154), .ZN(\mult_22/ab[2][7] ) );
  NOR3_X1 U14872 ( .A1(n835), .A2(n3510), .A3(n2422), .ZN(\mult_22/n53 ) );
  CLKBUF_X1 U14873 ( .A(n1809), .Z(n2697) );
  NOR2_X1 U14874 ( .A1(n2521), .A2(n2148), .ZN(\mult_22/ab[2][23] ) );
  NOR3_X1 U14875 ( .A1(n858), .A2(n3511), .A3(n2518), .ZN(\mult_22/n39 ) );
  NOR2_X1 U14876 ( .A1(n2515), .A2(n2150), .ZN(\mult_22/ab[2][22] ) );
  NOR3_X1 U14877 ( .A1(n856), .A2(n3503), .A3(n2512), .ZN(\mult_22/n40 ) );
  NOR2_X1 U14878 ( .A1(n2449), .A2(n2150), .ZN(\mult_22/ab[2][11] ) );
  NOR2_X1 U14879 ( .A1(n2473), .A2(n2148), .ZN(\mult_22/ab[2][15] ) );
  NOR3_X1 U14880 ( .A1(n843), .A2(n3511), .A3(n2470), .ZN(\mult_22/n46 ) );
  NOR2_X1 U14881 ( .A1(n2461), .A2(n2157), .ZN(\mult_22/ab[2][13] ) );
  NOR3_X1 U14882 ( .A1(n841), .A2(n3509), .A3(n2458), .ZN(\mult_22/n47 ) );
  NOR2_X1 U14883 ( .A1(n2557), .A2(n2154), .ZN(\mult_22/ab[2][29] ) );
  NOR2_X1 U14884 ( .A1(n2539), .A2(n2149), .ZN(\mult_22/ab[2][26] ) );
  NOR2_X1 U14885 ( .A1(n2525), .A2(n2147), .ZN(\mult_22/ab[2][24] ) );
  NOR2_X1 U14886 ( .A1(n2479), .A2(n2147), .ZN(\mult_22/ab[2][16] ) );
  NOR3_X1 U14887 ( .A1(n845), .A2(n3503), .A3(n2476), .ZN(\mult_22/n45 ) );
  NOR2_X1 U14888 ( .A1(n2455), .A2(n2149), .ZN(\mult_22/ab[2][12] ) );
  NOR3_X1 U14889 ( .A1(n894), .A2(n3497), .A3(n2458), .ZN(\mult_22/n48 ) );
  NOR2_X1 U14890 ( .A1(n2441), .A2(n2151), .ZN(\mult_22/ab[2][10] ) );
  NOR3_X1 U14891 ( .A1(n2446), .A2(n3497), .A3(n891), .ZN(\mult_22/n50 ) );
  NOR2_X1 U14892 ( .A1(n2405), .A2(n2148), .ZN(\mult_22/ab[2][4] ) );
  NOR2_X1 U14893 ( .A1(n2551), .A2(n2156), .ZN(\mult_22/ab[2][28] ) );
  NOR3_X1 U14894 ( .A1(n2554), .A2(n3497), .A3(n899), .ZN(\mult_22/n34 ) );
  NOR2_X1 U14895 ( .A1(n2545), .A2(n2157), .ZN(\mult_22/ab[2][27] ) );
  NOR2_X1 U14896 ( .A1(n2533), .A2(n2155), .ZN(\mult_22/ab[2][25] ) );
  NOR3_X1 U14897 ( .A1(n2536), .A2(n3497), .A3(n896), .ZN(\mult_22/n37 ) );
  NOR2_X1 U14898 ( .A1(n2509), .A2(n2151), .ZN(\mult_22/ab[2][21] ) );
  NOR3_X1 U14899 ( .A1(n854), .A2(n3511), .A3(n2506), .ZN(\mult_22/n41 ) );
  NOR2_X1 U14900 ( .A1(n2503), .A2(n2147), .ZN(\mult_22/ab[2][20] ) );
  NOR3_X1 U14901 ( .A1(n852), .A2(n3503), .A3(n2500), .ZN(\mult_22/n42 ) );
  NOR2_X1 U14902 ( .A1(n2497), .A2(n2153), .ZN(\mult_22/ab[2][19] ) );
  NOR3_X1 U14903 ( .A1(n868), .A2(n3503), .A3(n2494), .ZN(\mult_22/n16 ) );
  NOR2_X1 U14904 ( .A1(n2491), .A2(n2154), .ZN(\mult_22/ab[2][18] ) );
  NOR3_X1 U14905 ( .A1(n849), .A2(n3511), .A3(n2488), .ZN(\mult_22/n43 ) );
  NOR2_X1 U14906 ( .A1(n2485), .A2(n2155), .ZN(\mult_22/ab[2][17] ) );
  NOR3_X1 U14907 ( .A1(n847), .A2(n3510), .A3(n2482), .ZN(\mult_22/n44 ) );
  NOR2_X1 U14908 ( .A1(n2467), .A2(n2156), .ZN(\mult_22/ab[2][14] ) );
  NOR3_X1 U14909 ( .A1(n866), .A2(n3510), .A3(n2464), .ZN(\mult_22/n17 ) );
  NOR2_X1 U14910 ( .A1(n2437), .A2(n2147), .ZN(\mult_22/ab[2][9] ) );
  NOR3_X1 U14911 ( .A1(n839), .A2(n3511), .A3(n2434), .ZN(\mult_22/n51 ) );
  NOR2_X1 U14912 ( .A1(n2431), .A2(n2153), .ZN(\mult_22/ab[2][8] ) );
  NOR3_X1 U14913 ( .A1(n837), .A2(n3503), .A3(n2428), .ZN(\mult_22/n52 ) );
  NOR2_X1 U14914 ( .A1(n2419), .A2(n2156), .ZN(\mult_22/ab[2][6] ) );
  NOR3_X1 U14915 ( .A1(n864), .A2(n3503), .A3(n2416), .ZN(\mult_22/n18 ) );
  NOR3_X1 U14916 ( .A1(n833), .A2(n3503), .A3(n2410), .ZN(\mult_22/n54 ) );
  NOR2_X1 U14917 ( .A1(n2401), .A2(n2155), .ZN(\mult_22/ab[2][3] ) );
  NOR3_X1 U14918 ( .A1(n862), .A2(n3503), .A3(n2398), .ZN(\mult_22/n19 ) );
  NOR2_X1 U14919 ( .A1(n2395), .A2(n2147), .ZN(\mult_22/ab[2][2] ) );
  NOR3_X1 U14920 ( .A1(n860), .A2(n3509), .A3(n2392), .ZN(\mult_22/n20 ) );
  NOR2_X1 U14921 ( .A1(n2389), .A2(n2149), .ZN(\mult_22/ab[2][1] ) );
  NOR3_X1 U14922 ( .A1(n831), .A2(n3511), .A3(n2386), .ZN(\mult_22/n56 ) );
  NOR2_X1 U14923 ( .A1(n2381), .A2(n2150), .ZN(\mult_22/ab[2][0] ) );
  NOR3_X1 U14924 ( .A1(n907), .A2(n3499), .A3(n2386), .ZN(\mult_22/n21 ) );
  BUF_X1 U14925 ( .A(n1857), .Z(n2864) );
  BUF_X1 U14926 ( .A(n1870), .Z(n2840) );
  BUF_X1 U14927 ( .A(n1867), .Z(n2834) );
  BUF_X1 U14928 ( .A(n1869), .Z(n2846) );
  BUF_X1 U14929 ( .A(n1848), .Z(n2828) );
  BUF_X1 U14930 ( .A(n1867), .Z(n2835) );
  BUF_X1 U14931 ( .A(n1849), .Z(n2822) );
  BUF_X1 U14932 ( .A(n1850), .Z(n2816) );
  BUF_X1 U14933 ( .A(n1859), .Z(n2858) );
  BUF_X1 U14934 ( .A(n1851), .Z(n2810) );
  BUF_X1 U14935 ( .A(n1870), .Z(n2841) );
  BUF_X1 U14936 ( .A(n1869), .Z(n2847) );
  BUF_X1 U14937 ( .A(n1859), .Z(n2857) );
  BUF_X1 U14938 ( .A(n1857), .Z(n2862) );
  BUF_X1 U14939 ( .A(n1857), .Z(n2865) );
  BUF_X1 U14940 ( .A(n1858), .Z(n2871) );
  BUF_X1 U14941 ( .A(n1852), .Z(n2853) );
  BUF_X1 U14942 ( .A(n1859), .Z(n2859) );
  BUF_X1 U14943 ( .A(n1858), .Z(n2869) );
  BUF_X1 U14944 ( .A(n1887), .Z(n2875) );
  BUF_X1 U14945 ( .A(n1858), .Z(n2870) );
  BUF_X1 U14946 ( .A(n1886), .Z(n2881) );
  BUF_X1 U14947 ( .A(n1887), .Z(n2877) );
  BUF_X1 U14948 ( .A(n1887), .Z(n2876) );
  BUF_X1 U14949 ( .A(n1893), .Z(n2887) );
  BUF_X1 U14950 ( .A(n1886), .Z(n2883) );
  BUF_X1 U14951 ( .A(n1886), .Z(n2882) );
  BUF_X1 U14952 ( .A(n1893), .Z(n2889) );
  BUF_X1 U14953 ( .A(n1893), .Z(n2888) );
  BUF_X1 U14954 ( .A(n1892), .Z(n2899) );
  BUF_X1 U14955 ( .A(n1860), .Z(n2895) );
  BUF_X1 U14956 ( .A(n1860), .Z(n2894) );
  BUF_X1 U14957 ( .A(n1892), .Z(n2901) );
  BUF_X1 U14958 ( .A(n1892), .Z(n2900) );
  BUF_X1 U14959 ( .A(n1891), .Z(n2906) );
  BUF_X1 U14960 ( .A(n1859), .Z(n2856) );
  BUF_X1 U14961 ( .A(n1858), .Z(n2868) );
  BUF_X1 U14962 ( .A(n1887), .Z(n2874) );
  BUF_X1 U14963 ( .A(n1857), .Z(n2866) );
  BUF_X1 U14964 ( .A(n1886), .Z(n2880) );
  BUF_X1 U14965 ( .A(n1857), .Z(n2863) );
  BUF_X1 U14966 ( .A(n1858), .Z(n2872) );
  BUF_X1 U14967 ( .A(n1893), .Z(n2886) );
  BUF_X1 U14968 ( .A(n1887), .Z(n2878) );
  BUF_X1 U14969 ( .A(n1886), .Z(n2884) );
  BUF_X1 U14970 ( .A(n1860), .Z(n2893) );
  BUF_X1 U14971 ( .A(n1855), .Z(n2388) );
  BUF_X1 U14972 ( .A(n1876), .Z(n2382) );
  BUF_X1 U14973 ( .A(n1860), .Z(n2892) );
  BUF_X1 U14974 ( .A(n1850), .Z(n2818) );
  BUF_X1 U14975 ( .A(n1849), .Z(n2824) );
  BUF_X1 U14976 ( .A(n1848), .Z(n2830) );
  BUF_X1 U14977 ( .A(n1867), .Z(n2836) );
  BUF_X1 U14978 ( .A(n1859), .Z(n2860) );
  BUF_X1 U14979 ( .A(n1870), .Z(n2842) );
  BUF_X1 U14980 ( .A(n1869), .Z(n2848) );
  BUF_X1 U14981 ( .A(n1852), .Z(n2854) );
  NOR2_X1 U14982 ( .A1(n2704), .A2(n3118), .ZN(\mult_22/ab[63][54] ) );
  NOR2_X1 U14983 ( .A1(n2699), .A2(n3094), .ZN(\mult_22/ab[59][53] ) );
  BUF_X1 U14984 ( .A(n1891), .Z(n2905) );
  BUF_X1 U14985 ( .A(n1891), .Z(n2907) );
  BUF_X1 U14986 ( .A(n1890), .Z(n2911) );
  BUF_X1 U14987 ( .A(n1890), .Z(n2913) );
  BUF_X1 U14988 ( .A(n1890), .Z(n2912) );
  BUF_X1 U14989 ( .A(n1889), .Z(n2917) );
  BUF_X1 U14990 ( .A(n1889), .Z(n2919) );
  BUF_X1 U14991 ( .A(n1889), .Z(n2918) );
  BUF_X1 U14992 ( .A(n1900), .Z(n2925) );
  BUF_X1 U14993 ( .A(n1900), .Z(n2923) );
  BUF_X1 U14994 ( .A(n1900), .Z(n2924) );
  BUF_X1 U14995 ( .A(n1888), .Z(n2931) );
  BUF_X1 U14996 ( .A(n1888), .Z(n2929) );
  BUF_X1 U14997 ( .A(n1888), .Z(n2930) );
  BUF_X1 U14998 ( .A(n1899), .Z(n2935) );
  BUF_X1 U14999 ( .A(n1899), .Z(n2936) );
  BUF_X1 U15000 ( .A(n1898), .Z(n2941) );
  BUF_X1 U15001 ( .A(n1898), .Z(n2942) );
  BUF_X1 U15002 ( .A(n1899), .Z(n2937) );
  BUF_X1 U15003 ( .A(n1897), .Z(n2947) );
  BUF_X1 U15004 ( .A(n1897), .Z(n2948) );
  BUF_X1 U15005 ( .A(n1894), .Z(n2953) );
  BUF_X1 U15006 ( .A(n1894), .Z(n2954) );
  BUF_X1 U15007 ( .A(n1892), .Z(n2898) );
  BUF_X1 U15008 ( .A(n1891), .Z(n2904) );
  BUF_X1 U15009 ( .A(n1890), .Z(n2910) );
  BUF_X1 U15010 ( .A(n1889), .Z(n2916) );
  BUF_X1 U15011 ( .A(n1900), .Z(n2922) );
  BUF_X1 U15012 ( .A(n1888), .Z(n2928) );
  BUF_X1 U15013 ( .A(n1899), .Z(n2934) );
  BUF_X1 U15014 ( .A(n1898), .Z(n2940) );
  BUF_X1 U15015 ( .A(n1893), .Z(n2890) );
  BUF_X1 U15016 ( .A(n1860), .Z(n2896) );
  BUF_X1 U15017 ( .A(n1892), .Z(n2902) );
  BUF_X1 U15018 ( .A(n1891), .Z(n2908) );
  BUF_X1 U15019 ( .A(n1890), .Z(n2914) );
  BUF_X1 U15020 ( .A(n1889), .Z(n2920) );
  BUF_X1 U15021 ( .A(n1900), .Z(n2926) );
  BUF_X1 U15022 ( .A(n1888), .Z(n2932) );
  AOI21_X1 U15023 ( .B1(\mult_22/SUMB[63][62] ), .B2(\mult_22/CARRYB[63][61] ), 
        .A(n1287), .ZN(n1285) );
  XNOR2_X1 U15024 ( .A(n1288), .B(\mult_22/CARRYB[63][62] ), .ZN(n1287) );
  NOR2_X1 U15025 ( .A1(n652), .A2(n1288), .ZN(n1281) );
  AND3_X1 U15026 ( .A1(\mult_22/CARRYB[63][61] ), .A2(\mult_22/SUMB[63][62] ), 
        .A3(n1289), .ZN(n1284) );
  AOI21_X1 U15027 ( .B1(n1288), .B2(n652), .A(n1281), .ZN(n1289) );
  INV_X1 U15028 ( .A(n1935), .ZN(n3514) );
  INV_X1 U15029 ( .A(n1936), .ZN(n3525) );
  INV_X1 U15030 ( .A(n1936), .ZN(n3524) );
  INV_X1 U15031 ( .A(n1935), .ZN(n3513) );
  BUF_X1 U15032 ( .A(n1898), .Z(n2943) );
  BUF_X1 U15033 ( .A(n1895), .Z(n2959) );
  BUF_X1 U15034 ( .A(n1895), .Z(n2960) );
  BUF_X1 U15035 ( .A(n1896), .Z(n2965) );
  BUF_X1 U15036 ( .A(n1896), .Z(n2966) );
  BUF_X1 U15037 ( .A(n1897), .Z(n2949) );
  BUF_X1 U15038 ( .A(n1927), .Z(n2971) );
  BUF_X1 U15039 ( .A(n1927), .Z(n2972) );
  BUF_X1 U15040 ( .A(n1894), .Z(n2955) );
  BUF_X1 U15041 ( .A(n1928), .Z(n2978) );
  BUF_X1 U15042 ( .A(n1928), .Z(n2977) );
  BUF_X1 U15043 ( .A(n1895), .Z(n2961) );
  BUF_X1 U15044 ( .A(n1929), .Z(n2984) );
  BUF_X1 U15045 ( .A(n1929), .Z(n2983) );
  BUF_X1 U15046 ( .A(n1896), .Z(n2967) );
  BUF_X1 U15047 ( .A(n1930), .Z(n2990) );
  BUF_X1 U15048 ( .A(n1930), .Z(n2989) );
  BUF_X1 U15049 ( .A(n1931), .Z(n2995) );
  BUF_X1 U15050 ( .A(n1932), .Z(n3001) );
  BUF_X1 U15051 ( .A(n1927), .Z(n2973) );
  BUF_X1 U15052 ( .A(n1928), .Z(n2979) );
  BUF_X1 U15053 ( .A(n1929), .Z(n2985) );
  BUF_X1 U15054 ( .A(n1894), .Z(n2956) );
  BUF_X1 U15055 ( .A(n1895), .Z(n2962) );
  BUF_X1 U15056 ( .A(n1896), .Z(n2968) );
  BUF_X1 U15057 ( .A(n1927), .Z(n2974) );
  BUF_X1 U15058 ( .A(n1928), .Z(n2980) );
  BUF_X1 U15059 ( .A(n1929), .Z(n2986) );
  BUF_X1 U15060 ( .A(n1897), .Z(n2946) );
  BUF_X1 U15061 ( .A(n1894), .Z(n2952) );
  BUF_X1 U15062 ( .A(n1895), .Z(n2958) );
  BUF_X1 U15063 ( .A(n1896), .Z(n2964) );
  BUF_X1 U15064 ( .A(n1927), .Z(n2970) );
  BUF_X1 U15065 ( .A(n1928), .Z(n2976) );
  BUF_X1 U15066 ( .A(n1929), .Z(n2982) );
  BUF_X1 U15067 ( .A(n1930), .Z(n2988) );
  BUF_X1 U15068 ( .A(n1931), .Z(n2994) );
  BUF_X1 U15069 ( .A(n1899), .Z(n2938) );
  BUF_X1 U15070 ( .A(n1898), .Z(n2944) );
  BUF_X1 U15071 ( .A(n1897), .Z(n2950) );
  OAI221_X1 U15072 ( .B1(n1635), .B2(n1636), .C1(n392), .C2(n1637), .A(n1638), 
        .ZN(N127) );
  INV_X1 U15073 ( .A(\mult_20/CARRYB[31][30] ), .ZN(n392) );
  OAI221_X1 U15074 ( .B1(n1109), .B2(n1110), .C1(n486), .C2(n1111), .A(n1112), 
        .ZN(N63) );
  INV_X1 U15075 ( .A(\mult_19/CARRYB[31][30] ), .ZN(n486) );
  BUF_X1 U15076 ( .A(n1923), .Z(n3310) );
  BUF_X1 U15077 ( .A(n1923), .Z(n3309) );
  BUF_X1 U15078 ( .A(n1924), .Z(n3124) );
  BUF_X1 U15079 ( .A(n1924), .Z(n3123) );
  BUF_X1 U15080 ( .A(n1991), .Z(n3313) );
  BUF_X1 U15081 ( .A(n1993), .Z(n3127) );
  BUF_X1 U15082 ( .A(n1992), .Z(n3316) );
  BUF_X1 U15083 ( .A(n1994), .Z(n3130) );
  BUF_X1 U15084 ( .A(n1926), .Z(n3121) );
  BUF_X1 U15085 ( .A(n1925), .Z(n3307) );
  BUF_X1 U15086 ( .A(n1925), .Z(n3306) );
  BUF_X1 U15087 ( .A(n1926), .Z(n3120) );
  NOR2_X1 U15088 ( .A1(n3465), .A2(n3307), .ZN(\mult_20/ab[2][23] ) );
  NOR3_X1 U15089 ( .A1(n3468), .A2(n978), .A3(n1935), .ZN(\mult_20/n9 ) );
  NOR2_X1 U15090 ( .A1(n3294), .A2(n3121), .ZN(\mult_19/ab[2][28] ) );
  NOR3_X1 U15091 ( .A1(n3297), .A2(n1936), .A3(n1090), .ZN(\mult_19/n4 ) );
  NOR2_X1 U15092 ( .A1(n3282), .A2(n3121), .ZN(\mult_19/ab[2][24] ) );
  NOR3_X1 U15093 ( .A1(n3285), .A2(n1936), .A3(n1040), .ZN(\mult_19/n8 ) );
  BUF_X1 U15094 ( .A(n1905), .Z(n3483) );
  BUF_X1 U15095 ( .A(n1908), .Z(n3297) );
  BUF_X1 U15096 ( .A(n1910), .Z(n3486) );
  BUF_X1 U15097 ( .A(n1907), .Z(n3462) );
  BUF_X1 U15098 ( .A(n1916), .Z(n3459) );
  BUF_X1 U15099 ( .A(n1966), .Z(n3456) );
  BUF_X1 U15100 ( .A(n1963), .Z(n3453) );
  BUF_X1 U15101 ( .A(n1967), .Z(n3450) );
  BUF_X1 U15102 ( .A(n1964), .Z(n3447) );
  BUF_X1 U15103 ( .A(n1968), .Z(n3444) );
  BUF_X1 U15104 ( .A(n1965), .Z(n3441) );
  BUF_X1 U15105 ( .A(n1937), .Z(n3438) );
  BUF_X1 U15106 ( .A(n1938), .Z(n3435) );
  BUF_X1 U15107 ( .A(n1939), .Z(n3432) );
  BUF_X1 U15108 ( .A(n1941), .Z(n3426) );
  BUF_X1 U15109 ( .A(n1911), .Z(n3300) );
  BUF_X1 U15110 ( .A(n1909), .Z(n3276) );
  BUF_X1 U15111 ( .A(n1922), .Z(n3273) );
  BUF_X1 U15112 ( .A(n1969), .Z(n3270) );
  BUF_X1 U15113 ( .A(n1970), .Z(n3267) );
  BUF_X1 U15114 ( .A(n1971), .Z(n3264) );
  BUF_X1 U15115 ( .A(n1972), .Z(n3261) );
  BUF_X1 U15116 ( .A(n1973), .Z(n3258) );
  BUF_X1 U15117 ( .A(n1974), .Z(n3255) );
  BUF_X1 U15118 ( .A(n1942), .Z(n3252) );
  BUF_X1 U15119 ( .A(n1943), .Z(n3249) );
  BUF_X1 U15120 ( .A(n1944), .Z(n3246) );
  BUF_X1 U15121 ( .A(n1946), .Z(n3240) );
  BUF_X1 U15122 ( .A(n1947), .Z(n3423) );
  BUF_X1 U15123 ( .A(n1948), .Z(n3420) );
  BUF_X1 U15124 ( .A(n1951), .Z(n3411) );
  BUF_X1 U15125 ( .A(n1940), .Z(n3429) );
  BUF_X1 U15126 ( .A(n1955), .Z(n3237) );
  BUF_X1 U15127 ( .A(n1956), .Z(n3234) );
  BUF_X1 U15128 ( .A(n1959), .Z(n3225) );
  BUF_X1 U15129 ( .A(n1945), .Z(n3243) );
  BUF_X1 U15130 ( .A(n1949), .Z(n3417) );
  BUF_X1 U15131 ( .A(n1950), .Z(n3414) );
  BUF_X1 U15132 ( .A(n1957), .Z(n3231) );
  BUF_X1 U15133 ( .A(n1958), .Z(n3228) );
  BUF_X1 U15134 ( .A(n1913), .Z(n3480) );
  BUF_X1 U15135 ( .A(n1912), .Z(n3477) );
  BUF_X1 U15136 ( .A(n1915), .Z(n3474) );
  BUF_X1 U15137 ( .A(n1914), .Z(n3471) );
  BUF_X1 U15138 ( .A(n1906), .Z(n3468) );
  BUF_X1 U15139 ( .A(n1917), .Z(n3294) );
  BUF_X1 U15140 ( .A(n1918), .Z(n3291) );
  BUF_X1 U15141 ( .A(n1920), .Z(n3288) );
  BUF_X1 U15142 ( .A(n1919), .Z(n3285) );
  BUF_X1 U15143 ( .A(n1921), .Z(n3282) );
  BUF_X1 U15144 ( .A(n1902), .Z(n3489) );
  BUF_X1 U15145 ( .A(n1903), .Z(n3303) );
  BUF_X1 U15146 ( .A(n1905), .Z(n3484) );
  BUF_X1 U15147 ( .A(n1908), .Z(n3298) );
  BUF_X1 U15148 ( .A(n1901), .Z(n3465) );
  BUF_X1 U15149 ( .A(n1904), .Z(n3279) );
  BUF_X1 U15150 ( .A(n1902), .Z(n3490) );
  BUF_X1 U15151 ( .A(n1903), .Z(n3304) );
  NOR2_X1 U15152 ( .A1(n3483), .A2(n3307), .ZN(\mult_20/ab[2][29] ) );
  NOR3_X1 U15153 ( .A1(n1034), .A2(n3517), .A3(n3483), .ZN(\mult_20/n3 ) );
  NOR2_X1 U15154 ( .A1(n3480), .A2(n3307), .ZN(\mult_20/ab[2][28] ) );
  NOR3_X1 U15155 ( .A1(n3483), .A2(n1935), .A3(n1029), .ZN(\mult_20/n4 ) );
  NOR2_X1 U15156 ( .A1(n3474), .A2(n3307), .ZN(\mult_20/ab[2][26] ) );
  NOR3_X1 U15157 ( .A1(n3477), .A2(n1935), .A3(n989), .ZN(\mult_20/n6 ) );
  NOR2_X1 U15158 ( .A1(n3468), .A2(n3307), .ZN(\mult_20/ab[2][24] ) );
  NOR3_X1 U15159 ( .A1(n3471), .A2(n1935), .A3(n979), .ZN(\mult_20/n8 ) );
  NOR2_X1 U15160 ( .A1(n3462), .A2(n3307), .ZN(\mult_20/ab[2][22] ) );
  NOR3_X1 U15161 ( .A1(n1025), .A2(n3522), .A3(n3462), .ZN(\mult_20/n10 ) );
  NOR2_X1 U15162 ( .A1(n3438), .A2(n3306), .ZN(\mult_20/ab[2][14] ) );
  NOR3_X1 U15163 ( .A1(n1008), .A2(n3520), .A3(n3438), .ZN(\mult_20/n18 ) );
  NOR2_X1 U15164 ( .A1(n3435), .A2(n3306), .ZN(\mult_20/ab[2][13] ) );
  NOR3_X1 U15165 ( .A1(n1006), .A2(n3520), .A3(n3435), .ZN(\mult_20/n19 ) );
  NOR2_X1 U15166 ( .A1(n3432), .A2(n3306), .ZN(\mult_20/ab[2][12] ) );
  NOR3_X1 U15167 ( .A1(n1004), .A2(n3520), .A3(n3432), .ZN(\mult_20/n20 ) );
  NOR2_X1 U15168 ( .A1(n3429), .A2(n3306), .ZN(\mult_20/ab[2][11] ) );
  NOR3_X1 U15169 ( .A1(n1002), .A2(n3520), .A3(n3429), .ZN(\mult_20/n21 ) );
  NOR2_X1 U15170 ( .A1(n3426), .A2(n3306), .ZN(\mult_20/ab[2][10] ) );
  NOR3_X1 U15171 ( .A1(n1000), .A2(n3519), .A3(n3426), .ZN(\mult_20/n22 ) );
  NOR2_X1 U15172 ( .A1(n3297), .A2(n3121), .ZN(\mult_19/ab[2][29] ) );
  NOR3_X1 U15173 ( .A1(n1095), .A2(n3528), .A3(n3297), .ZN(\mult_19/n3 ) );
  NOR2_X1 U15174 ( .A1(n3276), .A2(n3121), .ZN(\mult_19/ab[2][22] ) );
  NOR3_X1 U15175 ( .A1(n1086), .A2(n3533), .A3(n3276), .ZN(\mult_19/n10 ) );
  NOR2_X1 U15176 ( .A1(n3252), .A2(n3120), .ZN(\mult_19/ab[2][14] ) );
  NOR3_X1 U15177 ( .A1(n1069), .A2(n3531), .A3(n3252), .ZN(\mult_19/n18 ) );
  NOR2_X1 U15178 ( .A1(n3249), .A2(n3120), .ZN(\mult_19/ab[2][13] ) );
  NOR3_X1 U15179 ( .A1(n1067), .A2(n3531), .A3(n3249), .ZN(\mult_19/n19 ) );
  NOR2_X1 U15180 ( .A1(n3246), .A2(n3120), .ZN(\mult_19/ab[2][12] ) );
  NOR3_X1 U15181 ( .A1(n1065), .A2(n3531), .A3(n3246), .ZN(\mult_19/n20 ) );
  NOR2_X1 U15182 ( .A1(n3243), .A2(n3120), .ZN(\mult_19/ab[2][11] ) );
  NOR3_X1 U15183 ( .A1(n1063), .A2(n3531), .A3(n3243), .ZN(\mult_19/n21 ) );
  NOR2_X1 U15184 ( .A1(n3240), .A2(n3120), .ZN(\mult_19/ab[2][10] ) );
  NOR3_X1 U15185 ( .A1(n1061), .A2(n3530), .A3(n3240), .ZN(\mult_19/n22 ) );
  NOR2_X1 U15186 ( .A1(n3423), .A2(n3308), .ZN(\mult_20/ab[2][9] ) );
  NOR3_X1 U15187 ( .A1(n998), .A2(n3519), .A3(n3423), .ZN(\mult_20/n23 ) );
  NOR2_X1 U15188 ( .A1(n3420), .A2(n3308), .ZN(\mult_20/ab[2][8] ) );
  NOR3_X1 U15189 ( .A1(n996), .A2(n3519), .A3(n3420), .ZN(\mult_20/n24 ) );
  NOR2_X1 U15190 ( .A1(n3417), .A2(n3308), .ZN(\mult_20/ab[2][7] ) );
  NOR3_X1 U15191 ( .A1(n994), .A2(n3519), .A3(n3417), .ZN(\mult_20/n25 ) );
  NOR2_X1 U15192 ( .A1(n3414), .A2(n3308), .ZN(\mult_20/ab[2][6] ) );
  NOR3_X1 U15193 ( .A1(n992), .A2(n3518), .A3(n3414), .ZN(\mult_20/n26 ) );
  NOR2_X1 U15194 ( .A1(n3411), .A2(n3308), .ZN(\mult_20/ab[2][5] ) );
  NOR3_X1 U15195 ( .A1(n990), .A2(n3518), .A3(n3411), .ZN(\mult_20/n27 ) );
  NOR2_X1 U15196 ( .A1(n3222), .A2(n3122), .ZN(\mult_19/ab[2][4] ) );
  NOR3_X1 U15197 ( .A1(n1048), .A2(n3529), .A3(n3222), .ZN(\mult_19/n28 ) );
  NOR2_X1 U15198 ( .A1(n3219), .A2(n3122), .ZN(\mult_19/ab[2][3] ) );
  NOR3_X1 U15199 ( .A1(n1046), .A2(n3529), .A3(n3219), .ZN(\mult_19/n29 ) );
  NOR2_X1 U15200 ( .A1(n3216), .A2(n3121), .ZN(\mult_19/ab[2][2] ) );
  NOR3_X1 U15201 ( .A1(n1044), .A2(n3528), .A3(n3216), .ZN(\mult_19/n30 ) );
  NOR2_X1 U15202 ( .A1(n3213), .A2(n3120), .ZN(\mult_19/ab[2][1] ) );
  NOR3_X1 U15203 ( .A1(n1042), .A2(n3528), .A3(n3213), .ZN(\mult_19/n31 ) );
  NOR2_X1 U15204 ( .A1(n3237), .A2(n3122), .ZN(\mult_19/ab[2][9] ) );
  NOR3_X1 U15205 ( .A1(n1059), .A2(n3530), .A3(n3237), .ZN(\mult_19/n23 ) );
  NOR2_X1 U15206 ( .A1(n3234), .A2(n3122), .ZN(\mult_19/ab[2][8] ) );
  NOR3_X1 U15207 ( .A1(n1057), .A2(n3530), .A3(n3234), .ZN(\mult_19/n24 ) );
  NOR2_X1 U15208 ( .A1(n3231), .A2(n3122), .ZN(\mult_19/ab[2][7] ) );
  NOR3_X1 U15209 ( .A1(n1055), .A2(n3530), .A3(n3231), .ZN(\mult_19/n25 ) );
  NOR2_X1 U15210 ( .A1(n3228), .A2(n3122), .ZN(\mult_19/ab[2][6] ) );
  NOR3_X1 U15211 ( .A1(n1053), .A2(n3529), .A3(n3228), .ZN(\mult_19/n26 ) );
  NOR2_X1 U15212 ( .A1(n3225), .A2(n3122), .ZN(\mult_19/ab[2][5] ) );
  NOR3_X1 U15213 ( .A1(n1051), .A2(n3529), .A3(n3225), .ZN(\mult_19/n27 ) );
  NOR2_X1 U15214 ( .A1(n3408), .A2(n3308), .ZN(\mult_20/ab[2][4] ) );
  NOR3_X1 U15215 ( .A1(n987), .A2(n3518), .A3(n3408), .ZN(\mult_20/n28 ) );
  NOR2_X1 U15216 ( .A1(n3405), .A2(n3308), .ZN(\mult_20/ab[2][3] ) );
  NOR3_X1 U15217 ( .A1(n985), .A2(n3518), .A3(n3405), .ZN(\mult_20/n29 ) );
  NOR2_X1 U15218 ( .A1(n3402), .A2(n3307), .ZN(\mult_20/ab[2][2] ) );
  NOR3_X1 U15219 ( .A1(n983), .A2(n3517), .A3(n3402), .ZN(\mult_20/n30 ) );
  NOR2_X1 U15220 ( .A1(n3399), .A2(n3306), .ZN(\mult_20/ab[2][1] ) );
  NOR3_X1 U15221 ( .A1(n981), .A2(n3517), .A3(n3399), .ZN(\mult_20/n31 ) );
  BUF_X1 U15222 ( .A(n1926), .Z(n3122) );
  BUF_X1 U15223 ( .A(n1925), .Z(n3308) );
  BUF_X1 U15224 ( .A(n1924), .Z(n3125) );
  BUF_X1 U15225 ( .A(n1923), .Z(n3311) );
  BUF_X1 U15226 ( .A(n1993), .Z(n3128) );
  BUF_X1 U15227 ( .A(n1902), .Z(n3491) );
  BUF_X1 U15228 ( .A(n1903), .Z(n3305) );
  NOR2_X1 U15229 ( .A1(n3486), .A2(n3307), .ZN(\mult_20/ab[2][30] ) );
  NOR2_X1 U15230 ( .A1(n3523), .A2(n3489), .ZN(\mult_20/ab[1][31] ) );
  NOR3_X1 U15231 ( .A1(n1036), .A2(n3517), .A3(n3486), .ZN(\mult_20/n33 ) );
  NOR2_X1 U15232 ( .A1(n3300), .A2(n3121), .ZN(\mult_19/ab[2][30] ) );
  NOR2_X1 U15233 ( .A1(n3534), .A2(n3303), .ZN(\mult_19/ab[1][31] ) );
  NOR3_X1 U15234 ( .A1(n1097), .A2(n3528), .A3(n3300), .ZN(\mult_19/n33 ) );
  NOR2_X1 U15235 ( .A1(n3477), .A2(n3307), .ZN(\mult_20/ab[2][27] ) );
  NOR3_X1 U15236 ( .A1(n3480), .A2(n1935), .A3(n1010), .ZN(\mult_20/n5 ) );
  NOR2_X1 U15237 ( .A1(n3471), .A2(n3307), .ZN(\mult_20/ab[2][25] ) );
  NOR3_X1 U15238 ( .A1(n3474), .A2(n1935), .A3(n980), .ZN(\mult_20/n7 ) );
  NOR2_X1 U15239 ( .A1(n3459), .A2(n3307), .ZN(\mult_20/ab[2][21] ) );
  NOR3_X1 U15240 ( .A1(n1023), .A2(n3522), .A3(n3459), .ZN(\mult_20/n11 ) );
  NOR2_X1 U15241 ( .A1(n3453), .A2(n3306), .ZN(\mult_20/ab[2][19] ) );
  NOR3_X1 U15242 ( .A1(n1019), .A2(n3522), .A3(n3453), .ZN(\mult_20/n13 ) );
  NOR2_X1 U15243 ( .A1(n3447), .A2(n3306), .ZN(\mult_20/ab[2][17] ) );
  NOR3_X1 U15244 ( .A1(n1015), .A2(n3521), .A3(n3447), .ZN(\mult_20/n15 ) );
  NOR2_X1 U15245 ( .A1(n3441), .A2(n3306), .ZN(\mult_20/ab[2][15] ) );
  NOR3_X1 U15246 ( .A1(n1011), .A2(n3521), .A3(n3441), .ZN(\mult_20/n17 ) );
  NOR2_X1 U15247 ( .A1(n3291), .A2(n3121), .ZN(\mult_19/ab[2][27] ) );
  NOR3_X1 U15248 ( .A1(n3294), .A2(n1936), .A3(n1071), .ZN(\mult_19/n5 ) );
  NOR2_X1 U15249 ( .A1(n3288), .A2(n3121), .ZN(\mult_19/ab[2][26] ) );
  NOR3_X1 U15250 ( .A1(n3291), .A2(n1936), .A3(n1050), .ZN(\mult_19/n6 ) );
  NOR2_X1 U15251 ( .A1(n3285), .A2(n3121), .ZN(\mult_19/ab[2][25] ) );
  NOR3_X1 U15252 ( .A1(n3288), .A2(n1936), .A3(n1041), .ZN(\mult_19/n7 ) );
  NOR2_X1 U15253 ( .A1(n3279), .A2(n3121), .ZN(\mult_19/ab[2][23] ) );
  NOR3_X1 U15254 ( .A1(n3282), .A2(n1039), .A3(n1936), .ZN(\mult_19/n9 ) );
  NOR2_X1 U15255 ( .A1(n3456), .A2(n3307), .ZN(\mult_20/ab[2][20] ) );
  NOR3_X1 U15256 ( .A1(n1021), .A2(n3522), .A3(n3456), .ZN(\mult_20/n12 ) );
  NOR2_X1 U15257 ( .A1(n3450), .A2(n3306), .ZN(\mult_20/ab[2][18] ) );
  NOR3_X1 U15258 ( .A1(n1017), .A2(n3521), .A3(n3450), .ZN(\mult_20/n14 ) );
  NOR2_X1 U15259 ( .A1(n3444), .A2(n3306), .ZN(\mult_20/ab[2][16] ) );
  NOR3_X1 U15260 ( .A1(n1013), .A2(n3521), .A3(n3444), .ZN(\mult_20/n16 ) );
  NOR2_X1 U15261 ( .A1(n3273), .A2(n3121), .ZN(\mult_19/ab[2][21] ) );
  NOR3_X1 U15262 ( .A1(n1084), .A2(n3533), .A3(n3273), .ZN(\mult_19/n11 ) );
  NOR2_X1 U15263 ( .A1(n3270), .A2(n3121), .ZN(\mult_19/ab[2][20] ) );
  NOR3_X1 U15264 ( .A1(n1082), .A2(n3533), .A3(n3270), .ZN(\mult_19/n12 ) );
  NOR2_X1 U15265 ( .A1(n3267), .A2(n3120), .ZN(\mult_19/ab[2][19] ) );
  NOR3_X1 U15266 ( .A1(n1080), .A2(n3533), .A3(n3267), .ZN(\mult_19/n13 ) );
  NOR2_X1 U15267 ( .A1(n3264), .A2(n3120), .ZN(\mult_19/ab[2][18] ) );
  NOR3_X1 U15268 ( .A1(n1078), .A2(n3532), .A3(n3264), .ZN(\mult_19/n14 ) );
  NOR2_X1 U15269 ( .A1(n3261), .A2(n3120), .ZN(\mult_19/ab[2][17] ) );
  NOR3_X1 U15270 ( .A1(n1076), .A2(n3532), .A3(n3261), .ZN(\mult_19/n15 ) );
  NOR2_X1 U15271 ( .A1(n3258), .A2(n3120), .ZN(\mult_19/ab[2][16] ) );
  NOR3_X1 U15272 ( .A1(n1074), .A2(n3532), .A3(n3258), .ZN(\mult_19/n16 ) );
  NOR2_X1 U15273 ( .A1(n3255), .A2(n3120), .ZN(\mult_19/ab[2][15] ) );
  NOR3_X1 U15274 ( .A1(n1072), .A2(n3532), .A3(n3255), .ZN(\mult_19/n17 ) );
  BUF_X1 U15275 ( .A(n1807), .Z(n3522) );
  BUF_X1 U15276 ( .A(n1807), .Z(n3521) );
  BUF_X1 U15277 ( .A(n1807), .Z(n3520) );
  BUF_X1 U15278 ( .A(n1808), .Z(n3533) );
  BUF_X1 U15279 ( .A(n1808), .Z(n3532) );
  BUF_X1 U15280 ( .A(n1808), .Z(n3531) );
  BUF_X1 U15281 ( .A(n1807), .Z(n3519) );
  BUF_X1 U15282 ( .A(n1808), .Z(n3528) );
  BUF_X1 U15283 ( .A(n1808), .Z(n3530) );
  BUF_X1 U15284 ( .A(n1808), .Z(n3529) );
  BUF_X1 U15285 ( .A(n1807), .Z(n3518) );
  BUF_X1 U15286 ( .A(n1807), .Z(n3517) );
  BUF_X1 U15287 ( .A(n1807), .Z(n3523) );
  BUF_X1 U15288 ( .A(n1808), .Z(n3534) );
  BUF_X1 U15289 ( .A(n1931), .Z(n2996) );
  BUF_X1 U15290 ( .A(n1934), .Z(n3007) );
  BUF_X1 U15291 ( .A(n1932), .Z(n3002) );
  BUF_X1 U15292 ( .A(n1933), .Z(n3013) );
  BUF_X1 U15293 ( .A(n1934), .Z(n3008) );
  BUF_X1 U15294 ( .A(n1995), .Z(n3019) );
  BUF_X1 U15295 ( .A(n1997), .Z(n3025) );
  BUF_X1 U15296 ( .A(n1996), .Z(n3031) );
  BUF_X1 U15297 ( .A(n1933), .Z(n3014) );
  BUF_X1 U15298 ( .A(n1998), .Z(n3037) );
  BUF_X1 U15299 ( .A(n1995), .Z(n3020) );
  BUF_X1 U15300 ( .A(n1999), .Z(n3043) );
  BUF_X1 U15301 ( .A(n1997), .Z(n3026) );
  BUF_X1 U15302 ( .A(n1996), .Z(n3032) );
  BUF_X1 U15303 ( .A(n1930), .Z(n2991) );
  BUF_X1 U15304 ( .A(n1931), .Z(n2997) );
  BUF_X1 U15305 ( .A(n1998), .Z(n3038) );
  BUF_X1 U15306 ( .A(n1932), .Z(n3003) );
  BUF_X1 U15307 ( .A(n1934), .Z(n3009) );
  BUF_X1 U15308 ( .A(n1933), .Z(n3015) );
  BUF_X1 U15309 ( .A(n1995), .Z(n3021) );
  BUF_X1 U15310 ( .A(n1930), .Z(n2992) );
  BUF_X1 U15311 ( .A(n1997), .Z(n3027) );
  BUF_X1 U15312 ( .A(n1931), .Z(n2998) );
  BUF_X1 U15313 ( .A(n1996), .Z(n3033) );
  BUF_X1 U15314 ( .A(n1932), .Z(n3004) );
  BUF_X1 U15315 ( .A(n1934), .Z(n3010) );
  BUF_X1 U15316 ( .A(n1998), .Z(n3039) );
  BUF_X1 U15317 ( .A(n1933), .Z(n3016) );
  BUF_X1 U15318 ( .A(n1995), .Z(n3022) );
  BUF_X1 U15319 ( .A(n1997), .Z(n3028) );
  BUF_X1 U15320 ( .A(n1932), .Z(n3000) );
  BUF_X1 U15321 ( .A(n1934), .Z(n3006) );
  BUF_X1 U15322 ( .A(n1933), .Z(n3012) );
  BUF_X1 U15323 ( .A(n1996), .Z(n3034) );
  BUF_X1 U15324 ( .A(n1998), .Z(n3040) );
  BUF_X1 U15325 ( .A(n1995), .Z(n3018) );
  BUF_X1 U15326 ( .A(n1997), .Z(n3024) );
  BUF_X1 U15327 ( .A(n1996), .Z(n3030) );
  BUF_X1 U15328 ( .A(n1998), .Z(n3036) );
  BUF_X1 U15329 ( .A(n1999), .Z(n3042) );
  BUF_X1 U15330 ( .A(n2000), .Z(n3048) );
  BUF_X1 U15331 ( .A(n1991), .Z(n3312) );
  BUF_X1 U15332 ( .A(n1993), .Z(n3126) );
  BUF_X1 U15333 ( .A(n1992), .Z(n3315) );
  BUF_X1 U15334 ( .A(n1994), .Z(n3129) );
  BUF_X1 U15335 ( .A(n1979), .Z(n3319) );
  BUF_X1 U15336 ( .A(n1979), .Z(n3318) );
  BUF_X1 U15337 ( .A(n1985), .Z(n3133) );
  BUF_X1 U15338 ( .A(n1985), .Z(n3132) );
  BUF_X1 U15339 ( .A(n1980), .Z(n3322) );
  BUF_X1 U15340 ( .A(n1980), .Z(n3321) );
  BUF_X1 U15341 ( .A(n1986), .Z(n3136) );
  BUF_X1 U15342 ( .A(n1986), .Z(n3135) );
  BUF_X1 U15343 ( .A(n1981), .Z(n3325) );
  BUF_X1 U15344 ( .A(n1981), .Z(n3324) );
  BUF_X1 U15345 ( .A(n1987), .Z(n3139) );
  BUF_X1 U15346 ( .A(n1987), .Z(n3138) );
  BUF_X1 U15347 ( .A(n1982), .Z(n3328) );
  BUF_X1 U15348 ( .A(n1982), .Z(n3327) );
  BUF_X1 U15349 ( .A(n1988), .Z(n3142) );
  BUF_X1 U15350 ( .A(n1988), .Z(n3141) );
  BUF_X1 U15351 ( .A(n1983), .Z(n3331) );
  BUF_X1 U15352 ( .A(n1983), .Z(n3330) );
  BUF_X1 U15353 ( .A(n1989), .Z(n3145) );
  BUF_X1 U15354 ( .A(n1989), .Z(n3144) );
  BUF_X1 U15355 ( .A(n1984), .Z(n3334) );
  BUF_X1 U15356 ( .A(n1984), .Z(n3333) );
  BUF_X1 U15357 ( .A(n1990), .Z(n3148) );
  BUF_X1 U15358 ( .A(n1990), .Z(n3147) );
  BUF_X1 U15359 ( .A(n2004), .Z(n3336) );
  BUF_X1 U15360 ( .A(n2005), .Z(n3150) );
  BUF_X1 U15361 ( .A(n2006), .Z(n3339) );
  BUF_X1 U15362 ( .A(n2007), .Z(n3153) );
  BUF_X1 U15363 ( .A(n2004), .Z(n3337) );
  BUF_X1 U15364 ( .A(n2005), .Z(n3151) );
  BUF_X1 U15365 ( .A(n2006), .Z(n3340) );
  BUF_X1 U15366 ( .A(n2007), .Z(n3154) );
  BUF_X1 U15367 ( .A(n1975), .Z(n3399) );
  BUF_X1 U15368 ( .A(n1976), .Z(n3213) );
  BUF_X1 U15369 ( .A(n1952), .Z(n3222) );
  BUF_X1 U15370 ( .A(n1960), .Z(n3408) );
  BUF_X1 U15371 ( .A(n1961), .Z(n3405) );
  BUF_X1 U15372 ( .A(n1953), .Z(n3219) );
  BUF_X1 U15373 ( .A(n1954), .Z(n3216) );
  BUF_X1 U15374 ( .A(n1962), .Z(n3402) );
  BUF_X1 U15375 ( .A(n1977), .Z(n3397) );
  BUF_X1 U15376 ( .A(n1978), .Z(n3211) );
  NOR2_X1 U15377 ( .A1(n3397), .A2(n3306), .ZN(\mult_20/ab[2][0] ) );
  NOR3_X1 U15378 ( .A1(n1038), .A2(n1935), .A3(n3399), .ZN(\mult_20/n32 ) );
  NOR2_X1 U15379 ( .A1(n3211), .A2(n3120), .ZN(\mult_19/ab[2][0] ) );
  NOR3_X1 U15380 ( .A1(n1099), .A2(n1936), .A3(n3213), .ZN(\mult_19/n32 ) );
  BUF_X1 U15381 ( .A(n1991), .Z(n3314) );
  BUF_X1 U15382 ( .A(n1994), .Z(n3131) );
  BUF_X1 U15383 ( .A(n1992), .Z(n3317) );
  BUF_X1 U15384 ( .A(n1985), .Z(n3134) );
  BUF_X1 U15385 ( .A(n1979), .Z(n3320) );
  BUF_X1 U15386 ( .A(n1986), .Z(n3137) );
  BUF_X1 U15387 ( .A(n1980), .Z(n3323) );
  BUF_X1 U15388 ( .A(n1987), .Z(n3140) );
  BUF_X1 U15389 ( .A(n1981), .Z(n3326) );
  BUF_X1 U15390 ( .A(n1988), .Z(n3143) );
  BUF_X1 U15391 ( .A(n1982), .Z(n3329) );
  BUF_X1 U15392 ( .A(n1989), .Z(n3146) );
  BUF_X1 U15393 ( .A(n1983), .Z(n3332) );
  BUF_X1 U15394 ( .A(n1990), .Z(n3149) );
  BUF_X1 U15395 ( .A(n1984), .Z(n3335) );
  BUF_X1 U15396 ( .A(n1905), .Z(n3485) );
  BUF_X1 U15397 ( .A(n1908), .Z(n3299) );
  BUF_X1 U15398 ( .A(n1976), .Z(n3215) );
  BUF_X1 U15399 ( .A(n1975), .Z(n3401) );
  BUF_X1 U15400 ( .A(n1941), .Z(n3428) );
  BUF_X1 U15401 ( .A(n1946), .Z(n3242) );
  BUF_X1 U15402 ( .A(n1910), .Z(n3488) );
  BUF_X1 U15403 ( .A(n1913), .Z(n3482) );
  BUF_X1 U15404 ( .A(n1912), .Z(n3479) );
  BUF_X1 U15405 ( .A(n1915), .Z(n3476) );
  BUF_X1 U15406 ( .A(n1914), .Z(n3473) );
  BUF_X1 U15407 ( .A(n1906), .Z(n3470) );
  BUF_X1 U15408 ( .A(n1907), .Z(n3464) );
  BUF_X1 U15409 ( .A(n1916), .Z(n3461) );
  BUF_X1 U15410 ( .A(n1966), .Z(n3458) );
  BUF_X1 U15411 ( .A(n1963), .Z(n3455) );
  BUF_X1 U15412 ( .A(n1967), .Z(n3452) );
  BUF_X1 U15413 ( .A(n1964), .Z(n3449) );
  BUF_X1 U15414 ( .A(n1968), .Z(n3446) );
  BUF_X1 U15415 ( .A(n1965), .Z(n3443) );
  BUF_X1 U15416 ( .A(n1937), .Z(n3440) );
  BUF_X1 U15417 ( .A(n1938), .Z(n3437) );
  BUF_X1 U15418 ( .A(n1939), .Z(n3434) );
  BUF_X1 U15419 ( .A(n1940), .Z(n3431) );
  BUF_X1 U15420 ( .A(n1911), .Z(n3302) );
  BUF_X1 U15421 ( .A(n1917), .Z(n3296) );
  BUF_X1 U15422 ( .A(n1918), .Z(n3293) );
  BUF_X1 U15423 ( .A(n1920), .Z(n3290) );
  BUF_X1 U15424 ( .A(n1919), .Z(n3287) );
  BUF_X1 U15425 ( .A(n1921), .Z(n3284) );
  BUF_X1 U15426 ( .A(n1909), .Z(n3278) );
  BUF_X1 U15427 ( .A(n1922), .Z(n3275) );
  BUF_X1 U15428 ( .A(n1969), .Z(n3272) );
  BUF_X1 U15429 ( .A(n1970), .Z(n3269) );
  BUF_X1 U15430 ( .A(n1971), .Z(n3266) );
  BUF_X1 U15431 ( .A(n1972), .Z(n3263) );
  BUF_X1 U15432 ( .A(n1973), .Z(n3260) );
  BUF_X1 U15433 ( .A(n1974), .Z(n3257) );
  BUF_X1 U15434 ( .A(n1942), .Z(n3254) );
  BUF_X1 U15435 ( .A(n1943), .Z(n3251) );
  BUF_X1 U15436 ( .A(n1944), .Z(n3248) );
  BUF_X1 U15437 ( .A(n1945), .Z(n3245) );
  BUF_X1 U15438 ( .A(n1951), .Z(n3413) );
  BUF_X1 U15439 ( .A(n1959), .Z(n3227) );
  BUF_X1 U15440 ( .A(n1947), .Z(n3425) );
  BUF_X1 U15441 ( .A(n1948), .Z(n3422) );
  BUF_X1 U15442 ( .A(n1949), .Z(n3419) );
  BUF_X1 U15443 ( .A(n1950), .Z(n3416) );
  BUF_X1 U15444 ( .A(n1952), .Z(n3224) );
  BUF_X1 U15445 ( .A(n1953), .Z(n3221) );
  BUF_X1 U15446 ( .A(n1954), .Z(n3218) );
  BUF_X1 U15447 ( .A(n1955), .Z(n3239) );
  BUF_X1 U15448 ( .A(n1956), .Z(n3236) );
  BUF_X1 U15449 ( .A(n1957), .Z(n3233) );
  BUF_X1 U15450 ( .A(n1958), .Z(n3230) );
  BUF_X1 U15451 ( .A(n1960), .Z(n3410) );
  BUF_X1 U15452 ( .A(n1961), .Z(n3407) );
  BUF_X1 U15453 ( .A(n1962), .Z(n3404) );
  BUF_X1 U15454 ( .A(n1977), .Z(n3398) );
  BUF_X1 U15455 ( .A(n1978), .Z(n3212) );
  BUF_X1 U15456 ( .A(n1901), .Z(n3467) );
  BUF_X1 U15457 ( .A(n1904), .Z(n3281) );
  BUF_X1 U15458 ( .A(n2000), .Z(n3049) );
  BUF_X1 U15459 ( .A(n2001), .Z(n3055) );
  BUF_X1 U15460 ( .A(n2003), .Z(n3061) );
  BUF_X1 U15461 ( .A(n2002), .Z(n3067) );
  BUF_X1 U15462 ( .A(n1999), .Z(n3044) );
  BUF_X1 U15463 ( .A(n2021), .Z(n3073) );
  BUF_X1 U15464 ( .A(n2000), .Z(n3050) );
  BUF_X1 U15465 ( .A(n2020), .Z(n3079) );
  BUF_X1 U15466 ( .A(n2027), .Z(n3085) );
  BUF_X1 U15467 ( .A(n2026), .Z(n3091) );
  BUF_X1 U15468 ( .A(n2001), .Z(n3056) );
  BUF_X1 U15469 ( .A(n2003), .Z(n3062) );
  BUF_X1 U15470 ( .A(n2002), .Z(n3068) );
  BUF_X1 U15471 ( .A(n2021), .Z(n3074) );
  BUF_X1 U15472 ( .A(n2020), .Z(n3080) );
  BUF_X1 U15473 ( .A(n1999), .Z(n3045) );
  BUF_X1 U15474 ( .A(n2027), .Z(n3086) );
  BUF_X1 U15475 ( .A(n2000), .Z(n3051) );
  BUF_X1 U15476 ( .A(n2001), .Z(n3057) );
  BUF_X1 U15477 ( .A(n2003), .Z(n3063) );
  BUF_X1 U15478 ( .A(n2026), .Z(n3092) );
  BUF_X1 U15479 ( .A(n2002), .Z(n3069) );
  BUF_X1 U15480 ( .A(n2021), .Z(n3075) );
  BUF_X1 U15481 ( .A(n2020), .Z(n3081) );
  BUF_X1 U15482 ( .A(n1999), .Z(n3046) );
  BUF_X1 U15483 ( .A(n2000), .Z(n3052) );
  BUF_X1 U15484 ( .A(n2027), .Z(n3087) );
  BUF_X1 U15485 ( .A(n2001), .Z(n3054) );
  BUF_X1 U15486 ( .A(n2026), .Z(n3093) );
  BUF_X1 U15487 ( .A(n2003), .Z(n3060) );
  BUF_X1 U15488 ( .A(n2001), .Z(n3058) );
  BUF_X1 U15489 ( .A(n2002), .Z(n3066) );
  BUF_X1 U15490 ( .A(n2025), .Z(n3099) );
  BUF_X1 U15491 ( .A(n2003), .Z(n3064) );
  BUF_X1 U15492 ( .A(n2021), .Z(n3072) );
  BUF_X1 U15493 ( .A(n2020), .Z(n3078) );
  BUF_X1 U15494 ( .A(n2002), .Z(n3070) );
  BUF_X1 U15495 ( .A(n2021), .Z(n3076) );
  BUF_X1 U15496 ( .A(n2027), .Z(n3084) );
  BUF_X1 U15497 ( .A(n2020), .Z(n3082) );
  BUF_X1 U15498 ( .A(n2026), .Z(n3090) );
  BUF_X1 U15499 ( .A(n2027), .Z(n3088) );
  BUF_X1 U15500 ( .A(n2026), .Z(n3094) );
  BUF_X1 U15501 ( .A(n2025), .Z(n3100) );
  BUF_X1 U15502 ( .A(n2008), .Z(n3342) );
  BUF_X1 U15503 ( .A(n2009), .Z(n3156) );
  BUF_X1 U15504 ( .A(n2010), .Z(n3345) );
  BUF_X1 U15505 ( .A(n2011), .Z(n3159) );
  BUF_X1 U15506 ( .A(n2012), .Z(n3348) );
  BUF_X1 U15507 ( .A(n2013), .Z(n3162) );
  BUF_X1 U15508 ( .A(n2014), .Z(n3351) );
  BUF_X1 U15509 ( .A(n2015), .Z(n3165) );
  BUF_X1 U15510 ( .A(n2016), .Z(n3354) );
  BUF_X1 U15511 ( .A(n2008), .Z(n3343) );
  BUF_X1 U15512 ( .A(n2017), .Z(n3168) );
  BUF_X1 U15513 ( .A(n2009), .Z(n3157) );
  BUF_X1 U15514 ( .A(n2018), .Z(n3357) );
  BUF_X1 U15515 ( .A(n2019), .Z(n3171) );
  BUF_X1 U15516 ( .A(n2028), .Z(n3360) );
  BUF_X1 U15517 ( .A(n2010), .Z(n3346) );
  BUF_X1 U15518 ( .A(n2029), .Z(n3174) );
  BUF_X1 U15519 ( .A(n2011), .Z(n3160) );
  BUF_X1 U15520 ( .A(n2030), .Z(n3363) );
  BUF_X1 U15521 ( .A(n2031), .Z(n3177) );
  BUF_X1 U15522 ( .A(n2012), .Z(n3349) );
  BUF_X1 U15523 ( .A(n2013), .Z(n3163) );
  BUF_X1 U15524 ( .A(n2014), .Z(n3352) );
  BUF_X1 U15525 ( .A(n2015), .Z(n3166) );
  BUF_X1 U15526 ( .A(n2016), .Z(n3355) );
  BUF_X1 U15527 ( .A(n2017), .Z(n3169) );
  BUF_X1 U15528 ( .A(n2018), .Z(n3358) );
  BUF_X1 U15529 ( .A(n2019), .Z(n3172) );
  BUF_X1 U15530 ( .A(n2028), .Z(n3361) );
  BUF_X1 U15531 ( .A(n2029), .Z(n3175) );
  BUF_X1 U15532 ( .A(n1978), .Z(n3210) );
  BUF_X1 U15533 ( .A(n1977), .Z(n3396) );
  BUF_X1 U15534 ( .A(n1906), .Z(n3469) );
  BUF_X1 U15535 ( .A(n1901), .Z(n3466) );
  BUF_X1 U15536 ( .A(n1941), .Z(n3427) );
  BUF_X1 U15537 ( .A(n1921), .Z(n3283) );
  BUF_X1 U15538 ( .A(n1904), .Z(n3280) );
  BUF_X1 U15539 ( .A(n1946), .Z(n3241) );
  BUF_X1 U15540 ( .A(n1907), .Z(n3463) );
  BUF_X1 U15541 ( .A(n1916), .Z(n3460) );
  BUF_X1 U15542 ( .A(n1966), .Z(n3457) );
  BUF_X1 U15543 ( .A(n1963), .Z(n3454) );
  BUF_X1 U15544 ( .A(n1967), .Z(n3451) );
  BUF_X1 U15545 ( .A(n1964), .Z(n3448) );
  BUF_X1 U15546 ( .A(n1968), .Z(n3445) );
  BUF_X1 U15547 ( .A(n1965), .Z(n3442) );
  BUF_X1 U15548 ( .A(n1937), .Z(n3439) );
  BUF_X1 U15549 ( .A(n1938), .Z(n3436) );
  BUF_X1 U15550 ( .A(n1939), .Z(n3433) );
  BUF_X1 U15551 ( .A(n1940), .Z(n3430) );
  BUF_X1 U15552 ( .A(n1909), .Z(n3277) );
  BUF_X1 U15553 ( .A(n1922), .Z(n3274) );
  BUF_X1 U15554 ( .A(n1969), .Z(n3271) );
  BUF_X1 U15555 ( .A(n1970), .Z(n3268) );
  BUF_X1 U15556 ( .A(n1971), .Z(n3265) );
  BUF_X1 U15557 ( .A(n1972), .Z(n3262) );
  BUF_X1 U15558 ( .A(n1973), .Z(n3259) );
  BUF_X1 U15559 ( .A(n1974), .Z(n3256) );
  BUF_X1 U15560 ( .A(n1942), .Z(n3253) );
  BUF_X1 U15561 ( .A(n1943), .Z(n3250) );
  BUF_X1 U15562 ( .A(n1944), .Z(n3247) );
  BUF_X1 U15563 ( .A(n1945), .Z(n3244) );
  BUF_X1 U15564 ( .A(n1912), .Z(n3478) );
  BUF_X1 U15565 ( .A(n1918), .Z(n3292) );
  BUF_X1 U15566 ( .A(n1915), .Z(n3475) );
  BUF_X1 U15567 ( .A(n1914), .Z(n3472) );
  BUF_X1 U15568 ( .A(n1913), .Z(n3481) );
  BUF_X1 U15569 ( .A(n1920), .Z(n3289) );
  BUF_X1 U15570 ( .A(n1919), .Z(n3286) );
  BUF_X1 U15571 ( .A(n1917), .Z(n3295) );
  BUF_X1 U15572 ( .A(n1910), .Z(n3487) );
  BUF_X1 U15573 ( .A(n1911), .Z(n3301) );
  BUF_X1 U15574 ( .A(n1951), .Z(n3412) );
  BUF_X1 U15575 ( .A(n1959), .Z(n3226) );
  BUF_X1 U15576 ( .A(n1947), .Z(n3424) );
  BUF_X1 U15577 ( .A(n1948), .Z(n3421) );
  BUF_X1 U15578 ( .A(n1949), .Z(n3418) );
  BUF_X1 U15579 ( .A(n1950), .Z(n3415) );
  BUF_X1 U15580 ( .A(n1952), .Z(n3223) );
  BUF_X1 U15581 ( .A(n1953), .Z(n3220) );
  BUF_X1 U15582 ( .A(n1954), .Z(n3217) );
  BUF_X1 U15583 ( .A(n1976), .Z(n3214) );
  BUF_X1 U15584 ( .A(n1955), .Z(n3238) );
  BUF_X1 U15585 ( .A(n1956), .Z(n3235) );
  BUF_X1 U15586 ( .A(n1957), .Z(n3232) );
  BUF_X1 U15587 ( .A(n1958), .Z(n3229) );
  BUF_X1 U15588 ( .A(n1960), .Z(n3409) );
  BUF_X1 U15589 ( .A(n1961), .Z(n3406) );
  BUF_X1 U15590 ( .A(n1962), .Z(n3403) );
  BUF_X1 U15591 ( .A(n1975), .Z(n3400) );
  BUF_X1 U15592 ( .A(n2005), .Z(n3152) );
  BUF_X1 U15593 ( .A(n2004), .Z(n3338) );
  BUF_X1 U15594 ( .A(n2007), .Z(n3155) );
  BUF_X1 U15595 ( .A(n2006), .Z(n3341) );
  BUF_X1 U15596 ( .A(n2009), .Z(n3158) );
  BUF_X1 U15597 ( .A(n2008), .Z(n3344) );
  BUF_X1 U15598 ( .A(n2011), .Z(n3161) );
  BUF_X1 U15599 ( .A(n2010), .Z(n3347) );
  BUF_X1 U15600 ( .A(n2013), .Z(n3164) );
  BUF_X1 U15601 ( .A(n2012), .Z(n3350) );
  BUF_X1 U15602 ( .A(n2015), .Z(n3167) );
  BUF_X1 U15603 ( .A(n2014), .Z(n3353) );
  BUF_X1 U15604 ( .A(n2017), .Z(n3170) );
  BUF_X1 U15605 ( .A(n2016), .Z(n3356) );
  BUF_X1 U15606 ( .A(n2019), .Z(n3173) );
  BUF_X1 U15607 ( .A(n2018), .Z(n3359) );
  BUF_X1 U15608 ( .A(n2029), .Z(n3176) );
  BUF_X1 U15609 ( .A(n2028), .Z(n3362) );
  BUF_X1 U15610 ( .A(n2030), .Z(n3365) );
  BUF_X1 U15611 ( .A(n2025), .Z(n3097) );
  BUF_X1 U15612 ( .A(n2024), .Z(n3103) );
  BUF_X1 U15613 ( .A(n2023), .Z(n3109) );
  BUF_X1 U15614 ( .A(n2022), .Z(n3115) );
  BUF_X1 U15615 ( .A(n2025), .Z(n3098) );
  BUF_X1 U15616 ( .A(n2024), .Z(n3104) );
  BUF_X1 U15617 ( .A(n2023), .Z(n3110) );
  BUF_X1 U15618 ( .A(n2022), .Z(n3116) );
  BUF_X1 U15619 ( .A(n2024), .Z(n3105) );
  BUF_X1 U15620 ( .A(n2023), .Z(n3111) );
  BUF_X1 U15621 ( .A(n2022), .Z(n3117) );
  BUF_X1 U15622 ( .A(n2025), .Z(n3096) );
  BUF_X1 U15623 ( .A(n2024), .Z(n3102) );
  BUF_X1 U15624 ( .A(n2023), .Z(n3108) );
  BUF_X1 U15625 ( .A(n2022), .Z(n3114) );
  BUF_X1 U15626 ( .A(n2024), .Z(n3106) );
  BUF_X1 U15627 ( .A(n2023), .Z(n3112) );
  BUF_X1 U15628 ( .A(n2022), .Z(n3118) );
  BUF_X1 U15629 ( .A(n2032), .Z(n3366) );
  BUF_X1 U15630 ( .A(n2033), .Z(n3180) );
  BUF_X1 U15631 ( .A(n2034), .Z(n3369) );
  BUF_X1 U15632 ( .A(n2035), .Z(n3183) );
  BUF_X1 U15633 ( .A(n2036), .Z(n3372) );
  BUF_X1 U15634 ( .A(n2037), .Z(n3186) );
  BUF_X1 U15635 ( .A(n2038), .Z(n3375) );
  BUF_X1 U15636 ( .A(n2039), .Z(n3189) );
  BUF_X1 U15637 ( .A(n2040), .Z(n3378) );
  BUF_X1 U15638 ( .A(n2041), .Z(n3192) );
  BUF_X1 U15639 ( .A(n2042), .Z(n3381) );
  BUF_X1 U15640 ( .A(n2030), .Z(n3364) );
  BUF_X1 U15641 ( .A(n2043), .Z(n3195) );
  BUF_X1 U15642 ( .A(n2031), .Z(n3178) );
  BUF_X1 U15643 ( .A(n2032), .Z(n3367) );
  BUF_X1 U15644 ( .A(n2033), .Z(n3181) );
  BUF_X1 U15645 ( .A(n2046), .Z(n3384) );
  BUF_X1 U15646 ( .A(n2047), .Z(n3198) );
  BUF_X1 U15647 ( .A(n2034), .Z(n3370) );
  BUF_X1 U15648 ( .A(n2035), .Z(n3184) );
  BUF_X1 U15649 ( .A(n2036), .Z(n3373) );
  BUF_X1 U15650 ( .A(n2037), .Z(n3187) );
  BUF_X1 U15651 ( .A(n2038), .Z(n3376) );
  BUF_X1 U15652 ( .A(n2039), .Z(n3190) );
  BUF_X1 U15653 ( .A(n2040), .Z(n3379) );
  BUF_X1 U15654 ( .A(n2041), .Z(n3193) );
  BUF_X1 U15655 ( .A(n2042), .Z(n3382) );
  BUF_X1 U15656 ( .A(n2043), .Z(n3196) );
  BUF_X1 U15657 ( .A(n2047), .Z(n3199) );
  BUF_X1 U15658 ( .A(n2046), .Z(n3385) );
  BUF_X1 U15659 ( .A(n2048), .Z(n3388) );
  BUF_X1 U15660 ( .A(n2049), .Z(n3202) );
  BUF_X1 U15661 ( .A(n2031), .Z(n3179) );
  BUF_X1 U15662 ( .A(n2033), .Z(n3182) );
  BUF_X1 U15663 ( .A(n2032), .Z(n3368) );
  BUF_X1 U15664 ( .A(n2035), .Z(n3185) );
  BUF_X1 U15665 ( .A(n2034), .Z(n3371) );
  BUF_X1 U15666 ( .A(n2037), .Z(n3188) );
  BUF_X1 U15667 ( .A(n2036), .Z(n3374) );
  BUF_X1 U15668 ( .A(n2039), .Z(n3191) );
  BUF_X1 U15669 ( .A(n2038), .Z(n3377) );
  BUF_X1 U15670 ( .A(n2041), .Z(n3194) );
  BUF_X1 U15671 ( .A(n2040), .Z(n3380) );
  BUF_X1 U15672 ( .A(n2043), .Z(n3197) );
  BUF_X1 U15673 ( .A(n2042), .Z(n3383) );
  BUF_X1 U15674 ( .A(n2047), .Z(n3200) );
  BUF_X1 U15675 ( .A(n2046), .Z(n3386) );
  BUF_X1 U15676 ( .A(n2049), .Z(n3203) );
  BUF_X1 U15677 ( .A(n2048), .Z(n3389) );
  BUF_X1 U15678 ( .A(n2048), .Z(n3387) );
  BUF_X1 U15679 ( .A(n2049), .Z(n3201) );
  BUF_X1 U15680 ( .A(n2050), .Z(n3390) );
  BUF_X1 U15681 ( .A(n2051), .Z(n3204) );
  BUF_X1 U15682 ( .A(n2044), .Z(n3393) );
  BUF_X1 U15683 ( .A(n2045), .Z(n3207) );
  BUF_X1 U15684 ( .A(n2050), .Z(n3391) );
  BUF_X1 U15685 ( .A(n2051), .Z(n3205) );
  BUF_X1 U15686 ( .A(n2044), .Z(n3394) );
  BUF_X1 U15687 ( .A(n2045), .Z(n3208) );
  BUF_X1 U15688 ( .A(n2050), .Z(n3392) );
  BUF_X1 U15689 ( .A(n2051), .Z(n3206) );
  BUF_X1 U15690 ( .A(n2044), .Z(n3395) );
  BUF_X1 U15691 ( .A(n2045), .Z(n3209) );
  NOR2_X1 U15692 ( .A1(n1935), .A2(n3396), .ZN(N64) );
  NOR2_X1 U15693 ( .A1(n1936), .A2(n3210), .ZN(N0) );
  NOR2_X1 U15694 ( .A1(n2707), .A2(n2764), .ZN(\mult_22/ab[4][55] ) );
  NAND2_X1 U15695 ( .A1(reg_mid_0[3]), .A2(reg_mid_1[56]), .ZN(n935) );
  XNOR2_X1 U15696 ( .A(n2355), .B(n2356), .ZN(n941) );
  NAND2_X1 U15697 ( .A1(reg_mid_0[25]), .A2(reg_mid_1[35]), .ZN(n2355) );
  XNOR2_X1 U15698 ( .A(\mult_22/SUMB[24][36] ), .B(\mult_22/CARRYB[24][35] ), 
        .ZN(n2356) );
  OAI211_X1 U15699 ( .C1(\mult_22/CARRYB[24][35] ), .C2(\mult_22/SUMB[24][36] ), .A(reg_mid_1[35]), .B(reg_mid_0[25]), .ZN(n967) );
  OAI211_X1 U15700 ( .C1(\mult_22/CARRYB[2][56] ), .C2(\mult_22/SUMB[2][57] ), 
        .A(reg_mid_1[56]), .B(reg_mid_0[3]), .ZN(n961) );
  OAI211_X1 U15701 ( .C1(\mult_22/CARRYB[27][30] ), .C2(\mult_22/SUMB[27][31] ), .A(reg_mid_1[30]), .B(reg_mid_0[28]), .ZN(n963) );
  OAI211_X1 U15702 ( .C1(\mult_22/CARRYB[23][32] ), .C2(\mult_22/SUMB[23][33] ), .A(reg_mid_1[32]), .B(reg_mid_0[24]), .ZN(n968) );
  NAND2_X1 U15703 ( .A1(reg_mid_1[36]), .A2(n3495), .ZN(n814) );
  NAND2_X1 U15704 ( .A1(reg_mid_1[34]), .A2(n3492), .ZN(n810) );
  OAI211_X1 U15705 ( .C1(\mult_22/CARRYB[7][50] ), .C2(\mult_22/SUMB[7][51] ), 
        .A(reg_mid_1[50]), .B(reg_mid_0[8]), .ZN(n959) );
  NAND2_X1 U15706 ( .A1(reg_mid_1[38]), .A2(n3492), .ZN(n818) );
  NAND2_X1 U15707 ( .A1(reg_mid_1[32]), .A2(n3495), .ZN(n870) );
  NOR2_X1 U15708 ( .A1(n2648), .A2(n2811), .ZN(\mult_22/ab[12][45] ) );
  NOR2_X1 U15709 ( .A1(n2605), .A2(n2870), .ZN(\mult_22/ab[22][37] ) );
  NOR2_X1 U15710 ( .A1(n2545), .A2(n2941), .ZN(\mult_22/ab[34][27] ) );
  NOR2_X1 U15711 ( .A1(n2570), .A2(n2888), .ZN(\mult_22/ab[25][31] ) );
  NOR2_X1 U15712 ( .A1(n2677), .A2(n2793), .ZN(\mult_22/ab[9][49] ) );
  NAND2_X1 U15713 ( .A1(reg_mid_0[8]), .A2(reg_mid_1[50]), .ZN(n931) );
  NOR2_X1 U15714 ( .A1(n2557), .A2(n2911), .ZN(\mult_22/ab[29][29] ) );
  NAND2_X1 U15715 ( .A1(reg_mid_0[28]), .A2(reg_mid_1[30]), .ZN(n939) );
  NOR2_X1 U15716 ( .A1(n2370), .A2(n2770), .ZN(\mult_22/ab[5][54] ) );
  NOR2_X1 U15717 ( .A1(n2611), .A2(n2876), .ZN(\mult_22/ab[23][38] ) );
  NOR2_X1 U15718 ( .A1(n2370), .A2(n2776), .ZN(\mult_22/ab[6][54] ) );
  NOR2_X1 U15719 ( .A1(n2374), .A2(n2764), .ZN(\mult_22/ab[4][56] ) );
  OAI21_X1 U15720 ( .B1(n741), .B2(n740), .A(n961), .ZN(
        \mult_22/CARRYB[3][56] ) );
  NOR2_X1 U15721 ( .A1(n2370), .A2(n2788), .ZN(\mult_22/ab[8][54] ) );
  NOR2_X1 U15722 ( .A1(n2370), .A2(n2782), .ZN(\mult_22/ab[7][54] ) );
  NAND2_X1 U15723 ( .A1(reg_mid_1[41]), .A2(n2139), .ZN(n873) );
  NAND2_X1 U15724 ( .A1(reg_mid_1[39]), .A2(n2139), .ZN(n820) );
  NAND2_X1 U15725 ( .A1(reg_mid_1[37]), .A2(n2139), .ZN(n816) );
  NAND2_X1 U15726 ( .A1(reg_mid_1[35]), .A2(n3495), .ZN(n812) );
  AND2_X1 U15727 ( .A1(reg_mid_0[4]), .A2(reg_mid_1[52]), .ZN(n2357) );
  XNOR2_X1 U15728 ( .A(n956), .B(n2358), .ZN(\mult_22/SUMB[18][40] ) );
  AND2_X1 U15729 ( .A1(reg_mid_0[18]), .A2(reg_mid_1[40]), .ZN(n2358) );
  NOR2_X1 U15730 ( .A1(n2599), .A2(n2870), .ZN(\mult_22/ab[22][36] ) );
  OAI21_X1 U15731 ( .B1(n975), .B2(n713), .A(n953), .ZN(
        \mult_22/CARRYB[21][36] ) );
  AOI21_X1 U15732 ( .B1(reg_mid_0[21]), .B2(reg_mid_1[36]), .A(
        \mult_22/CARRYB[20][36] ), .ZN(n975) );
  NOR2_X1 U15733 ( .A1(n2370), .A2(n2794), .ZN(\mult_22/ab[9][54] ) );
  INV_X1 U15734 ( .A(reg_mid_1[55]), .ZN(n753) );
  NAND2_X1 U15735 ( .A1(reg_mid_1[38]), .A2(n3502), .ZN(n821) );
  INV_X1 U15736 ( .A(reg_mid_1[62]), .ZN(n746) );
  INV_X1 U15737 ( .A(reg_mid_1[60]), .ZN(n748) );
  OR2_X1 U15738 ( .A1(n2359), .A2(n3498), .ZN(n914) );
  INV_X1 U15739 ( .A(reg_mid_1[54]), .ZN(n754) );
  NAND2_X1 U15740 ( .A1(reg_mid_1[44]), .A2(n2371), .ZN(n918) );
  NAND2_X1 U15741 ( .A1(reg_mid_1[42]), .A2(n3492), .ZN(n916) );
  NAND2_X1 U15742 ( .A1(reg_mid_1[42]), .A2(n3502), .ZN(n825) );
  NAND2_X1 U15743 ( .A1(reg_mid_1[36]), .A2(n3502), .ZN(n817) );
  NAND2_X1 U15744 ( .A1(reg_mid_1[35]), .A2(n3502), .ZN(n815) );
  OR2_X1 U15745 ( .A1(n2360), .A2(n3499), .ZN(n878) );
  NAND2_X1 U15746 ( .A1(reg_mid_1[46]), .A2(n3493), .ZN(n917) );
  OR2_X1 U15747 ( .A1(n2361), .A2(n3511), .ZN(n879) );
  OR2_X1 U15748 ( .A1(n2362), .A2(n3511), .ZN(n875) );
  OR2_X1 U15749 ( .A1(n2363), .A2(n3511), .ZN(n892) );
  NAND2_X1 U15750 ( .A1(reg_mid_1[47]), .A2(n3494), .ZN(n915) );
  OR2_X1 U15751 ( .A1(n2372), .A2(n2142), .ZN(n2364) );
  INV_X1 U15752 ( .A(reg_mid_1[56]), .ZN(n752) );
  NAND2_X1 U15753 ( .A1(reg_mid_1[21]), .A2(n3495), .ZN(n852) );
  NAND2_X1 U15754 ( .A1(reg_mid_1[17]), .A2(n3492), .ZN(n845) );
  NAND2_X1 U15755 ( .A1(reg_mid_1[14]), .A2(n2139), .ZN(n841) );
  NAND2_X1 U15756 ( .A1(reg_mid_1[24]), .A2(n3492), .ZN(n858) );
  NAND2_X1 U15757 ( .A1(reg_mid_1[23]), .A2(n2139), .ZN(n856) );
  NAND2_X1 U15758 ( .A1(reg_mid_1[19]), .A2(n2371), .ZN(n849) );
  NAND2_X1 U15759 ( .A1(reg_mid_1[16]), .A2(n3492), .ZN(n843) );
  NAND2_X1 U15760 ( .A1(reg_mid_1[8]), .A2(n3492), .ZN(n835) );
  NAND2_X1 U15761 ( .A1(reg_mid_1[22]), .A2(n3495), .ZN(n854) );
  NAND2_X1 U15762 ( .A1(reg_mid_1[10]), .A2(n2371), .ZN(n839) );
  NAND2_X1 U15763 ( .A1(reg_mid_1[28]), .A2(n3502), .ZN(n899) );
  NAND2_X1 U15764 ( .A1(reg_mid_1[12]), .A2(n3502), .ZN(n894) );
  NAND2_X1 U15765 ( .A1(reg_mid_1[0]), .A2(n3501), .ZN(n907) );
  NAND2_X1 U15766 ( .A1(reg_mid_1[12]), .A2(n3495), .ZN(n921) );
  NAND2_X1 U15767 ( .A1(reg_mid_1[11]), .A2(n2139), .ZN(n920) );
  NAND2_X1 U15768 ( .A1(reg_mid_1[26]), .A2(n3502), .ZN(n897) );
  NAND2_X1 U15769 ( .A1(reg_mid_1[24]), .A2(n3500), .ZN(n895) );
  NAND2_X1 U15770 ( .A1(reg_mid_1[18]), .A2(n3494), .ZN(n847) );
  NAND2_X1 U15771 ( .A1(reg_mid_1[6]), .A2(n3493), .ZN(n833) );
  NAND2_X1 U15772 ( .A1(reg_mid_1[9]), .A2(n3494), .ZN(n837) );
  NAND2_X1 U15773 ( .A1(reg_mid_1[2]), .A2(n2371), .ZN(n831) );
  NAND2_X1 U15774 ( .A1(reg_mid_1[23]), .A2(n3502), .ZN(n859) );
  NAND2_X1 U15775 ( .A1(reg_mid_1[22]), .A2(n3502), .ZN(n857) );
  NAND2_X1 U15776 ( .A1(reg_mid_1[16]), .A2(n3502), .ZN(n846) );
  NAND2_X1 U15777 ( .A1(reg_mid_1[7]), .A2(n3502), .ZN(n836) );
  NAND2_X1 U15778 ( .A1(reg_mid_1[18]), .A2(n3501), .ZN(n850) );
  NAND2_X1 U15779 ( .A1(reg_mid_1[13]), .A2(n3500), .ZN(n842) );
  NAND2_X1 U15780 ( .A1(reg_mid_1[9]), .A2(n3502), .ZN(n840) );
  NAND2_X1 U15781 ( .A1(reg_mid_1[5]), .A2(n2188), .ZN(n834) );
  NAND2_X1 U15782 ( .A1(reg_mid_1[13]), .A2(n3493), .ZN(n922) );
  NAND2_X1 U15783 ( .A1(reg_mid_1[5]), .A2(n3495), .ZN(n919) );
  NOR2_X1 U15784 ( .A1(n2370), .A2(n3088), .ZN(\mult_22/ab[58][54] ) );
  NOR2_X1 U15785 ( .A1(n2370), .A2(n3094), .ZN(\mult_22/ab[59][54] ) );
  NOR2_X1 U15786 ( .A1(n2370), .A2(n3100), .ZN(\mult_22/ab[60][54] ) );
  NOR2_X1 U15787 ( .A1(n2370), .A2(n3106), .ZN(\mult_22/ab[61][54] ) );
  NOR2_X1 U15788 ( .A1(n2370), .A2(n3112), .ZN(\mult_22/ab[62][54] ) );
  NAND2_X1 U15789 ( .A1(reg_mid_0[23]), .A2(reg_mid_1[37]), .ZN(n948) );
  NAND2_X1 U15790 ( .A1(n3515), .A2(reg_ini_3[23]), .ZN(n1025) );
  NAND2_X1 U15791 ( .A1(n3526), .A2(reg_ini_1[23]), .ZN(n1086) );
  NAND2_X1 U15792 ( .A1(reg_ini_3[22]), .A2(n3515), .ZN(n1023) );
  NAND2_X1 U15793 ( .A1(reg_ini_3[21]), .A2(n3515), .ZN(n1021) );
  NAND2_X1 U15794 ( .A1(reg_ini_3[20]), .A2(n3515), .ZN(n1019) );
  NAND2_X1 U15795 ( .A1(reg_ini_3[19]), .A2(n3515), .ZN(n1017) );
  NAND2_X1 U15796 ( .A1(reg_ini_3[18]), .A2(n3515), .ZN(n1015) );
  NAND2_X1 U15797 ( .A1(reg_ini_3[17]), .A2(n3515), .ZN(n1013) );
  NAND2_X1 U15798 ( .A1(reg_ini_1[22]), .A2(n3526), .ZN(n1084) );
  NAND2_X1 U15799 ( .A1(reg_ini_1[21]), .A2(n3526), .ZN(n1082) );
  NAND2_X1 U15800 ( .A1(reg_ini_1[20]), .A2(n3526), .ZN(n1080) );
  NAND2_X1 U15801 ( .A1(reg_ini_1[19]), .A2(n3526), .ZN(n1078) );
  NAND2_X1 U15802 ( .A1(reg_ini_1[18]), .A2(n3526), .ZN(n1076) );
  NAND2_X1 U15803 ( .A1(reg_ini_1[17]), .A2(n3526), .ZN(n1074) );
  NAND2_X1 U15804 ( .A1(reg_ini_3[31]), .A2(n3513), .ZN(n1036) );
  NAND2_X1 U15805 ( .A1(reg_ini_3[30]), .A2(n3513), .ZN(n1034) );
  NAND2_X1 U15806 ( .A1(reg_ini_3[16]), .A2(n3514), .ZN(n1011) );
  NAND2_X1 U15807 ( .A1(reg_ini_3[15]), .A2(n3514), .ZN(n1008) );
  NAND2_X1 U15808 ( .A1(reg_ini_3[14]), .A2(n3514), .ZN(n1006) );
  NAND2_X1 U15809 ( .A1(reg_ini_3[13]), .A2(n3514), .ZN(n1004) );
  NAND2_X1 U15810 ( .A1(reg_ini_3[12]), .A2(n3514), .ZN(n1002) );
  NAND2_X1 U15811 ( .A1(reg_ini_1[31]), .A2(n3524), .ZN(n1097) );
  NAND2_X1 U15812 ( .A1(reg_ini_1[30]), .A2(n3524), .ZN(n1095) );
  NAND2_X1 U15813 ( .A1(reg_ini_1[16]), .A2(n3525), .ZN(n1072) );
  NAND2_X1 U15814 ( .A1(reg_ini_1[15]), .A2(n3525), .ZN(n1069) );
  NAND2_X1 U15815 ( .A1(reg_ini_1[14]), .A2(n3525), .ZN(n1067) );
  NAND2_X1 U15816 ( .A1(reg_ini_1[13]), .A2(n3525), .ZN(n1065) );
  NAND2_X1 U15817 ( .A1(reg_ini_1[12]), .A2(n3525), .ZN(n1063) );
  NAND2_X1 U15818 ( .A1(reg_ini_3[11]), .A2(n3514), .ZN(n1000) );
  NAND2_X1 U15819 ( .A1(reg_ini_3[10]), .A2(n3514), .ZN(n998) );
  NAND2_X1 U15820 ( .A1(reg_ini_3[9]), .A2(n3514), .ZN(n996) );
  NAND2_X1 U15821 ( .A1(reg_ini_3[8]), .A2(n3514), .ZN(n994) );
  NAND2_X1 U15822 ( .A1(reg_ini_3[7]), .A2(n3514), .ZN(n992) );
  NAND2_X1 U15823 ( .A1(reg_ini_1[5]), .A2(n3524), .ZN(n1048) );
  NAND2_X1 U15824 ( .A1(reg_ini_1[4]), .A2(n3524), .ZN(n1046) );
  NAND2_X1 U15825 ( .A1(reg_ini_1[11]), .A2(n3525), .ZN(n1061) );
  NAND2_X1 U15826 ( .A1(reg_ini_1[10]), .A2(n3525), .ZN(n1059) );
  NAND2_X1 U15827 ( .A1(reg_ini_1[9]), .A2(n3525), .ZN(n1057) );
  NAND2_X1 U15828 ( .A1(reg_ini_1[8]), .A2(n3525), .ZN(n1055) );
  NAND2_X1 U15829 ( .A1(reg_ini_1[7]), .A2(n3525), .ZN(n1053) );
  NAND2_X1 U15830 ( .A1(reg_ini_1[6]), .A2(n3525), .ZN(n1051) );
  NAND2_X1 U15831 ( .A1(reg_ini_3[6]), .A2(n3514), .ZN(n990) );
  NAND2_X1 U15832 ( .A1(reg_ini_3[5]), .A2(n3513), .ZN(n987) );
  NAND2_X1 U15833 ( .A1(reg_ini_3[4]), .A2(n3513), .ZN(n985) );
  NAND2_X1 U15834 ( .A1(reg_ini_3[28]), .A2(n1806), .ZN(n1029) );
  NAND2_X1 U15835 ( .A1(reg_ini_3[27]), .A2(n1806), .ZN(n1010) );
  NAND2_X1 U15836 ( .A1(reg_ini_3[26]), .A2(n1806), .ZN(n989) );
  NAND2_X1 U15837 ( .A1(reg_ini_3[25]), .A2(n1806), .ZN(n980) );
  NAND2_X1 U15838 ( .A1(reg_ini_3[24]), .A2(n1806), .ZN(n979) );
  NAND2_X1 U15839 ( .A1(reg_ini_1[28]), .A2(n1805), .ZN(n1090) );
  NAND2_X1 U15840 ( .A1(reg_ini_1[27]), .A2(n1805), .ZN(n1071) );
  NAND2_X1 U15841 ( .A1(reg_ini_1[26]), .A2(n1805), .ZN(n1050) );
  NAND2_X1 U15842 ( .A1(reg_ini_1[25]), .A2(n1805), .ZN(n1041) );
  NAND2_X1 U15843 ( .A1(reg_ini_1[24]), .A2(n1805), .ZN(n1040) );
  NAND2_X1 U15844 ( .A1(reg_ini_3[23]), .A2(n1806), .ZN(n978) );
  NAND2_X1 U15845 ( .A1(reg_ini_1[23]), .A2(n1805), .ZN(n1039) );
  NAND2_X1 U15846 ( .A1(reg_ini_3[7]), .A2(n3516), .ZN(n995) );
  NAND2_X1 U15847 ( .A1(reg_ini_3[6]), .A2(n3516), .ZN(n993) );
  NAND2_X1 U15848 ( .A1(reg_ini_1[5]), .A2(n3527), .ZN(n1052) );
  NAND2_X1 U15849 ( .A1(reg_ini_1[4]), .A2(n3527), .ZN(n1049) );
  NAND2_X1 U15850 ( .A1(reg_ini_1[3]), .A2(n3527), .ZN(n1047) );
  NAND2_X1 U15851 ( .A1(reg_ini_1[2]), .A2(n3527), .ZN(n1045) );
  NAND2_X1 U15852 ( .A1(reg_ini_1[7]), .A2(n3527), .ZN(n1056) );
  NAND2_X1 U15853 ( .A1(reg_ini_1[6]), .A2(n3527), .ZN(n1054) );
  NAND2_X1 U15854 ( .A1(reg_ini_3[5]), .A2(n3516), .ZN(n991) );
  NAND2_X1 U15855 ( .A1(reg_ini_3[4]), .A2(n3516), .ZN(n988) );
  NAND2_X1 U15856 ( .A1(reg_ini_3[3]), .A2(n3516), .ZN(n986) );
  NAND2_X1 U15857 ( .A1(reg_ini_3[2]), .A2(n3516), .ZN(n984) );
  NAND2_X1 U15858 ( .A1(reg_ini_3[29]), .A2(n3513), .ZN(n1033) );
  NAND2_X1 U15859 ( .A1(reg_ini_3[28]), .A2(n3513), .ZN(n1032) );
  NAND2_X1 U15860 ( .A1(reg_ini_3[27]), .A2(n3513), .ZN(n1031) );
  NAND2_X1 U15861 ( .A1(reg_ini_3[26]), .A2(n3513), .ZN(n1030) );
  NAND2_X1 U15862 ( .A1(reg_ini_3[25]), .A2(n3513), .ZN(n1028) );
  NAND2_X1 U15863 ( .A1(reg_ini_3[24]), .A2(n3514), .ZN(n1027) );
  NAND2_X1 U15864 ( .A1(reg_ini_1[29]), .A2(n3524), .ZN(n1094) );
  NAND2_X1 U15865 ( .A1(reg_ini_1[28]), .A2(n3524), .ZN(n1093) );
  NAND2_X1 U15866 ( .A1(reg_ini_1[27]), .A2(n3524), .ZN(n1092) );
  NAND2_X1 U15867 ( .A1(reg_ini_1[26]), .A2(n3524), .ZN(n1091) );
  NAND2_X1 U15868 ( .A1(reg_ini_1[25]), .A2(n3524), .ZN(n1089) );
  NAND2_X1 U15869 ( .A1(reg_ini_1[24]), .A2(n3525), .ZN(n1088) );
  NAND2_X1 U15870 ( .A1(reg_ini_3[30]), .A2(n1806), .ZN(n1037) );
  NAND2_X1 U15871 ( .A1(reg_ini_3[29]), .A2(n1806), .ZN(n1035) );
  NAND2_X1 U15872 ( .A1(reg_ini_3[22]), .A2(n1806), .ZN(n1026) );
  NAND2_X1 U15873 ( .A1(reg_ini_3[21]), .A2(n1806), .ZN(n1024) );
  NAND2_X1 U15874 ( .A1(reg_ini_3[20]), .A2(n3516), .ZN(n1022) );
  NAND2_X1 U15875 ( .A1(reg_ini_3[19]), .A2(n3516), .ZN(n1020) );
  NAND2_X1 U15876 ( .A1(reg_ini_3[18]), .A2(n3516), .ZN(n1018) );
  NAND2_X1 U15877 ( .A1(reg_ini_3[17]), .A2(n3516), .ZN(n1016) );
  NAND2_X1 U15878 ( .A1(reg_ini_3[16]), .A2(n3516), .ZN(n1014) );
  NAND2_X1 U15879 ( .A1(reg_ini_3[15]), .A2(n3516), .ZN(n1012) );
  NAND2_X1 U15880 ( .A1(reg_ini_3[14]), .A2(n3516), .ZN(n1009) );
  NAND2_X1 U15881 ( .A1(reg_ini_3[13]), .A2(n3516), .ZN(n1007) );
  NAND2_X1 U15882 ( .A1(reg_ini_3[12]), .A2(n3516), .ZN(n1005) );
  NAND2_X1 U15883 ( .A1(reg_ini_3[11]), .A2(n3516), .ZN(n1003) );
  NAND2_X1 U15884 ( .A1(reg_ini_1[30]), .A2(n1805), .ZN(n1098) );
  NAND2_X1 U15885 ( .A1(reg_ini_1[29]), .A2(n1805), .ZN(n1096) );
  NAND2_X1 U15886 ( .A1(reg_ini_1[22]), .A2(n1805), .ZN(n1087) );
  NAND2_X1 U15887 ( .A1(reg_ini_1[21]), .A2(n1805), .ZN(n1085) );
  NAND2_X1 U15888 ( .A1(reg_ini_1[20]), .A2(n3527), .ZN(n1083) );
  NAND2_X1 U15889 ( .A1(reg_ini_1[19]), .A2(n3527), .ZN(n1081) );
  NAND2_X1 U15890 ( .A1(reg_ini_1[18]), .A2(n3527), .ZN(n1079) );
  NAND2_X1 U15891 ( .A1(reg_ini_1[17]), .A2(n3527), .ZN(n1077) );
  NAND2_X1 U15892 ( .A1(reg_ini_1[16]), .A2(n3527), .ZN(n1075) );
  NAND2_X1 U15893 ( .A1(reg_ini_1[15]), .A2(n3527), .ZN(n1073) );
  NAND2_X1 U15894 ( .A1(reg_ini_1[14]), .A2(n3527), .ZN(n1070) );
  NAND2_X1 U15895 ( .A1(reg_ini_1[13]), .A2(n3527), .ZN(n1068) );
  NAND2_X1 U15896 ( .A1(reg_ini_1[12]), .A2(n3527), .ZN(n1066) );
  NAND2_X1 U15897 ( .A1(reg_ini_1[11]), .A2(n3527), .ZN(n1064) );
  NAND2_X1 U15898 ( .A1(reg_ini_3[10]), .A2(n3516), .ZN(n1001) );
  NAND2_X1 U15899 ( .A1(reg_ini_3[9]), .A2(n3516), .ZN(n999) );
  NAND2_X1 U15900 ( .A1(reg_ini_3[8]), .A2(n3516), .ZN(n997) );
  NAND2_X1 U15901 ( .A1(reg_ini_1[10]), .A2(n3527), .ZN(n1062) );
  NAND2_X1 U15902 ( .A1(reg_ini_1[9]), .A2(n3527), .ZN(n1060) );
  NAND2_X1 U15903 ( .A1(reg_ini_1[8]), .A2(n3527), .ZN(n1058) );
  NAND2_X1 U15904 ( .A1(reg_ini_1[3]), .A2(n3524), .ZN(n1044) );
  NAND2_X1 U15905 ( .A1(reg_ini_3[3]), .A2(n3513), .ZN(n983) );
  NAND2_X1 U15906 ( .A1(reg_ini_3[2]), .A2(n3513), .ZN(n981) );
  NAND2_X1 U15907 ( .A1(reg_ini_1[2]), .A2(n3524), .ZN(n1042) );
  NAND2_X1 U15908 ( .A1(reg_ini_1[0]), .A2(n3527), .ZN(n1099) );
  NAND2_X1 U15909 ( .A1(reg_ini_3[0]), .A2(n3516), .ZN(n1038) );
  NAND2_X1 U15910 ( .A1(reg_ini_3[1]), .A2(n3516), .ZN(n982) );
  NAND2_X1 U15911 ( .A1(reg_ini_1[1]), .A2(n3527), .ZN(n1043) );
  NAND2_X1 U15912 ( .A1(reg_ini_3[1]), .A2(n3513), .ZN(n1108) );
  NAND2_X1 U15913 ( .A1(reg_ini_1[1]), .A2(n3524), .ZN(n1799) );
  NAND2_X1 U15914 ( .A1(reg_ini_2[31]), .A2(reg_ini_3[31]), .ZN(n1637) );
  NAND2_X1 U15915 ( .A1(reg_ini_0[31]), .A2(reg_ini_1[31]), .ZN(n1111) );
  NAND2_X1 U15916 ( .A1(reg_mid_0[63]), .A2(reg_mid_1[63]), .ZN(n1288) );
  NAND2_X1 U15917 ( .A1(n594), .A2(n2169), .ZN(n1631) );
  AOI21_X1 U15918 ( .B1(n2087), .B2(n590), .A(n591), .ZN(n1532) );
  XNOR2_X1 U15919 ( .A(n1282), .B(n1281), .ZN(N255) );
  CLKBUF_X1 U15920 ( .A(n1471), .Z(n2365) );
  CLKBUF_X1 U15921 ( .A(n1809), .Z(n2367) );
  CLKBUF_X1 U15922 ( .A(n1809), .Z(n2698) );
  NOR2_X1 U15923 ( .A1(n3497), .A2(n2380), .ZN(N128) );
  NOR3_X1 U15924 ( .A1(n890), .A2(n3497), .A3(n2410), .ZN(\mult_22/n55 ) );
  NOR3_X1 U15925 ( .A1(n2452), .A2(n3499), .A3(n893), .ZN(\mult_22/n49 ) );
  NOR3_X1 U15926 ( .A1(n2530), .A2(n3499), .A3(n895), .ZN(\mult_22/n38 ) );
  NOR3_X1 U15927 ( .A1(n2542), .A2(n3497), .A3(n897), .ZN(\mult_22/n36 ) );
  NOR3_X1 U15928 ( .A1(n2548), .A2(n3497), .A3(n898), .ZN(\mult_22/n35 ) );
  NOR3_X1 U15929 ( .A1(n2560), .A2(n3497), .A3(n900), .ZN(\mult_22/n33 ) );
  NOR3_X1 U15930 ( .A1(n905), .A2(n3497), .A3(n2566), .ZN(\mult_22/n32 ) );
  NOR3_X1 U15931 ( .A1(n906), .A2(n3497), .A3(n2577), .ZN(\mult_22/n31 ) );
  NOR3_X1 U15932 ( .A1(n888), .A2(n3497), .A3(n2630), .ZN(\mult_22/n58 ) );
  NAND2_X1 U15933 ( .A1(reg_mid_1[1]), .A2(n3500), .ZN(n832) );
  NAND2_X1 U15934 ( .A1(reg_mid_1[8]), .A2(n3500), .ZN(n838) );
  NAND2_X1 U15935 ( .A1(reg_mid_1[11]), .A2(n3500), .ZN(n893) );
  NAND2_X1 U15936 ( .A1(reg_mid_1[20]), .A2(n3500), .ZN(n853) );
  NAND2_X1 U15937 ( .A1(reg_mid_1[25]), .A2(n3500), .ZN(n896) );
  NAND2_X1 U15938 ( .A1(reg_mid_1[29]), .A2(n3500), .ZN(n900) );
  NAND2_X1 U15939 ( .A1(reg_mid_1[44]), .A2(n3500), .ZN(n827) );
  NOR2_X1 U15940 ( .A1(n2698), .A2(n2157), .ZN(\mult_22/ab[2][53] ) );
  NOR2_X1 U15941 ( .A1(n2709), .A2(n2154), .ZN(\mult_22/ab[2][55] ) );
  NOR2_X1 U15942 ( .A1(n2374), .A2(n2151), .ZN(\mult_22/ab[2][56] ) );
  NOR2_X1 U15943 ( .A1(n751), .A2(n2156), .ZN(\mult_22/ab[2][57] ) );
  NOR2_X1 U15944 ( .A1(n2720), .A2(n2155), .ZN(\mult_22/ab[2][58] ) );
  NOR2_X1 U15945 ( .A1(n2726), .A2(n2150), .ZN(\mult_22/ab[2][59] ) );
  NOR2_X1 U15946 ( .A1(n2413), .A2(n2157), .ZN(\mult_22/ab[2][5] ) );
  NOR2_X1 U15947 ( .A1(n748), .A2(n2153), .ZN(\mult_22/ab[2][60] ) );
  NOR2_X1 U15948 ( .A1(n2742), .A2(n2149), .ZN(\mult_22/ab[2][62] ) );
  NOR2_X1 U15949 ( .A1(n2751), .A2(n2148), .ZN(\mult_22/ab[2][63] ) );
  BUF_X1 U15950 ( .A(n2368), .Z(n2369) );
  NOR2_X1 U15951 ( .A1(n2703), .A2(n2950), .ZN(\mult_22/ab[35][54] ) );
  NOR2_X1 U15952 ( .A1(n2703), .A2(n2944), .ZN(\mult_22/ab[34][54] ) );
  NOR2_X1 U15953 ( .A1(n2703), .A2(n2938), .ZN(\mult_22/ab[33][54] ) );
  NOR2_X1 U15954 ( .A1(n2703), .A2(n2932), .ZN(\mult_22/ab[32][54] ) );
  NOR2_X1 U15955 ( .A1(n2703), .A2(n2926), .ZN(\mult_22/ab[31][54] ) );
  NOR2_X1 U15956 ( .A1(n2703), .A2(n2920), .ZN(\mult_22/ab[30][54] ) );
  NOR2_X1 U15957 ( .A1(n2703), .A2(n2155), .ZN(\mult_22/ab[2][54] ) );
  NOR2_X1 U15958 ( .A1(n2703), .A2(n2914), .ZN(\mult_22/ab[29][54] ) );
  NOR2_X1 U15959 ( .A1(n2703), .A2(n2908), .ZN(\mult_22/ab[28][54] ) );
  NOR2_X1 U15960 ( .A1(n2703), .A2(n2902), .ZN(\mult_22/ab[27][54] ) );
  NOR2_X1 U15961 ( .A1(n2703), .A2(n2896), .ZN(\mult_22/ab[26][54] ) );
  NOR2_X1 U15962 ( .A1(n2703), .A2(n2890), .ZN(\mult_22/ab[25][54] ) );
  OAI21_X1 U15963 ( .B1(n718), .B2(n717), .A(n976), .ZN(
        \mult_22/CARRYB[18][40] ) );
  NAND2_X1 U15964 ( .A1(reg_mid_1[10]), .A2(n3501), .ZN(n891) );
  NAND2_X1 U15965 ( .A1(reg_mid_1[15]), .A2(n3501), .ZN(n844) );
  NAND2_X1 U15966 ( .A1(reg_mid_1[17]), .A2(n3501), .ZN(n848) );
  NAND2_X1 U15967 ( .A1(reg_mid_1[21]), .A2(n3501), .ZN(n855) );
  NAND2_X1 U15968 ( .A1(reg_mid_1[27]), .A2(n3501), .ZN(n898) );
  NAND2_X1 U15969 ( .A1(reg_mid_1[30]), .A2(n3501), .ZN(n905) );
  NAND2_X1 U15970 ( .A1(reg_mid_1[32]), .A2(n3501), .ZN(n906) );
  NAND2_X1 U15971 ( .A1(reg_mid_1[34]), .A2(n3501), .ZN(n813) );
  NAND2_X1 U15972 ( .A1(reg_mid_1[37]), .A2(n3501), .ZN(n819) );
  NAND2_X1 U15973 ( .A1(reg_mid_1[39]), .A2(n3501), .ZN(n823) );
  NAND2_X1 U15974 ( .A1(reg_mid_1[48]), .A2(n2188), .ZN(n829) );
  NAND2_X1 U15975 ( .A1(reg_mid_1[58]), .A2(n2189), .ZN(n911) );
  INV_X1 U15976 ( .A(n2322), .ZN(n3512) );
  NAND2_X1 U15977 ( .A1(reg_mid_1[49]), .A2(n2120), .ZN(n828) );
  NAND2_X1 U15978 ( .A1(reg_mid_1[51]), .A2(n2120), .ZN(n882) );
  NAND2_X1 U15979 ( .A1(reg_mid_1[53]), .A2(n2293), .ZN(n883) );
  NOR3_X1 U15980 ( .A1(n2699), .A2(n3496), .A3(n872), .ZN(\mult_22/n7 ) );
  NOR2_X1 U15981 ( .A1(n2700), .A2(n2800), .ZN(\mult_22/ab[10][53] ) );
  NOR2_X1 U15982 ( .A1(n2697), .A2(n2794), .ZN(\mult_22/ab[9][53] ) );
  NOR2_X1 U15983 ( .A1(n2697), .A2(n2787), .ZN(\mult_22/ab[8][53] ) );
  NOR2_X1 U15984 ( .A1(n2697), .A2(n2782), .ZN(\mult_22/ab[7][53] ) );
  NOR2_X1 U15985 ( .A1(n2696), .A2(n2776), .ZN(\mult_22/ab[6][53] ) );
  NOR2_X1 U15986 ( .A1(n2700), .A2(n3118), .ZN(\mult_22/ab[63][53] ) );
  NOR2_X1 U15987 ( .A1(n2695), .A2(n3112), .ZN(\mult_22/ab[62][53] ) );
  NOR2_X1 U15988 ( .A1(n2697), .A2(n3106), .ZN(\mult_22/ab[61][53] ) );
  NOR2_X1 U15989 ( .A1(n2696), .A2(n3100), .ZN(\mult_22/ab[60][53] ) );
  NOR2_X1 U15990 ( .A1(n2696), .A2(n2770), .ZN(\mult_22/ab[5][53] ) );
  OAI21_X1 U15991 ( .B1(n727), .B2(n726), .A(n977), .ZN(
        \mult_22/CARRYB[11][46] ) );
  OAI211_X1 U15992 ( .C1(\mult_22/CARRYB[10][46] ), .C2(\mult_22/SUMB[10][47] ), .A(reg_mid_1[46]), .B(reg_mid_0[11]), .ZN(n977) );
  INV_X1 U15993 ( .A(n3499), .ZN(n2371) );
  INV_X1 U15994 ( .A(n3498), .ZN(n3494) );
  INV_X1 U15995 ( .A(n3497), .ZN(n3492) );
  INV_X1 U15996 ( .A(n3497), .ZN(n3495) );
  NOR2_X1 U15997 ( .A1(n911), .A2(n912), .ZN(\mult_22/CARRYB[1][58] ) );
  NOR2_X1 U15998 ( .A1(n903), .A2(n912), .ZN(\mult_22/n163 ) );
  OAI21_X1 U15999 ( .B1(n738), .B2(n737), .A(n960), .ZN(
        \mult_22/CARRYB[4][52] ) );
  INV_X1 U16000 ( .A(n3511), .ZN(n3500) );
  INV_X1 U16001 ( .A(n3511), .ZN(n3501) );
  CLKBUF_X1 U16002 ( .A(n3512), .Z(n3506) );
  CLKBUF_X1 U16003 ( .A(n3512), .Z(n3504) );
  CLKBUF_X1 U16004 ( .A(n3512), .Z(n3505) );
  CLKBUF_X1 U16005 ( .A(n3512), .Z(n3507) );
  CLKBUF_X1 U16006 ( .A(n3512), .Z(n3508) );
  CLKBUF_X1 U16007 ( .A(n3512), .Z(n3509) );
  CLKBUF_X1 U16008 ( .A(n3512), .Z(n3510) );
  CLKBUF_X1 U16009 ( .A(n3512), .Z(n3503) );
  OR2_X1 U16010 ( .A1(n2372), .A2(n2368), .ZN(n913) );
  OAI211_X1 U16011 ( .C1(\mult_22/SUMB[21][39] ), .C2(n2183), .A(reg_mid_1[38]), .B(reg_mid_0[22]), .ZN(n973) );
  XNOR2_X1 U16012 ( .A(\mult_22/SUMB[20][39] ), .B(\mult_22/CARRYB[20][38] ), 
        .ZN(n950) );
  OAI211_X1 U16013 ( .C1(\mult_22/CARRYB[3][52] ), .C2(\mult_22/SUMB[3][53] ), 
        .A(reg_mid_1[52]), .B(reg_mid_0[4]), .ZN(n960) );
  INV_X1 U16014 ( .A(\mult_22/CARRYB[3][52] ), .ZN(n737) );
  NOR2_X1 U16015 ( .A1(n887), .A2(n2364), .ZN(\mult_22/n59 ) );
  NAND2_X1 U16016 ( .A1(reg_mid_1[3]), .A2(n3494), .ZN(n860) );
  NAND2_X1 U16017 ( .A1(reg_mid_1[4]), .A2(n3492), .ZN(n862) );
  NAND2_X1 U16018 ( .A1(reg_mid_1[7]), .A2(n2139), .ZN(n864) );
  NAND2_X1 U16019 ( .A1(reg_mid_1[15]), .A2(n2139), .ZN(n866) );
  NAND2_X1 U16020 ( .A1(reg_mid_1[20]), .A2(n3493), .ZN(n868) );
  NAND2_X1 U16021 ( .A1(reg_mid_1[40]), .A2(n3495), .ZN(n822) );
  NAND2_X1 U16022 ( .A1(reg_mid_1[43]), .A2(n2371), .ZN(n824) );
  NAND2_X1 U16023 ( .A1(reg_mid_1[45]), .A2(n3493), .ZN(n826) );
  NAND2_X1 U16024 ( .A1(reg_mid_0[0]), .A2(reg_mid_1[63]), .ZN(n901) );
  NAND2_X1 U16025 ( .A1(reg_mid_1[60]), .A2(reg_mid_0[0]), .ZN(n910) );
  NAND2_X1 U16026 ( .A1(reg_mid_0[0]), .A2(reg_mid_1[58]), .ZN(n886) );
  INV_X1 U16027 ( .A(reg_mid_1[56]), .ZN(n2374) );
  CLKBUF_X1 U16028 ( .A(n752), .Z(n2715) );
  OR2_X1 U16029 ( .A1(n2142), .A2(n2376), .ZN(n876) );
  OAI211_X1 U16030 ( .C1(n1418), .C2(n1419), .A(n2121), .B(n1421), .ZN(n2378)
         );
  NOR3_X1 U16031 ( .A1(n884), .A2(n2369), .A3(n2698), .ZN(\mult_22/n6 ) );
  NAND2_X1 U16032 ( .A1(reg_mid_1[54]), .A2(reg_mid_0[0]), .ZN(n884) );
  NOR2_X1 U16033 ( .A1(n2712), .A2(n2860), .ZN(\mult_22/ab[20][56] ) );
  NOR2_X1 U16034 ( .A1(n2712), .A2(n2854), .ZN(\mult_22/ab[19][56] ) );
  NOR2_X1 U16035 ( .A1(n2712), .A2(n2848), .ZN(\mult_22/ab[18][56] ) );
  NOR2_X1 U16036 ( .A1(n2712), .A2(n2842), .ZN(\mult_22/ab[17][56] ) );
  NOR2_X1 U16037 ( .A1(n2712), .A2(n2836), .ZN(\mult_22/ab[16][56] ) );
  NOR2_X1 U16038 ( .A1(n2712), .A2(n2830), .ZN(\mult_22/ab[15][56] ) );
  NOR2_X1 U16039 ( .A1(n2712), .A2(n2824), .ZN(\mult_22/ab[14][56] ) );
  NOR2_X1 U16040 ( .A1(n2712), .A2(n2818), .ZN(\mult_22/ab[13][56] ) );
  NOR2_X1 U16041 ( .A1(n2712), .A2(n2812), .ZN(\mult_22/ab[12][56] ) );
  NOR2_X1 U16042 ( .A1(n2712), .A2(n2806), .ZN(\mult_22/ab[11][56] ) );
  NOR2_X1 U16043 ( .A1(n2715), .A2(n2800), .ZN(\mult_22/ab[10][56] ) );
  NAND2_X1 U16044 ( .A1(reg_mid_1[1]), .A2(n3492), .ZN(n1634) );
  NAND2_X1 U16045 ( .A1(reg_mid_1[25]), .A2(n2371), .ZN(n923) );
  NAND2_X1 U16046 ( .A1(reg_mid_1[26]), .A2(n3493), .ZN(n924) );
  NAND2_X1 U16047 ( .A1(reg_mid_1[27]), .A2(n3495), .ZN(n925) );
  NAND2_X1 U16048 ( .A1(reg_mid_1[28]), .A2(n2139), .ZN(n926) );
  NAND2_X1 U16049 ( .A1(reg_mid_1[29]), .A2(n2139), .ZN(n927) );
  NAND2_X1 U16050 ( .A1(reg_mid_1[30]), .A2(n2371), .ZN(n928) );
  NAND2_X1 U16051 ( .A1(reg_mid_1[31]), .A2(n3495), .ZN(n929) );
  NAND2_X1 U16052 ( .A1(reg_mid_1[33]), .A2(n3495), .ZN(n930) );
  NAND2_X1 U16053 ( .A1(reg_mid_1[52]), .A2(n2293), .ZN(n880) );
  NAND2_X1 U16054 ( .A1(reg_mid_0[0]), .A2(reg_mid_1[59]), .ZN(n912) );
  NOR2_X1 U16055 ( .A1(n2375), .A2(n2377), .ZN(\mult_22/ab[0][56] ) );
  NOR2_X1 U16056 ( .A1(n2706), .A2(n3118), .ZN(\mult_22/ab[63][55] ) );
  NOR2_X1 U16057 ( .A1(n2706), .A2(n3112), .ZN(\mult_22/ab[62][55] ) );
  NOR2_X1 U16058 ( .A1(n2706), .A2(n3106), .ZN(\mult_22/ab[61][55] ) );
  NOR2_X1 U16059 ( .A1(n2706), .A2(n3100), .ZN(\mult_22/ab[60][55] ) );
  NOR2_X1 U16060 ( .A1(n2706), .A2(n3094), .ZN(\mult_22/ab[59][55] ) );
  NOR2_X1 U16061 ( .A1(n2706), .A2(n3088), .ZN(\mult_22/ab[58][55] ) );
  NOR2_X1 U16062 ( .A1(n2706), .A2(n2800), .ZN(\mult_22/ab[10][55] ) );
  NOR2_X1 U16063 ( .A1(n2706), .A2(n2788), .ZN(\mult_22/ab[8][55] ) );
  NOR2_X1 U16064 ( .A1(n2706), .A2(n2782), .ZN(\mult_22/ab[7][55] ) );
  NOR2_X1 U16065 ( .A1(n2706), .A2(n2776), .ZN(\mult_22/ab[6][55] ) );
  NOR2_X1 U16066 ( .A1(n2706), .A2(n2770), .ZN(\mult_22/ab[5][55] ) );
  NOR2_X1 U16067 ( .A1(n2376), .A2(n2373), .ZN(\mult_22/ab[1][55] ) );
  XNOR2_X1 U16068 ( .A(\mult_22/SUMB[10][47] ), .B(\mult_22/CARRYB[10][46] ), 
        .ZN(n958) );
  NOR3_X1 U16069 ( .A1(n876), .A2(n2369), .A3(n2370), .ZN(\mult_22/n324 ) );
  INV_X1 U16070 ( .A(\mult_22/CARRYB[7][50] ), .ZN(n731) );
  OAI21_X1 U16071 ( .B1(n732), .B2(n731), .A(n959), .ZN(
        \mult_22/CARRYB[8][50] ) );
  NAND2_X1 U16072 ( .A1(n1471), .A2(n2348), .ZN(n1469) );
  INV_X1 U16073 ( .A(n1467), .ZN(n603) );
  INV_X1 U16074 ( .A(n1482), .ZN(n601) );
  OAI211_X1 U16075 ( .C1(n1400), .C2(n1401), .A(n1402), .B(n1403), .ZN(n1398)
         );
  AND2_X1 U16076 ( .A1(n2089), .A2(n2379), .ZN(n1422) );
  AOI21_X1 U16077 ( .B1(n1616), .B2(n622), .A(n623), .ZN(n1609) );
  OAI21_X1 U16078 ( .B1(n1332), .B2(n1331), .A(n1333), .ZN(n1325) );
  NAND2_X1 U16079 ( .A1(n594), .A2(n622), .ZN(n1615) );
  OAI21_X1 U16080 ( .B1(n1342), .B2(n1341), .A(n1343), .ZN(n1335) );
  OAI211_X1 U16081 ( .C1(n1467), .C2(n1468), .A(n1469), .B(n1470), .ZN(n1465)
         );
  NAND2_X1 U16082 ( .A1(reg_mid_1[4]), .A2(n3502), .ZN(n890) );
  NAND2_X1 U16083 ( .A1(reg_mid_1[41]), .A2(n3501), .ZN(n888) );
  NAND2_X1 U16084 ( .A1(reg_mid_1[43]), .A2(n3500), .ZN(n889) );
  NAND2_X1 U16085 ( .A1(reg_mid_1[49]), .A2(n2189), .ZN(n830) );
  NAND2_X1 U16086 ( .A1(reg_mid_1[59]), .A2(n2188), .ZN(n909) );
  NAND2_X1 U16087 ( .A1(reg_mid_1[52]), .A2(n2189), .ZN(n872) );
  NAND2_X1 U16088 ( .A1(reg_mid_1[56]), .A2(n2189), .ZN(n887) );
  NAND2_X1 U16089 ( .A1(reg_mid_1[53]), .A2(n2188), .ZN(n885) );
  NOR2_X1 U16090 ( .A1(n612), .A2(n1422), .ZN(n1433) );
  OAI21_X1 U16091 ( .B1(n1322), .B2(n1321), .A(n1323), .ZN(n1316) );
  OAI211_X1 U16092 ( .C1(n708), .C2(\mult_22/CARRYB[22][37] ), .A(
        reg_mid_1[37]), .B(reg_mid_0[23]), .ZN(n969) );
  INV_X1 U16093 ( .A(\mult_22/CARRYB[10][46] ), .ZN(n726) );
  OAI21_X1 U16094 ( .B1(n1549), .B2(n1548), .A(n1550), .ZN(n1542) );
  OAI211_X1 U16095 ( .C1(n1563), .C2(n1564), .A(n1565), .B(n1566), .ZN(n1561)
         );
  OAI21_X1 U16096 ( .B1(n1453), .B2(n1452), .A(n1454), .ZN(n1446) );
  OAI21_X1 U16097 ( .B1(n1362), .B2(n1361), .A(n1363), .ZN(n1355) );
  OAI211_X1 U16098 ( .C1(\mult_22/SUMB[20][39] ), .C2(\mult_22/CARRYB[20][38] ), .A(reg_mid_1[38]), .B(reg_mid_0[21]), .ZN(n974) );
  OAI21_X1 U16099 ( .B1(n2083), .B2(n1442), .A(n1444), .ZN(n1439) );
  OAI221_X1 U16100 ( .B1(n1371), .B2(n1372), .C1(n1374), .C2(n1373), .A(n1375), 
        .ZN(n1365) );
  AOI21_X1 U16101 ( .B1(n1295), .B2(n646), .A(n1296), .ZN(n1290) );
  OAI22_X1 U16102 ( .A1(n1290), .A2(n650), .B1(n1291), .B2(n1292), .ZN(n1283)
         );
  AOI21_X1 U16103 ( .B1(n1561), .B2(n584), .A(n1562), .ZN(n1560) );
  AOI21_X1 U16104 ( .B1(n1465), .B2(n604), .A(n1466), .ZN(n1464) );
  AOI21_X1 U16105 ( .B1(\mult_22/CARRYB[63][1] ), .B2(\mult_22/SUMB[63][2] ), 
        .A(n2354), .ZN(n1629) );
  INV_X1 U16106 ( .A(\mult_22/CARRYB[17][40] ), .ZN(n717) );
  OAI21_X1 U16107 ( .B1(n1352), .B2(n1351), .A(n1353), .ZN(n1345) );
  OAI211_X1 U16108 ( .C1(n1583), .C2(n1584), .A(n1586), .B(n1585), .ZN(n1567)
         );
  INV_X1 U16109 ( .A(n974), .ZN(n712) );
  OAI22_X1 U16110 ( .A1(n1311), .A2(n643), .B1(n1312), .B2(n1313), .ZN(n1304)
         );
  AOI21_X1 U16111 ( .B1(n1316), .B2(n642), .A(n1317), .ZN(n1311) );
  AOI21_X1 U16112 ( .B1(n1283), .B2(n651), .A(n1284), .ZN(n1282) );
  AOI21_X1 U16113 ( .B1(n2232), .B2(n626), .A(n627), .ZN(n1389) );
  AOI21_X1 U16114 ( .B1(n582), .B2(n2341), .A(n581), .ZN(n1576) );
  AOI21_X1 U16115 ( .B1(n617), .B2(n2378), .A(n618), .ZN(n1412) );
  AOI21_X1 U16116 ( .B1(n1491), .B2(n1507), .A(n1498), .ZN(n1505) );
  OAI21_X1 U16117 ( .B1(n1629), .B2(n1613), .A(n2169), .ZN(n1625) );
  AOI21_X1 U16118 ( .B1(n2366), .B2(n1604), .A(n1594), .ZN(n1601) );
  AOI21_X1 U16119 ( .B1(n1365), .B2(n631), .A(n1366), .ZN(n1362) );
  NAND2_X1 U16120 ( .A1(n1376), .A2(n626), .ZN(n1374) );
  AOI21_X1 U16121 ( .B1(n1456), .B2(n606), .A(n1457), .ZN(n1453) );
  INV_X1 U16122 ( .A(n1629), .ZN(n594) );
  INV_X1 U16123 ( .A(\mult_22/SUMB[32][29] ), .ZN(n687) );
  OAI211_X1 U16124 ( .C1(\mult_22/CARRYB[32][28] ), .C2(\mult_22/SUMB[32][29] ), .A(reg_mid_1[28]), .B(reg_mid_0[33]), .ZN(n962) );
  OAI21_X1 U16125 ( .B1(n941), .B2(n698), .A(n696), .ZN(
        \mult_22/CARRYB[26][34] ) );
  INV_X1 U16126 ( .A(n964), .ZN(n696) );
  AOI211_X1 U16127 ( .C1(n698), .C2(n941), .A(n2588), .B(n2892), .ZN(n964) );
  INV_X1 U16128 ( .A(n946), .ZN(n708) );
  XNOR2_X1 U16129 ( .A(n947), .B(n946), .ZN(\mult_22/SUMB[23][37] ) );
  INV_X1 U16130 ( .A(\mult_22/SUMB[17][41] ), .ZN(n718) );
  OAI211_X1 U16131 ( .C1(\mult_22/CARRYB[17][40] ), .C2(\mult_22/SUMB[17][41] ), .A(reg_mid_1[40]), .B(reg_mid_0[18]), .ZN(n976) );
  NAND2_X1 U16132 ( .A1(reg_mid_1[2]), .A2(n3500), .ZN(n861) );
  NAND2_X1 U16133 ( .A1(reg_mid_1[3]), .A2(n3501), .ZN(n863) );
  NAND2_X1 U16134 ( .A1(reg_mid_1[6]), .A2(n3501), .ZN(n865) );
  NAND2_X1 U16135 ( .A1(reg_mid_1[14]), .A2(n3500), .ZN(n867) );
  NAND2_X1 U16136 ( .A1(reg_mid_1[19]), .A2(n3501), .ZN(n869) );
  NAND2_X1 U16137 ( .A1(reg_mid_1[31]), .A2(n3502), .ZN(n871) );
  NAND2_X1 U16138 ( .A1(reg_mid_1[33]), .A2(n3502), .ZN(n811) );
  NAND2_X1 U16139 ( .A1(reg_mid_1[40]), .A2(n3502), .ZN(n874) );
  NAND2_X1 U16140 ( .A1(reg_mid_1[51]), .A2(n2188), .ZN(n881) );
  NAND2_X1 U16141 ( .A1(reg_mid_1[50]), .A2(n2189), .ZN(n851) );
  NAND2_X1 U16142 ( .A1(reg_mid_1[54]), .A2(n2188), .ZN(n877) );
  CLKBUF_X1 U16143 ( .A(n1876), .Z(n2385) );
  CLKBUF_X1 U16144 ( .A(n1855), .Z(n2391) );
  CLKBUF_X1 U16145 ( .A(n1854), .Z(n2397) );
  CLKBUF_X1 U16146 ( .A(n1853), .Z(n2403) );
  CLKBUF_X1 U16147 ( .A(n1875), .Z(n2409) );
  CLKBUF_X1 U16148 ( .A(n1847), .Z(n2415) );
  CLKBUF_X1 U16149 ( .A(n1846), .Z(n2421) );
  CLKBUF_X1 U16150 ( .A(n1832), .Z(n2427) );
  CLKBUF_X1 U16151 ( .A(n1845), .Z(n2433) );
  CLKBUF_X1 U16152 ( .A(n1844), .Z(n2439) );
  CLKBUF_X1 U16153 ( .A(n1874), .Z(n2445) );
  CLKBUF_X1 U16154 ( .A(n1861), .Z(n2451) );
  CLKBUF_X1 U16155 ( .A(n1863), .Z(n2457) );
  CLKBUF_X1 U16156 ( .A(n1837), .Z(n2463) );
  CLKBUF_X1 U16157 ( .A(n1843), .Z(n2469) );
  CLKBUF_X1 U16158 ( .A(n1835), .Z(n2475) );
  CLKBUF_X1 U16159 ( .A(n1836), .Z(n2481) );
  CLKBUF_X1 U16160 ( .A(n1842), .Z(n2487) );
  CLKBUF_X1 U16161 ( .A(n1841), .Z(n2493) );
  CLKBUF_X1 U16162 ( .A(n1840), .Z(n2499) );
  CLKBUF_X1 U16163 ( .A(n1839), .Z(n2505) );
  CLKBUF_X1 U16164 ( .A(n1838), .Z(n2511) );
  CLKBUF_X1 U16165 ( .A(n1834), .Z(n2517) );
  CLKBUF_X1 U16166 ( .A(n1833), .Z(n2523) );
  CLKBUF_X1 U16167 ( .A(n1873), .Z(n2529) );
  CLKBUF_X1 U16168 ( .A(n1864), .Z(n2535) );
  CLKBUF_X1 U16169 ( .A(n1862), .Z(n2541) );
  CLKBUF_X1 U16170 ( .A(n1865), .Z(n2547) );
  CLKBUF_X1 U16171 ( .A(n1868), .Z(n2553) );
  CLKBUF_X1 U16172 ( .A(n1856), .Z(n2559) );
  CLKBUF_X1 U16173 ( .A(n1823), .Z(n2565) );
  CLKBUF_X1 U16174 ( .A(n1816), .Z(n2571) );
  CLKBUF_X1 U16175 ( .A(n1817), .Z(n2582) );
  CLKBUF_X1 U16176 ( .A(n1819), .Z(n2588) );
  CLKBUF_X1 U16177 ( .A(n1811), .Z(n2594) );
  CLKBUF_X1 U16178 ( .A(n1815), .Z(n2600) );
  CLKBUF_X1 U16179 ( .A(n1814), .Z(n2606) );
  CLKBUF_X1 U16180 ( .A(n1820), .Z(n2617) );
  CLKBUF_X1 U16181 ( .A(n1812), .Z(n2623) );
  CLKBUF_X1 U16182 ( .A(n1824), .Z(n2629) );
  CLKBUF_X1 U16183 ( .A(n1818), .Z(n2635) );
  CLKBUF_X1 U16184 ( .A(n1825), .Z(n2641) );
  CLKBUF_X1 U16185 ( .A(n1813), .Z(n2647) );
  CLKBUF_X1 U16186 ( .A(n2362), .Z(n2653) );
  CLKBUF_X1 U16187 ( .A(n2363), .Z(n2659) );
  CLKBUF_X1 U16188 ( .A(n2361), .Z(n2665) );
  CLKBUF_X1 U16189 ( .A(n2360), .Z(n2671) );
  CLKBUF_X1 U16190 ( .A(n1826), .Z(n2677) );
  CLKBUF_X1 U16191 ( .A(n2359), .Z(n2683) );
  CLKBUF_X1 U16192 ( .A(n1821), .Z(n2689) );
  CLKBUF_X1 U16193 ( .A(n754), .Z(n2705) );
  CLKBUF_X1 U16194 ( .A(n753), .Z(n2711) );
  CLKBUF_X1 U16195 ( .A(n1822), .Z(n2724) );
  CLKBUF_X1 U16196 ( .A(n2140), .Z(n2730) );
  CLKBUF_X1 U16197 ( .A(n748), .Z(n2736) );
  CLKBUF_X1 U16198 ( .A(n746), .Z(n2747) );
  CLKBUF_X1 U16199 ( .A(n2111), .Z(n2753) );
  CLKBUF_X1 U16200 ( .A(n1810), .Z(n2759) );
  CLKBUF_X1 U16201 ( .A(n1827), .Z(n2765) );
  CLKBUF_X1 U16202 ( .A(n1829), .Z(n2771) );
  CLKBUF_X1 U16203 ( .A(n1828), .Z(n2777) );
  CLKBUF_X1 U16204 ( .A(n1878), .Z(n2783) );
  CLKBUF_X1 U16205 ( .A(n1877), .Z(n2789) );
  CLKBUF_X1 U16206 ( .A(n1866), .Z(n2795) );
  CLKBUF_X1 U16207 ( .A(n1872), .Z(n2801) );
  CLKBUF_X1 U16208 ( .A(n1871), .Z(n2807) );
  CLKBUF_X1 U16209 ( .A(n1851), .Z(n2813) );
  CLKBUF_X1 U16210 ( .A(n1850), .Z(n2819) );
  CLKBUF_X1 U16211 ( .A(n1849), .Z(n2825) );
  CLKBUF_X1 U16212 ( .A(n1848), .Z(n2831) );
  CLKBUF_X1 U16213 ( .A(n1867), .Z(n2837) );
  CLKBUF_X1 U16214 ( .A(n1870), .Z(n2843) );
  CLKBUF_X1 U16215 ( .A(n1869), .Z(n2849) );
  CLKBUF_X1 U16216 ( .A(n1852), .Z(n2855) );
  CLKBUF_X1 U16217 ( .A(n1859), .Z(n2861) );
  CLKBUF_X1 U16218 ( .A(n1857), .Z(n2867) );
  CLKBUF_X1 U16219 ( .A(n1858), .Z(n2873) );
  CLKBUF_X1 U16220 ( .A(n1887), .Z(n2879) );
  CLKBUF_X1 U16221 ( .A(n1886), .Z(n2885) );
  CLKBUF_X1 U16222 ( .A(n1893), .Z(n2891) );
  CLKBUF_X1 U16223 ( .A(n1860), .Z(n2897) );
  CLKBUF_X1 U16224 ( .A(n1892), .Z(n2903) );
  CLKBUF_X1 U16225 ( .A(n1891), .Z(n2909) );
  CLKBUF_X1 U16226 ( .A(n1890), .Z(n2915) );
  CLKBUF_X1 U16227 ( .A(n1889), .Z(n2921) );
  CLKBUF_X1 U16228 ( .A(n1900), .Z(n2927) );
  CLKBUF_X1 U16229 ( .A(n1888), .Z(n2933) );
  CLKBUF_X1 U16230 ( .A(n1899), .Z(n2939) );
  CLKBUF_X1 U16231 ( .A(n1898), .Z(n2945) );
  CLKBUF_X1 U16232 ( .A(n1897), .Z(n2951) );
  CLKBUF_X1 U16233 ( .A(n1894), .Z(n2957) );
  CLKBUF_X1 U16234 ( .A(n1895), .Z(n2963) );
  CLKBUF_X1 U16235 ( .A(n1896), .Z(n2969) );
  CLKBUF_X1 U16236 ( .A(n1927), .Z(n2975) );
  CLKBUF_X1 U16237 ( .A(n1928), .Z(n2981) );
  CLKBUF_X1 U16238 ( .A(n1929), .Z(n2987) );
  CLKBUF_X1 U16239 ( .A(n1930), .Z(n2993) );
  CLKBUF_X1 U16240 ( .A(n1931), .Z(n2999) );
  CLKBUF_X1 U16241 ( .A(n1932), .Z(n3005) );
  CLKBUF_X1 U16242 ( .A(n1934), .Z(n3011) );
  CLKBUF_X1 U16243 ( .A(n1933), .Z(n3017) );
  CLKBUF_X1 U16244 ( .A(n1995), .Z(n3023) );
  CLKBUF_X1 U16245 ( .A(n1997), .Z(n3029) );
  CLKBUF_X1 U16246 ( .A(n1996), .Z(n3035) );
  CLKBUF_X1 U16247 ( .A(n1998), .Z(n3041) );
  CLKBUF_X1 U16248 ( .A(n1999), .Z(n3047) );
  CLKBUF_X1 U16249 ( .A(n2000), .Z(n3053) );
  CLKBUF_X1 U16250 ( .A(n2001), .Z(n3059) );
  CLKBUF_X1 U16251 ( .A(n2003), .Z(n3065) );
  CLKBUF_X1 U16252 ( .A(n2002), .Z(n3071) );
  CLKBUF_X1 U16253 ( .A(n2021), .Z(n3077) );
  CLKBUF_X1 U16254 ( .A(n2020), .Z(n3083) );
  CLKBUF_X1 U16255 ( .A(n2027), .Z(n3089) );
  CLKBUF_X1 U16256 ( .A(n2026), .Z(n3095) );
  CLKBUF_X1 U16257 ( .A(n2025), .Z(n3101) );
  CLKBUF_X1 U16258 ( .A(n2024), .Z(n3107) );
  CLKBUF_X1 U16259 ( .A(n2023), .Z(n3113) );
  CLKBUF_X1 U16260 ( .A(n2022), .Z(n3119) );
  INV_X1 U16261 ( .A(n1935), .ZN(n3515) );
  INV_X1 U16262 ( .A(n1936), .ZN(n3526) );
endmodule

